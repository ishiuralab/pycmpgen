module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [10:0] src12;
    reg [9:0] src13;
    reg [8:0] src14;
    reg [7:0] src15;
    reg [6:0] src16;
    reg [5:0] src17;
    reg [4:0] src18;
    reg [3:0] src19;
    reg [2:0] src20;
    reg [1:0] src21;
    reg [0:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3])<<19) + ((src20[0] + src20[1] + src20[2])<<20) + ((src21[0] + src21[1])<<21) + ((src22[0])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5da8b71eabc896107e14dd93766a46e0cefe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22808a17a999039cad23f2f6c07543ce5368;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h727a7d1f69c5bf73badd52f09469bd1b9201;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6486d4335a38ccb12e6d85b4b7dd6ce800e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5c14a673b71af299f792a5b09f1c62640ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb572ab553b43cf046e119d9dc70b4a660;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35e02984a18fa094d2dc2459f1087c14e503;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd824f43e558d2d9b9fe989ccbfcbd1d36c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbee0405c59258d41f2cd957a989616f99ed4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e290ecf58e499a32e41002f784cd181bcef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd34d00e20140dfda26a0af035afe1a107af4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4065b9c3f27839781cd05445bcbc5ea7e02b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53234d3533f14e6e2a9170c2db93e0aae0de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51a24c3dc14f2153594bb11e6da1edf5356b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3127f6bb5316a8655a442362a5372e095e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcaf9e1e9e616ee0a92dcfe708c484ffc6f68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aa041c4457012605345eca94639754286ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dc228bf5fdb1294873628e10569d457aac7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56799ea8145bdb3aadb402b218564014a015;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefc5bcb4b630b741fb4c375f8015c6c394f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h998199e0c25f910174b2cacf7ab1ec4def1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e85f1e2638440bb887061236a8f5472adc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae6437d319d52a8d2374683808ffbdf5b2ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc19291443a82033382c4be3ef16dc2d4e26e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h767f368c259f9a6a29171e446610b9587bca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c9748a1bba201526f0a9c9ca6920899d03a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha65c9112f6d660bbed132d57f9d6d1aaaacf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he31311cb1994be203afa417a64ededd8f525;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h529795df8d2bcbc7b4575bd0115937306410;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e12172d8f4e2d9d5ceb787cc07bc127571c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha86c13af4a4f28a1c591cf375304ed3459f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb29f36b947dcdfd6e1ba2eee54ade97fa85d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb13defc2673d3bd347b58001b57091f66138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90ba3a47ca38851a8d54e38044a376b24f1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d989e881beb0a4e3809d993acb992ef2819;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he042b892fcf12e0cd2871de2629238127511;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd071d742d10e7d9ff39deb3c1b7cf6e5c499;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf581a9f4c350170dbb45a830cb043395f6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10d1eaa6ab80f4d17023e6b404745cd4b1ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c0c5cc8df31b517316cc9318d8e893e7a62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf993e51308d7a10bf9900dc0b8910e56514c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a331075c9a182eb3add4d5912e8151fcfca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he26f61450b1b7390d5d920e573d51b74fe83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hace464320afd6caaf6d0e0f3d537d2731335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1142e44c39b63613b0a8458f8e20b92a94d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb42b987d614090e1ea1cda35b4e1b8ad710a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he663ca8392265a00769d3f9e132f70359111;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h506cdecb5806b73d8e62dc65a851799084d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc670935c365c280ac44d47a0b26e222a908;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h721e62ad11c1c6f3932f98faa1714ecfcb61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha483bd69f5b8577f64842036a451ddf34182;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ffc23dd1dea597f505ad230e9d8882bad99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2896f90d4ebabb04c4142acb7ada4e4d1fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7930be806b28329de95bf716dcf0693d1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7e43db5e8409d1fe1de1f0e08bd9c7016f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72f2b22245707599d4c4b9e37682040b7170;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafec8dd04f65d824e64c6689790e82d83b0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10653bd3364e1a9dc11195d945447039534b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65027868cf3e4d44edcfed2ad2d2e79bdceb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67fc2f8bd3706053b3bb370ae3ba5d0b60ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3d51522f183e2e2fab4fadec53c24488c71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9e7428781d531f7463c6ae2fc29cad002fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d94c2af2742d8cf0997a93398b491c2ea05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0f2b32b22548ac8aa222f85697268dc397;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97415d6fb39cc30a25a00d9b87de2fc12335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h271730f6a55a9f9fd09d4576d973c015a17c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1458f63eeb1595f216d9678691e077936c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c453b84bed67533d19869b4319683151eb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7dd2358b80fa67206c8bd46a7d91c216dd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d1dee0d42737d167bfff5e29e7f91475b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3592f46836e97908c235c9b178f5204757b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3bf2b13589aeb7ea497d020590c911b9d6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d40c21c1e0296e926ad0822f0f3ea09e54e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee9ade52e378fa7b244654399090f0439e35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h309b195b030f2f3b5a027a17dbff9df4f47c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb40ff751dd09ddbc26fb55ed77dae1f2c28a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7fb16946a084c7bd7caeb81924bafbbe213;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25dc7fbb921bf4573366410c883e2a4bdad3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb96b154882ea4d83216a335c6e3dedda47a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd76320da45ac904f8abd363479ed5b4f2f48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h228182d1fea074f1a2eb3b73f8f0ed518e2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f2f055caeecde16a03ecdb8f70d189280ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f7923b50c6b7246e7cc5c32716796aab838;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c35aa29649f04b58c0838da0356aa561945;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae3d262a6e546072cbed519c3c800abaa412;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41292e8b3a2ac655589a1ddfd1c51c48c031;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd206c0e73b345b204af7b7a25ce350ae1fcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6764b24a583aa72ebf417c053f1e850f8190;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd6729a37ca7d81314e929e54330f26fe931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8352903439517b87a29662054ae99f2f464;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4159f853303cfce1c0fcfad1b5172b32c716;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ee71ef64da15bc851a18fd4d16953df0e37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c2639021a93aa87eec60347c44950a093fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb21dc2bf957d0cbb33998a20778a6d270cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h960ba0307136d7a49b2f1e274203f4e9ef80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd201a9dbc27a3070315af8a6858f811fb16c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76f43a4ce690b534be016e630566b166970f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62d5ca0fc2e277366f4450b75707babafaf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9887f59ad12ebc1bede3e510b3e6000b9f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49f8ad8e3de7b4bf95a4bf6d949be209a958;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99646ca2351457f28dc121aeb0b538aa06fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcd2965caf182dd6c2285ca8df785f6e4d56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2434a168393348ace14d96d02182119ecaff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cd93f107f0fe15de0d25a5fd5f0b2f8ea9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h773ee75f9386c673a0c802f538a7522fb074;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbeaa0889826cdd0eba4ea5b3beaadd779504;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf82759fea0a46c011f052f9f767d3c3b647f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42a79da751b1cb4a125e0d78aeed8fa4c6f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbaa5656a2ce4a7c0459474b51d6b7ed8ab19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe745703ca8d9fd1c0e22d767edf6464163;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cbbe56f84e39add1607d559c7258788557a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfbd25cedaccb7118d50bc203ce879d8853c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5379f34ec148638aec8e8028998ba45317b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4623e9d2c285fb49440bff73ed3c64789ca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ae10490a5f8436afc3e4c98c9c58ae4e08d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc961f9e06348c4697993b4882b95f5c0f52e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3d9153d14657b31167795b05f4da3e3063d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b838ed541cf4d10dbf74aa99442fbc50a28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49bb6ecbeeee6d980af392528ca19f90f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ad5a1e0dd5bc61b1187942a7ef85ed82c5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6e3abe49c55e9c58795fa00e05af10f8ee1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h125ef0d7e749e209f3c13631cbc15f60f0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ba9d7d93c89513968761615e30d0e5584f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c718f708f39fe32954381c763e4778b1e3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9cdd153694c40c4fc441270c8eed3ca9e8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aa3b4b6cc36387e1949576752af93d9836d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc86e0341b707d997521fbf03e2c2d1c5016e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3d926796c1da63282bd39882f325919cef8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28a5a4e808af88769ed53f6cb84cca4a0400;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b8e6b60485b4e6e50edb70b48c330bdde3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd223b6ace3cf41f1a46951e8cd74d5ec47e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59daad7d0ac74600f9c88225f936eed816e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6701b9b439e6ef24aba376af4e56c37d9e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3246efcaaef1ce3670af3e50ac0b6a1f938b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf144d66225452f4b6ffae90717eadf00dda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4d304e1dbb67bda6f22dbba6bfccd8a651b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32204c567f8077722afdcda73a9fe96d488b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h353e9de30dca55dbbd7c561198d09712614a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d627bc5820e2f8308a915b18c1f60ce8ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c32c31826e8d1479dc8d6171e0dc0b7081a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h301b0d74e942d2de449dabc6f3843641a439;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h750d878c0e0595ffd70e032f5c40306db90b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1594a03b9b2047c25b179369d8f250ea13d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2317b203e8887f8eb412a43cac73455b55c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97ba8bf7a72cb72ace4cb6f55a5ee464d2da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b9fb5656ca68c6dbf74cf38445a6fde34c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2c157d4b8ba1af95a029e8e7c5bd06e5a32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h214b441bf4ee730e78509c6cc5f75f846580;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81ce7d777481b9a02cc7ba6f0dd9944703df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b7d5c5cd2b6a0f076e1ac50b79e737b4bf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24caeaa1046eb9b246cc2a796d332ebe8e2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf968e96566f9a8bace96224939d6e4b3faa0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e33b09b19e438b5ce9007d63e8c0fe36208;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd54ae5b6d3bb82903f60837a0076db409f73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heed7b4451e2070514e2ed79200138b0d13ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha93f62cb1ec820d291d27d005d8a7f31b3ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f061eb0851df3e0015aed4aa904794861db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf236efcab34c1b7b07ad11b23c74149b738c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ecbac5bedc4ffb4d9c56e90ce6d69b57884;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he101eebf7183ec3b89151e5e6853c9877374;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeb0d7ac2a98b848daf453f2704bd7ee1ffb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd68edbc173583fd8882019cdbfa4512b87b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6492ec8b24ea808b23ca7e80fb3af0c85ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea56faa47b4abfee80f9e907c48396851030;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fe3ed7de11f894823f21ff6d1bb317104d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66c76d0773f09eb70f0b4620c7825dc88939;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10bb6927bd10272a91eedbb3d386f8a2c91d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a6049515cec6d5ae156d435e15b7c57cc0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h684b168a8c2829d47cc7956cfaf0ed42757b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d57be8e738d26842c9e86d9f38f70c4237f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f5482967a554975b6c1bcdb5545f15afff7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd3e08f159d903eac0c26d51058c78f98a69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b01859bac7152a98f5103b06d9f4c24527f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8314e1b10f60aa7fd52d867379b48b1af93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fd217831e29d7a1b4752149d86385951e9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fb2091c834dbd97e0772cd562cf16b64bd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d3787ea10963ddffb10e29b5f9ed168d63d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29368bdada4a8ded0092567e5ba34eb7b0ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c24cf77ba12087c00f58e7b7c46743a520e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ccab9fd9a05bbb5c96530dc552d2674514;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf895849a37e20054ea6f2598ddc6085843cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bdcd9c3743988b3faf5ab30d3c5e5ed7c9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60a261506037635b372d7e13b2cf2b335b41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h373253b5be7d933269495a35101bb60d317d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7adfadc9a5de79354cade644b175da6e7741;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d49acc6531b487a08b8fb8ccf5631da7731;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0e01a8e7e17fdee95979ab6bbc60f2f999;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h466d14f1602dc3db9cc23ca4dff483dba63b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ad1424a808ebc7f50a551f6271e41c4b096;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82865f6bac66a6412375efe962b190d691cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58dbbc1050e9f099b443d8ae400f7928c849;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96644b585bcfefc9ebd6ea5c3cd7f110fbdd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb323ec64be2546933bda073a392705c494d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56c978e30d6ea1ee597210d01946fa81caed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h960828d9b316ecf1d732d04e418cfd79d2c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cc3ef739770fc101756f2308052786d4bbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8560797004bdb449c395fa53b073fb3c8a00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58d08e868a43fdbd0d81a9298b7218b652ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfad6f1cf33615540fd0dd2c863d7df7be5c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1f510ef7cb900b341e12ce986383916a192;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68041141704c4f69bd7c3e9b9bdc7f4e51f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he034219e62649ca90e048e02a4eab56c7a94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62f7a4d00600140b6b7f8ca066ea8dda711;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0b26b5c49a7de9467464b289f4bbe46f113;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haca1ade9f9ca35cf7fe7e808921a0f80ac4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f52c45a11839f8f2719dda3ee83e672eabe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dd9956f27756d3dd9ba40e1ce3665fee738;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1dd536e00abd33a7fe5285c15f0b6f19a7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc66e2b41c9f13fe238c44a255f1a74e9764a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e0f74e84467bc6c38e34f18ff96245e9b60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8804965cccb73629f7c67027c996f07dce4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8788d99cb678426b5758f07f4bb34fefcfa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8241200ad29117fbc762581046f407e74b8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h997ced34e9663e720e1cef385f0094489879;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65b8ed81470a41038cbe3a366881e58bae5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf25fe4dcadfad551338115a3095250a06a9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff09196754c3e4ca134ab7ad716692eb479f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45ea03172c011bd96fb2d02cfe25d813348d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3fdae01f9f98a1f33f3486b7449dfd41e0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4e98f888b9dcaea51d7f2206676bf2b505a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35661352b9ad2448032d5b61fd13d4b89bb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f441f7fee8ed4e329a2e9279fdefbaa9b9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ef14015b8cc73e44321346e81510a352534;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a7f0fe8e45910808b61be421c8d12c1404c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he41f2f3968c24340bdcaf522aa512743d122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h397301f9402b3c209c6769555d4832e2e390;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e0b78ef4ad99cf07c12b0eabf9d8818d0f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e8f55dcad3f8bf265e7741df7f39fafc9df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0950ce7cc479099bb7894718d5d5d701d56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9529966f26d20ffb39a86ab8a2ce4eb63bc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd93bcf079764dee96bc55d89d9ee38ca9a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b9a0e8e185b93182c21864dc12ceea68fea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ff8ef2a9187767ba8d83cc7f45bc39e5fe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43a72e001622da0e22e6f50f58d16161aafa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1237103fd87b887c56d46cddaf2e3af23202;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h191b90e2e4e67b2701af945ec1e13dc78b5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90b1b5b6a91effb48b5b2d2e1464d4568b34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h679b9554949f45e9297aa63656fab925cd54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13930108ffa453255f08f7236c6e218278e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a055c3f8ee82b4c4d0c7b33c356775fac75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a03132d1e1080ff8b449e1d78698b51f26d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb0d63b0e2babd465f7f760d3275457d35b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he08f18def102de12edd9b6651455e6ee6a8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd80818c2fd349c8ba8d67c5d0d16c1f8fb47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ef3ea712b432b407a1a4057a0bbc73ec463;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfab554f356fe6780ff04c7a8bfeeccce125b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39bc59dfc15ba5c700827fa28ea0ecb7fe83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde77b279ba124124f4ae5647ac4796ea49e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b6760ced6a722c93caf8adbc2079e805e75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2db0feb2d84232d5b684aeb6c291da68d49d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had586e70d75538ea0dfb000a3ffeaa368e0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha803823523ff180221c631c547b674c9c8d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4429137014f4aa3916e96aa44bf1b6e74d35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6982425f54589df0124355ccf862a0655ee2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda83a5af4d58d6ed882a25e5a5aa00244c8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h106534b9b13bde121decd545d73e9dd623e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ae32b6eb7ded2a6f329ab8003adac69a1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8401c0ee0ca70e8f09bb5f44d05cdd85b61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3aca22c633fe846badc146624e84b0758950;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd60ab2ba140dda5d7fc888295962619525c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ed39bf470188ef36789376d16793af4be95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88ee0602a5966dc9c34ed423a9561cee7b12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1847310bf8ff0ae750dd4e1c2d846e11868;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8613865fba0fb4325bd2751ca7a988ab040f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0df53d17faea85b33f30817a4e535808288;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7c393af17bb712e8d4b0bc3d63d64cd205f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10a62ea5308dd04d1aa661da95d9aa302288;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b9d4da5c4d5386c6523a2bbbbe3e952fa5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b8d4cd418f514b4eb254404d058bdc5ba95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce2ec8ad585273bbbaae3efbc993bbe5c964;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf49cd152099101ceb9966006f94148fc3182;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4dc9e5140d1500d455e7c4d2a0a5588202cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h540d4f684479b4613a9eaecc2c802286d472;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h542d28d1df66bc5cdcc67426dfb6a2c1038d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb786669765fe1bd76e105b8548c1e80fef69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77e5314be147cc10830f2bae088b91120e23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcef34b50692f4e86273f41df2c6c7683c0bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66771bb4e041775fbbf81a1c0f8a50f109f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f8437ceb51391643b3c8720797189d4f75d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bab1a169f6fa52ab3acd59c2fd88993b19b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1446def657045ef4193f5e2dc93db4551e26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3919fd0d260213b1fdfb8a5581e050174959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63232b1a60e2a862850a1a1e169faf6c44af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2c562d4fed2952f1ef85e42822cd0d638c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd293aa82e2f9ee52378f1c25480da6503da2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5963dfedbb64d8fb40893adaab4c5f0009d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76eecaa5333bde64fbd6a6e1faef419ba01c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50eefe462c0bd7c11fe2bd0d424a2e7d85fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa1db4d30a2ff6262ae7faa7beaebb64bdfe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd227f13554bebf062140040032d645563701;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h948b1f44befe854093ad0ef7f9f6ea17bbf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd28d0cc14f432b7d3776398a6ac78d89b98e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dcedc520e8a92d35db1257d76448ac5327f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37426175e6418976b04736c04408c690247;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d6c3829a2718fa1f9ea22c50481a0c80c65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e8a5f85ef44e29474a1df9b87283b271f0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7eb425b4173b065b37a16515292c7d2951b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37713e1a72914689ced08d9b19f91a2a7674;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc64b30bee30126fc789b54efbb2b82a93d02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b06dd23689e04817808289913fd15f67c7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d5f34d757b5762adcce41b75a3ba09aed86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h990ccb3b80a2b0ac4c0cc1e443daa2f1fb3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0cd1992bec2f51d9a7a44764fd5d8098d98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e50420d8fb23f95874cbc6d06f5400e2b7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha92f7263ec93463414ba79f5c4d64097c975;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10e10e3d2662954b442f6e50c2b23380ff75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30ed9667e5c2450d68d89f29b91771905965;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb38778f69be31559b6bac13fab753aa750fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h297e4df03fe7a6bc01d8ffc0729c0eaef109;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16e914631b7a1ee34d1419a98e8d57262f0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8422e65e46023735a29bcfbea150350d7bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfc3ea02e837b5c92dee1f66dfb54b848cd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3ae141cc824e600fbca4fad4daf0b9cab87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea3b11fafd2663b7ba56a88fea79d98c87a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f35a6341c13286950ce3e261d7d2a5ffb30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d9ff22d8c58d77e78bf0b3b7e950975a08b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c31f710becb2346a061cbea5bd1474d871;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha44ce9c72d37c0aacf686df48541d6ce4d4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1349f2be2473dcefd064686f1b7753cf68bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdafeab3b4fc6fb79eea6df5efcabec48a497;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc46b15c1f3910a2520cc1bf00f5a551b5e6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46bd9405d79e035063f00230d5e191b900fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7256c0def1c32da10020b9a70b4bf92b63f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73094987bb7f8f7a53fee4541c7d22fbdeef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h719dc3a89c5935f19aabec4e067ae36c845b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fcbdc31bcc2c94882badb68187227424eb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf13c180bb03f4cf6c54cf3de394ec91e968a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64ce40b27488c69d1363965ee8ec2f56f59e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h881630ad5d218dd2071a05f202ca40f59049;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h840ddd0b2afd1783ffd751c012413040afb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbef9219203c5ed2f29c38e613ac1964763d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde50dcf0df86728339440b7eaf17c030c24b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e8bcc24a197626bd39075c39cbd20f13db6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d7b675e68e4e342b8ea366dcc93628f9beb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha01e6a0ef18f775746f740ca05c95d41e1ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97735027c5fcda0cf5475e05c26630399079;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha19221a1d74d6bb110c4ff480068c968299;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f81e99db0c482193b9a6008aa747e2e0c47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb3c39991386a0f072d6c7ca683d6727a7c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecd262554ba36789ba8e74aac141250ecc8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cd625948647f07a38b82cb9b1818b6527c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h180b68cc13d0836af57832206cdf1051e271;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45f6fc62813633be854d28a2a46aea6c053f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcab29f7408787c75e946fa28df64e3585358;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b737fa29fa349c4cdb6ed0e2e0ef1c864c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2080b31158a8427ead04731f2d3aa4916ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d87db1d132dc8c4161fe13a23ae78311dbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefa81d5d98592138e350b41c2a893104baac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6cf056d0c68d3bec66a88459b330f9fc39a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6edf5035205980f6f322a9eac2794ec7ea65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd039855b249f89b464df5e3b2ba33f4b7360;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4610a9b4be75f23df08f7fcb103c7d8422ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d2245384c8ab38cb1674633d0e3c18e940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h296d44850c933c43fd3d3e715da9fff71662;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7af0a09716d3cae98881f987a129ccb1c2be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84f3da36720861930944273d04ddd5e4ec50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a45f9873bf995b7f9a8c4f0054ce49e1820;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e9f7858b16ba12338493ff737583cab9531;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ce031da092dbf70aebed6bf6acf38aec9c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h485d5b95dc8ba97bb0e4a1642c284e415408;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a2eeb231ab2e5af97e232658b68a8c7a03e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2413e6217851ea1636488bcc3773eccebfd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac5085ae6d091b358757691d9f97d7299a76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46a5c4cf931fb29282e375ac519e7b61dbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2d6f43ef57d27514253d76d1770373c9674;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h420987781a68bbc1986534fbc13185646f25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64b13aa54c46f0c0e622fdf47903d61d73be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dfc4622d46f7104e64918aea4a04bce164e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ba9799ca6acbae494fa152c6a261885d748;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c8c4b0614fb8f698effda5b48d23fb6c816;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafbe1607e0cafb0891395f8ef6bb4fd88aff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h993d03197e0e75523fb0d8c512268c290cde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98564062ad2f685dce725ffe58ff0b81521c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h760a72279dc0f7886352d68d125300ad8ac0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3339bd1c08abb2e125d3f8717f4004af8ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3158d88597207ea2b1e9e55e536a9c41b084;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5181e1237280b619fb7df0afd081716d4814;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39bf010d5e62c2e2159ef8d0e58262421c0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h360a6a4c5e9d8c928a4c534bd633f141a70e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b6dc7baa16ccfdad58eba10658c4ef5c8ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5170f6aabb2b08995482b4cac4f2681e9f7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb58b8bc9da8df016301e3f4f5782c8bc017;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0c6f78cf91e452261b7bd006cce93728ec9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd848647f3ef200e5fe2d67c68e2eb9fd330c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73264a6c0562aa4bc5b040d10f25f6a45618;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h313871523b0b6be394a74853511a8b5d5480;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h393ca20f4074b926b38cff12e09c51d2ebd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he614b8d3a372a220bfa5d86ed6a9a5b622a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2cc64992a9ae8a43c561d211b39dd9a91d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca41d1069c759bead4d837e896834ee48d87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bfa5382d570cfdfafc9a09ae9a5f232a57b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c500d613b0b642c0208e79a81117c1415b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cc161f129f51ec59c1947394e687877f792;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10e79ca9347be3a937cbd0522bd36692b490;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf0f81410f317ada65462fa1bca1821f59f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4860c8869469a4ecd3f7907e3393b46a4d80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bc84a24167dd98277303cb7208b01044fbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71888ff5be2a7e64f953e20c9c6cc11d155a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ea7c5ee3f6e3a55039799549fcdccb42a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3aa5b69f13d9e3ffb07cef50f7aa41828b8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4105a0d556baef2fec3f722aff7a44246725;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b76353a01b464c3a7632fafb938ff0ba082;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8cf607cb00d23a29836e6853fd6a4df98b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6788a78f56ab7a3ae0e00ca2b3aa05765d0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55c214d468716c6fe45e8502a2811256095;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f39aa873bfe9ba005f72a89cfbbe0e858d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9cf7698f5bc0b7af70086874a47ecce01ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4461bdb4fa78401fdf7ebc1c1cf3a0143a21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d6b96bae62fe2faf2391952f32762209773;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57b4b140ae710916fd01f9baa42c6fa56c11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb0a559844c47db4b92886faa40011aa0b2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef9909881c30878aab7ed5f535eb527812d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f2dfb04732b245180cdb94121f303bedb65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefb432bb0374bd48e19368af09534b20a78f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ebfa086260b9f61484103cdbf5f3bb322b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4daaacf8afc44ab9c9d3c0c07384ed076280;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e2cd07b27fcd63f0aee3b340520eaad1a6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57fbe956bd5ca5abb871b3a12b779a52a9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38c9846f91dbbf1bdedfe61ecf26d7ad5cdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e9a2e4208951169239b60570803a92f6a1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d9d873e7812b878e4a82f776a4a05673c9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e2539296159670b77ce0795f133d85658a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf394982f5b6fee558872278039fc3edcabb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7cfbbb548abaa418de20a52f53792a6e65d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53476139de5f9cbc3c034388c506aefaa377;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa7d2c4c6141bf53918a7bfa538c3dbf2952;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc062d919b31af4d813b19fd151ed0ba6481;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5aad1457f8e50a9c648f9453354956aadddf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee967bd9060778757c3874ec34ff8b279e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a7f99292c164440b315c04b3c53b64b47ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h900a06154418a97110c775e2208dc85cc74b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b5f4d920a3f96e9a31e23cc43704f8e9270;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd534aa44a050fc9dbf59be134a1bc3d94d2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4cb94fb46f135b8b7565252da6661c174cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d06f1d15b206593d795285ccc4f7e5d4cce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39d2d91b1ffa29143eeb382bbb702d8072b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b8d11c018ee29bd14ed54928a837657d350;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23011109a1652d84137814df3728ab9095d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8827b2d46759268d05d9cfb749a2a987e24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haffd3ec2f3458158ba3a9cbb04067335ad15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he16366d977384a64b2a2542daf11ea1c7594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbaf527a75828a2ade3ee518c6dbfda1b5fbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e04cbf40f2cb0628e2e0270fbaf4449650c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h124111552d1746cd63352941c51e4457ea09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74867cb1bae7987d1068c1913dbb94b7689;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he000acce93d26614357eda2e59f299e65f79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74db3fefe05ff11626e119d693f3482e185d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca56a71091af8dac7149595078eff6ed85b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33371a8fc2331ca6487970426c25e61fdfc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bbb5ef064ec25fd9d050657b3e43bcd1f52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haae55ce8e6dcce707695dda62666684125f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h439620538106e5ab47b68a4584323db4285;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a95fc730f3868de31e3b02199c657de3bee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f44f393a60fdaabcc9c62bcc499ca4a43f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6e068770c29b03c65258c21f41874413aa5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h218441e20a8ddadc9e0c27794785a883aae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf21cbce73530b1cc3fb0cac6780643bcd334;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a67f481fdc6cbcfacbeb9ae7d90cdfc6a5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1f1fbc92fe0802557fa5f7d23e0294dd044;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8dbd146525d78d1812095446a360525dfa9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcedcaa90b297793beb18adcee4a3551943;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0ac2aee680e5e1a0c3145a9b521f3bf06f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1972b1ba3243cd362cf5bca7d51b5fa0817;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4ee2e7703cfe2a31cc6195ddc4a2a98180;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72b8a006d59166fcc3f546f50fc5154ab9df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf328e4a9431eb0e82230a03ab060eb9cec4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50095a1e943934afe9547d42b5a7db6f79fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff4f76c4af471ad22e45da3a4c3d81b528a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha88152f10988c51968299b1e53ca091456bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he614ab904dccf1d6d6d6c38e7edde6722cec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5d1b4c6ebbdde5b0823490167bc0eabddff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51ac0ca6c247602b0529c62a8f9e5089998;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd70def88c1e4ea8b25fcc393bd7321f8e7f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12a69f5fb43bb83df6b8b66454bfd552038c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6be721e3edcd936045ac0f840e2185657c2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dac1712e35a2bc84eccee0805218362d19f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49f2357bdefb8de381b242c5e911b8915b90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb74a6f554db782060062980e1e99a04a6abd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d0c4e9d0a8fa76949bdbcc5f7cd84361e05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1078958db7a0c72c72598413fd03345cb5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf78329a754e748a095fc39d172fffb94c7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aa6fd08bb520716f83d6a12ebbaa00234c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7221cf8d82e846daef701b15005d71d3fb3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6912b62b426757ffd77f0c963551eee1197b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h545dc9e8a2659fe5463ad7893daf5d466813;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3e221cb79787861c621a68fe5d682e74ff0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3fbdac250afaf2e75a0717e69d8e9bbaa94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda73358c5de129686e38a3df4f1c23ccba42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4328f966216bef282cf1412a353aef420430;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde126c9d11d3ce736b17318861a23bcbaded;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc570e694859c62b32cada3c9ab601e298d11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0762bd6bfd8c63908d9c484ec382d67cfb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fa5f72407a6cd4607adf9440184e93f8066;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2122d9bdce96e7e90ba6885278ecff0b862f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee3dd306a2fb53e125dc4880fa7ca17f35bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb592545ba50bdfecbb0d9c3e3dd418fde80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb994c09e712a18acf8aba9b37c2b273d3e65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h246a33768154a8d9251a700e58c6b75b6000;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1ef8d8f9f2bfc0463fd56bfb1a06737c3f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb8b843dc7cb8abba754b692be1944109fcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfbe01ea4a3d5c92a039d3f803c1759d9a9a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8cf8735943b001f5f726c7b780637fd7b65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd09b1ed9916e6ef460bf4abb175eab9243be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83964546795594a616e90879bd493923ad45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadc76d22814c727af3840bc8bd866bad5503;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf037cf44f0fd07d4c6aaa61afd094ff66f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haeb736833f8da5bb438aeaaf8cef7e7c49b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63c8bb5df2ab681b3e3c92eae5c15c724668;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b5782f4c6497123e828e0d6b35a7da643a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dba90c32cb87a46933772d82f494ae03c83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f4ac07d028f3114d2125a4c5fa422ef4eff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7da4d8f004c904212a6a0fd3513bb5eb5297;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2337606c0ec001bb0dc0f10f4db49fa29c5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4489e62bb6930e39997a2d7eaa8813e9915;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9501545cc1b3b30e3a42bc6c0353ef044b2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8319d130be81fa0c17cc059de51bc3ec488;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5be3d265358e0ec53734f05583ec57a32150;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e78e55e8c9a959eef480d97364cdb187b23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h968cabcee6da37e9dbc27efa5e3ff5ce1f2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25e62a5c2b0bc72fc1cce8e45ce3f50f441d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dd42f2dc499ca4191deb9104b8c9cb69f05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee14bd14778af565173c3502cac52490f1d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h779bb772848ef7c94394fd3d56c81f6563bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f0e3099cf1d4a14242bc00b71c66ce0b6d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3639c215b69b4eec2817f66be1a80aed325d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55c6b9108c70f8ea3b07e3e2dfa204883953;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c8a4b0a37f3523b11e45dc1e68704296069;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f2f60c7b814f90c301f707e550e99c0763a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5543ba5b379871a7c9c1d9bb48c775292497;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had3daecab61da159a96004f7c34d11db9eba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8eafc79f45851c6b693d5d616d83a4aa577a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5e6099857ebff7dad1d39566a7a11fb10a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cde698ccba3556774266d5d8fa5d1ca3ad8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3ee4122f21841b552a3716fd59c1d1b31d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75c28817aa3d13c6c87ed8ea1253bf404b23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha38abf65590b90ca2176a55b923f6d635a29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ae32a63ede8e753955244ab053ac46b59db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4809a3fda65c4eec8c3262eb5f90ed431fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h201a11db0e64caca8498234dc5c0a61b0e40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h763e09ec77df82e4a4087b29698db2baefc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a38ae75c6022814511607fb142f35cfa141;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68eb683d3a261dd203af252af6fb8f4b1807;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3031532b60b50973c76ffdb46d01677ee28c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d64aca3641bac89c0d3259192cdadecf020;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hceb7a015964123f4d10b935b911acf7639ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ac70e933e2519ce94a968501e90f486f904;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90d187470835b8a5661a7976c25b4b1143fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a5301a6498df37069b1e7afc57c06c5c180;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcea46e8566f6b1381d066fb82d5617956fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7241eb5374d05ca8170478a34b61b118ab31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3ed765ab66ef82cb58f25d9400c19fc3449;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28e6e4ff89bced811b684ea58b6abba9713a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5eebed7c16602f637ba38940211cb88a04a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5562c395cde6fe2dd82445014192b34bb6a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80850ff422fb9fdc093c06f919f0a7cd21da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf16c9acb84ddf5ded6bb27320d697ac37a9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f1ab876e6b7835ea2dee2aa76e5808f4ae7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e7c0fefbcfac5d6d6cf41a51eb7f2eddbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78f981c2744ad76fd183b2e07a2046912c35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h981fdd96b6a84a001bb303607c993477a75d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fc6ca115a245fb3144519279724a60b32ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha369ff71b4f509f4d3e3ef682afc61cd8fe7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f2f0fa16358aea4d6642d639a47a914aa45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h402447c5822f9940f1ce6106cff86bbd3039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88b44edfc3765aae3d41c6680a1184031bd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45e7108e6b2e291893ffb5b14d7b52199d13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f1e375b8772cf58439372b93a5307f71130;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he21589203a6821a65a15f2d13869de157251;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68d4d97e7bfb92dd5d53a16dc3e71af1e4f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf203a72abc8f900fd6a4d6e3ad3f4fb294e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dcf1c672552fb1a4d73a662fd0193d90d2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha985a3ca9c4334f18aee9b131a2379dae86a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccf80e3a259c89d67e8a7354bbff855276b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2d5602ad8a4bedf5a555a6c3be341a50f30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4255f625b862e1a6de13e3073ecb2c98d72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbf9ab8282d015be92c78a115a0c255d30eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha76aee7db8480a3ef311e9c43464011038bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ca43348d54fb421315656ce70a2a6a52b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f3b1bfd7de030202716a5b9eaf5d783bf61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35a71a594e30ab26149be6f091fa041df40e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4daed9ea34e4ef66afd1873316ecd7a12ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed1014c028705d86e06baf4991045cbeb888;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd140aa55a5ffb53bc4a58acd9bb663c585e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bd40e242aad063d83135ae58133fdf8e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2b9890331123a33eef1b24965c5d3f0c7f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e2a2135ad1b0e429626bbb0fca10e3f4d93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h650c60cc703806f0dc13aa673b53a482864d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c8c0e301ee2241766af121b7dd1515d0689;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5854cbab5393ce824e2c430f1e1d55b0217c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he79644ac708c31f1806262205934efa29fcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbeee6b3d40e917aefad4bc0e1e6c8db668f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdac88d3ef49124b12326a38e66d9b62d205;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a30cecbc3b209450d49890df37c70e2615f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc921b5c5934b21389a16effeba98d98e4b1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc785e2b8a3fab33c25443b9c182437cc6f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7b3d4c15857af4521b61ddc265005f45db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3cfa334a530c2c16309cc5028db095576d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1b0db2a66a5f0c2244e490d18f48cbc6eda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha63e138b38e3ad49470ab21741386e45c3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h133e0a9daf0571291587a2be55445befeb38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a5fba50de9c631fd9cbce335161a634fe74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89422fd308968b8b1b46eef4f8d227209cf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60f213388aba98010c2825d1d5d1ff5a054d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20eedfbd4077da2f6213f28b22df9392f6de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h802980358a5a4f77cf30ddd38a1341dc3332;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4530912c0447afa3119e523a84eba6f1413a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb7a289f9dd2111b014563f4b9a47e98d96f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6f507d172b02268211f9992cf917d3ad625;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc21e9c31c1b9abde6cd260f6f1ec71163675;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h934c0eb4d8e7aaf73570d9eaebce7052fdb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5082a8c1f8ce60e6d9e4bc8bc42f30824b65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36950322eddd95cc961aeaed114caffec4df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb32ce7eef34490a9edc76dcff41c33030cee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92ad3e75125b17dac739dcf9be7857ec535f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab5629974bf7aeed5d104c1c0a9e0a81fb3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h125fd31e00b168872eb8f7ce07106f9b5f77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2924005cbf4b26b9a5aa2708e4b6e26aa824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3d8fb6ad641100f71ecc4ee2ad168b5a5bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h220680e66f236c521dc787d775fc6ce1a455;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88da661b855885b3985275232480f682a34a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2737765759492a9330bcf847b263c8bff166;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4f3ebfddbea59863dcd73601d8f00804fc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb4c97ea23aad22f4b0185337e011c0159df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha57dd6f09e6732780a2a4442d0845afd3ca2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d6ea052d19d1c19ae4f63e38c1189210756;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95a70b0b0c76385a5c8e7cf1fda21982ca86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e876eca769e4108e637995f89fb0760dab8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heee5dae989fd85c41a80e885173fafcce89e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f4d64651f5618c75e2758a5864e772b3449;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h256cafbfb8e184d8cf9752eb77d3eb8d51d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h124fdd230574d59b101a4d3f34f4fe79874;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h608425d1125088778e117f335a8dbf2ec1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb26cb458ddcedf9f878aa4956ed9cfd5f40f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f4c7eb96dafd7c15b6192c31515462422e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff6add2050d0c0a0b1e87eb3fc75db266549;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b47ef942e7c4e580e33965b4d0d115d6c20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h865d30148761fe2bbb7826c30762786aa11b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e8c95996336c2ac7bfe4d563f9a34afe2ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h612dce1baf84e4bfeb33259e18876ab950d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70c4ddeebe4c0939054cdef69c8876ddd278;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87e093dd6e269e36ffddb305cadca4d1c8fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23674527cf187836746ebd653cb2e0094211;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf113eac42c29bde562c62a8a6bb72e249fce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d38e7314bb1787121f5d90074a6aa2f0a16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc90a678b743bbed4a6ef14a21bc130c7d01e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d92dc48f88420ee10ed29eea23ed99ae576;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h322de341cd7b759fede3286e451b96815291;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd543ca0dba776ee5ddb77dcd6e2bd46b523;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfece28267e8093c9a56e34396b75af25b3a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58a3ba8066590884d38f17a6899b2006e0f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc0f9aef6b230d35014f06bff62d394e298e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf449a59735cd088c7ef43b0481c474d7a4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h277dc8eb02fa8c92b674bc97724f74ffba8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8723c80bfe6a06f16a863ee571c5ea2de3fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h416ffe79b1f1d5207f209d9d81c99f86abc8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf447982041d68f89543acfbd7adbf74df17f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef45e1448f76ea0ca7f6ce0bb9774ded31eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf94e7241f933575efeda2521746934630d75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h350149084ccbb3354fb89b90b4b4e716cf3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5590226a4c90fe66b59cbc0f7a2c5f7238ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18e29c087ebc5e25d8e1e7f16a18079aa2fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83725cc6326a7113dab82de4789916bdc167;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6647747f11460334925938128e53a6a534a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95ec56d960f4578ffda732cf47bb153da564;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h314ae6357be29dea92a7b503e78f14d96ade;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4049aede11806674ed8a2a68bb5db52d94a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h560a8ec014758b2a9426bccfd1f820933c0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd9ceb5dfd8e75767da19d8da00a0f8f3138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f266fee1b521343d87fcdadd7defa3fead1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54a3943f266a4d9ff38eb1f94b9b370a4e1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c231755fa7e785853a383e397f43ffe9dc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59a9b4c32b54effa53611fefe11d44011c40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92cc0ad406cad00b6b7b77dde0f4e460f661;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2bc4d93fa8b0c0d0965474be440d4bb09fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1609140b330f2bd9393d33ce86eeba42915;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd61e3f9519179708ae5be135073bb4d02d0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69c6f1055699d5bdc304acf911cf0844b215;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60c5871f3f5c873f82e1d2011f7a5246ee73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b3485faccbb2fb5854998ffb129f61ca46d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45e43c2f5ae7e8f3967db9cfef772bea13eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3607202dcca333564a48eb9204e24e007d08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6129d95b1d802e8e16f0d5b3413686a67deb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe2630dc8c900ad16b61852c61d039129fa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3af1cdc3fbf00c3bc8ac7c7c8a31cbe72030;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78f3435b2479361dd12cd99093dc4787bf9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bdff9e9d312c390a26a0537281f0396e93a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde6e9d0c317c9bb57c6b5b6ede56596ec850;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34d4a173f8d6b96a380a72b8204d7a263999;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3582a35865af5858ef053e0eaa84805c50c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3af89d4ae1b8a96a6e9d2815d680a182276d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h581efd436dd7887857fcf18a64fa5d4a17b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5724e08e6e8c0a08a0ba8a08ae2d3d541d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40451a4840cfd3789869b6f9bd6abbe2e985;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h343c8855cbdcd4633523d1cc46a67dd07a95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59e80d1dd14ce39091cf9f1c3f15b42ef7cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea7db4df8fc7f466e03cc26fa7b598f584bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd613bf03b0e39934d68ad3954ce14958c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e3c77aa7dca11fd345a5eabc44aa7f8d9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd43a8533505834f7edf02704e7489e0c2765;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6dd4bf5905a19a3f10e8ef2fa74bb4223d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0899809e9e753abb061ed55f2b5fd74a4cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8fcda787ee5c49f57b7a0525f18b0072bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7371b36a4420d598f73b65ec50770559866;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8593d17ceb735081e2d717a5ed58a4a14060;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h190c6aa3847b7a97cac69cf9df1fbba8979c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87aeab25a6fa1648b68f68af80fdce3dc4d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17bb2e7dbb04af70fa2b14e9fe157b0b681f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h329056cd2bcf77f930fb5a6101dbf689c082;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e440a1cafc4e070c735ace1d4f737992a98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd25d71cf15529633498f42744b5327cdb6a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a0fed765b68d5db36366b3953a25add3551;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd2a8b55a08ee143e7216264f6591d92c0b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec322a5fcdb8f8ee3a8a2a5aa3da4108d12d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aeb1f810585ce330498e41a73ffa16c0fba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50060b5f0501085de4d1e1981da891fe97a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd7ee4b9726f0e0d17c7f7169d0e1ff15c11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f3206aad806d89e2943fe1af164e97bed4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc123ee0897718525ba3c5e3b4efe99aac948;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9374d437b3ea742ba308ed65048d9693f48b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b7d86975d0d1201cf7a7faecd5dd8b50039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b7ac953277465ed82cb559fafe64530ed53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55237ce21cf2fb61b769bb4eca1a716e27d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e3d3e94f78cd94201c1d02e27ee5f6bbdd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3e353c9d0e4d49a95b0a98d78b4e9dda370;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5009877db805bff6d568bc8738b846318f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cf8afd4eed89d5968ca1a42c0b25fce8c99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h910c7614e7c731c5624cf362c04e929fcbe0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h977fad76be0e48db0ec521317ba6a37488ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d9d38fb517ca6f39859d1e3a4b1e18c9a2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec55e01646ecaa7f29687c38e72698ad6992;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc781592baa7a146b580f63b7341a84b6f65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b7a725592fdb2b6d084fc6dda91a06678eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44368dabb1fbeeff1eeb0d9fa43c9e62be2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he85ac547fe0f72deef778d6f071d988a6ac6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2158dfa947f375a7df3414ded08080caef10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf361f5135e2ddd4bcbe0a1f8d0af9a8d7e62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e00334a986ccc6973533355b7c30e9eed66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc060f1ee20456ee071aefd95cca6178bd4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6031114270cc114fb8b4e57f5594625951;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcae93b279a09389050fb4e18c6055f894856;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he89636eb21d77b3f14fd1007544f59350b32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2710c3ee1e81ab637ed0aa1e8b72deff6461;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21c765682ed453fb65d256b3e5faae4e0e9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99d4cb741a9e03f44a9bfe4af400da21069e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7a974b80cd73b0a1c716ea581d61adcbb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha242749d0dc15758540448be0d0a9450c39f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h272cf01c5baffa8ffd6e5be32f7e06c71d19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha161ff2cf196c0ee4b5e605469314229ef61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d026f9953b60fcf711d78571396e12a7b83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97a53a289f24ae581b421e19372c71157987;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he16d60a60b86655bd8bc471275b21bfbd4ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd426359df92bf2e88ec24d39048a20a11e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8d34820c7d8781f74d7e22468c318321c26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7eff90f2a89728603225f616d46b118e8e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf049686d338bd83580005e80c3ca2bfb59b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb642c09f531aa9f8d8175ee01b97a1f694a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h436b62c9a7bfdf0f2302e3c4e61e9a583d8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e8fd82cf52bd9870e2e6c882e953b623fb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23c41fa7162392e0ac7562a377bca298544c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf0fefd20bc604d6e5247cf8b33a05204667;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea5f11bba8fbbd3e0d1cafc22fa4f15b698f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h330e77fdb8bcea7f2dbad4ea35029811522b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84c8c8d2539745fe3d4337c5cd477927daec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1542c327e8b84d6ee943fce4aec5cfedde9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h252fc9b99aaa92a9b2e5ef8299256c32f617;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1e95b590b6f53bc887f2ff6a370394ef22c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h527128d2f9bd51976579d44fa37a60694248;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71f25740696f15644581eeebb3c8e0bb12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20ab3644bbc57ee65714ef48b1aa4ee521d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c2aa73ff26182fb17e1ce9bca859e16a95e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef49a3c4abe4c6b63fd3e682a9dd3462873f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha565300bef21a88bd87f193a3701d97d0ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd792c2d156fe172ed2ad69bf5dc901634ce1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had532b006d7477f5a520ec26409eecce8c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc16130bf7a10bcf1d83a93155e4e08167ed7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53bc8d4cb43d1ca1f6d701782f31a5e2e186;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e98a93e5d49f232174ee0b6066b7681c712;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd07ba56d80ffe3d655cc25428ddaed55ed7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf1c8e8f6d1386d944dfeb6f9337c4a47fe0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h701b0debc41781ed645d8a1350878f141a57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff6e09442420f1a7aa43f1b2e60c21ef8db7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96ece91056672039ed5f7477449c0bdccfcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67e6a320226d96c9ccfac26b185a8711b896;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5dc6c8baf96ff670b3d2a497f4f36203e965;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3acb3d6191c891a302a0881b4fd63d58845;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he96167c0cc73abe7f545b172b4b8e16d5a83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c6e046ac266b694920ab3af005e4cc66515;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14a55d18feefc7c89988d35852fdb28dc28c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30859b6ce12daced099ba135d741af45c4d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d7444dfbc5becf3e251cd33e02aa77afb02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb948cd089bf247a3f64c2c3e53213d008494;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdac582625c42ab0f78035fbf3f77865e0705;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20b61172243406f68993a9e448247c5060cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b9a0b5442cba0a76588b446b986c157f38c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88be2db67d85fbab378d3d3001c0bbc9ea51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3eb00cefec4ea9e2c100bc329a1c3cb65f4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd316773fd5d00c56f4b6bfe77a5ddeb1aa86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2194090a436aba5d010a880a10e51673dbc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h613fbef4ff4772391b2a5b122ac86427b85f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h264b64281f055ee5b6b88d7cc0decc2da8b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb03a999b0ef7de04013e54b3786e95eb6d86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d7aa33e9d84b39d8da7fddd90882af35e9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h199eeb689011ccf4a6e6996b73cc5c5e3105;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f002f1d37d6fa211cbae7fb0c6c50aa04d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99c73c86d3cf1523197fa848bd60e12f6d85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67261c956679f2c0a2ee566744e31ba48c96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4c9097c184f926287a55c34c91fafc8e0d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9d0b2b7ad8f3dffebd8a0fb7f1dd050ef07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5dadb1066f9cc9751102a6191bc1f110b16c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9192f2ceb3170c8cce8d6a084969cbb207f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf815924ce7b4f74dafc76a2fa34371a935b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81ef5c42a69d18c0b91f7f835e9c3a92454e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2504b78b16a4ab382343aad8de8b5c43971;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf3b4601d3bec5687c874bf96eccf1e579ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11af3a42f934919290dd81d942b63db1862c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cbe2e36e995e36bffa54d7577033e6a8215;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb10935c9eb776f72b167612a17b5c68e7c7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17f46a1612fc8c13024803aceaacfe4ddb71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffc1f674c1d741f4258ccbe310512cc528ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7126556e72b8e9292523b6202e1635dc21b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h133659cd8c1b20703f7f8778f3a540cd0753;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ccf5a5dad8d7fe61eeaf90c07ac55ac26ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf941e33dd6524533013f330c36602d6a2bef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h438f05536777de4fc75fb3317c1574ae8749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbd5f80aba9185b4e3d0ebcdda6010d12dab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h211b0d7227c2f31914c325d06c3cbfca304b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbdb9e0a1ecbca58f49447b9e0a2ed84b022;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb07b971ad29b2b7b6f2c458ce76fc00537da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2746d490a0c0b767b9f122bdf072e226f58c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b0982123112eca805593318a622c3d521f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he686d6ac937d96f6da7a7fcdef42e178bbc8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfbf414af539e9787ff5296745ffd6a2b09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2af8d507d5935d0cf0cdb479bc92c16841b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h492eecbe82354c98e0cdcb466d2bd94c3d7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habeca1eca69fedc0cd6e8e99b45c5fcb3d69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h553d0b9f00cff8d0bd01a6cc78cb5dab2edb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7766714a0b2184862a60ae9b2912bcec068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86e50ad60f1021bb9247feeff76d6b7bf1f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf69083546b9f1e6d5250068dee1939f5dbe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf8ab7f7dd0263402ab2a27ace3b0dfeada1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94b53e13d83b06db5b8c706671d591549094;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfd4d16a8f10b1e5ea3cdd61c715427924af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec6dbed9476b6f30baff462fa00db04ac4b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf5b67b0bbc0ac212d7687c41bc85b224e26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b92b5dbec62859738eae76c65faf23d0dcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he26b358e3b40408252d42111ce155ac88d20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafe006e6a1df5b21c2d30a4fc21412c18eee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f41e2548f1768782547878f2e837fdea6fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29edd509c92303676cb5342dd1a7d55c8f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9d56d444bd8657e9766ff3b17d8ed73764f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfed84ed98dd06bafe340596213aaa3d7d86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5751d5c2702281a2f2bdf3d3c33809091b7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb2c09881f0267f759fc9735352bdc628313;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b4ade52f7cff4eeb67d052f950be99c8a7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c49eb5aebd9e090d8741df33af7a2d2751a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7e123eb15231577880a7577e77f71ecffa2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d16cd53b7a7150adeac0f6e1e6693b1381f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec25fb4cdda4854da95234d1d36fbbd00560;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heebf39283d31deacd434b9c3958ce67866b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdde12dac574f5c18f4768b64a5504da9fb4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafa35ba0df76293b1c194796b277659babda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63701b5014b9e22931ced459ba0a8f90c151;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1d141199e9a5d2a7c07af6da620c7630877;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91c7bfc58b4397e166fb921c9f73257ce636;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff9f6a108465c341378fc54cb9a30a31d487;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c57e88ba62ef1ba92dca47b4efe98356b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf54fa56628176677f994b71627c5e2ca1ae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde7159c8c4b535520fbb420c4602f121f9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h691be912abe0972317b9964b0c45ffdc4f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40132ed99aea3d294ccae41d745b69291bea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58c193ee00ea0e440f8e51ef4006337882fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc02276c9c3ae0af40543a4d81be8dae0ff95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73ba4e6aced05f1aa7cab8d2b8a507181d63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd74d396c504c60ab324a458572ff3d60612f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde42ea6ecdffbe68306a486daa5b9c192fbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf040bda0047666cebe01a1e0f6da5d66d37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef478c7e0682075ab03bbcfcba49254475c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bc384ba4ae08bf50a62dbd4869bf745cf5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h277ea81df27c98c7f1ddf22dcf93e6893e93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69816aa0403b44dbfa88a96ee95cbb7b0dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2d62deb44a0d9f9e5171375e88b49f63577;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2068fb801ed095bd1dea369e066ab34a1178;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf17e253c79223c81fca6144c7e10951b550f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddd1a1a5cb2aeb5f31cf1d870afbcbdbeb56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d35a89bda4e1d2c9be831c4495a5264362e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he50a04967c1c68379016b6789d2d9dd0b488;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7600facca36b4c092268fdacbe66e4f8485;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7bbdc65dd2f584bcbff94ef6425dc175eb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h205c87e38d88620db1fb4d17934b6f9a1ed0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1d12016858ce2fd94958e862ea520d5ec30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f2c8011f0c65842910eafebe7c01474d639;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34fbca4bc7ab7acf45a55a95c13789f306b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bba29c50d936e07a3fbe8f94c5d7855d48a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3597790fa349c8b6a6d6eabc69f72bfbe58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e60cb897275cf08e9b83ded80cb6e25c3c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aac923d9d2f3cb0bfe4c436a7e58361feab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h963817fa847cd3529ec3f5e12ba05e4c8674;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d22688a373615137c97b9dc8b74388ff3bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6624eea3d6fc7bf6dc24b88027a5461c21d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4a4dc6ef31929c0c3b5eb2d4a942d1c277c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2abca74c1e54b1404a0f3a3654fbdf543a60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c6fcfdde34b497cc45d2b466bc0b7406b14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26ae2401fd32c33c6143393f751b2bb73284;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e432ee3c4e82c917e94a5f8d1b85a5cdeb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h214f9585983bd0b5c617dd42e5d94306d052;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f1778ceadc86fce92a5d963b53541663fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h203558fb8617cbe456855dd9abab10d659ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc880960dcf90592d4499b153b116f1d91478;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8646284e7d4cbcf36e28b6cc1309cbf69256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c5c01a6f5e8749dad077bb9116cd7d656f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc600489bff9b75ddd40f97bd19d14e73c5bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd92e675ba1699f835b3a5648021d400a7918;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c3cd60a2792454de74cb9901e1c7b5f0c11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e80f3b7accbc23e436ec06a57d6e597f13d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a98f2a1ba265385f99db8cd819a8eca9552;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31beb2bcbccd766268d0430d85cd465ef498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8350f8d2edd3b4d53ab58e87f466aa05cbcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41751a0a6ba50c5a5834cbb0228028fc2c89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92f3c536722e23a71613e589614aa5714812;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54c791d37cf2678caddc99fa40268b93c03c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33df6f21bf4628c42b04363dd88fbb36a0bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he796a4f0257979c0bb2eb2addafaf21bfd35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92841702defe6c1998179f21da7fbca941ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4dccab2a883db38f4112ef6b09f19691090;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51265a26152437d826c38b2f339f01f188d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f66c36f4ac4f5f83665c3c47cce55700a48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h546f05a524e591afead7ab44ef9a6a1ba4a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0ceb26f4525bc14f1462a8bd3c66bc9ec34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c4107c5538caed07f371d2457298e2e9ebe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ed9685f70135af737e0d6ba0a2d4518c71f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4c4a7e2a8bca56e6b3e006c117e08e25a39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4662723112343c7203e9c6cce3449ad8a216;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcfd39a282186f1cb8ebb42b7868f8e722ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53d44308f6e7b41a6e8c5d808c35007c1820;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d0496980fd54c79e94be78aa32c5493872;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62ee120fc2831ca3114cc80ad1d73704e17e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b3814f12f0ed666480f49d1f7ec45afc50a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h436b59ad667049c09fbe61c454dbbfb24a35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hced1b773b0e1a42f9e08d2aa176fde1e18f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67320f85ebc6bb28d1c487d7efba7f58021c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0d46c88d9a15b4d3cfa7a9e7e15f414ad12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72bfd9657f41cb424d5769cfb601cfabe106;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ce22a296b32e00f4fae6326113c86d1194a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa24fba2456b663b6e2c5980f37b555141f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcb08f7247b976c34d4a7d75eb917bdc732d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29b6a750f023c252563267aa1c4dbe08cf5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha19e4fdbf0de4cfaacee7c034fb6e034324;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f77d8e67d5e72ad36dba9f9ac2485434cb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3983f2e41afc7f886d93fa7e57ed61a63267;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc50aff98c6ca9685bebb4779b8cec8fb1448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd41f3837b84678e770b4139daa61de3e5c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9e43610327df4f2ed99e082727a0b1f6962;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h534782e792f176373f9a8a9f094a4b1d10ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ea4190c83ae82e59019122af55bfeeed713;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31bbdcc4fc2f6e3b9964da7e455864ca5144;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf12b87b251745d1be1a350e25b99422a26a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf063592fd46cf59887abb53b043544e826cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5db6f5566773ba124392ff04b4e6125dff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h247a14e24c2f5d9ab338d670a316897ad18f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2509b3bcf7e7c21ffeaffa3a98f3892da757;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16b7c6e1fbd56a07fae97d79a79f413bce87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3889a1cc161ab0968ab4471293f0ed8421fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c584ff0a423e43438232085f0ce0b845e75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h205510b5db04e443652cda7a896f2431a38e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5b4712a7a6624396d1ffabaaea5dadd8241;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d02a57d6dd51c9a69beebaa411080100866;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6378a525f15accc31db3c7639acfbe7119f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f84e7298768ef62866ae9d5b402bd515746;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4151e382648d1a4bf7feb71a57f9c819c13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1532eb71878a62472306734a1cb7fe0f389;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6217cfa6d13a7e3c6c3152813a441795722a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e27d6897b6d7e2fdb40628091a5aac89448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5fd85509aa357c3ca8861f50abca5856e2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ecbf6a5847e775b7015e03347513bcffeeb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2af96838a464272c977edc40ae806c84ce7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd2de5e7291591a3c3d2bacb55a11f8afd0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23797ef8c8aa4ad35d00f48cc75618b36cad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79dd2beef4321dd15e93e1b60929deae628d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7efda7a65c52699d005e5be9e3ee97cb7574;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5afe4bcce6dc1a0ddae8ba4155362475356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc09e6d935a8edfd9f39551cf895ef799589;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd94a59344ff5fa4802efc40b203f5b80b577;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe51f38cbdcf915039224fb3ba71e8d286d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50ed5d263ad64634314bbc090a030faf93f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b38acda5513c16ad3e8c2bf00d78fa6fb71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1d59d7996a35637cf47de293b20db5c75fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc59654b1307639118d2ea64d1f101c77f60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc26dc1b0100af295d8f7c0adff092d3f140a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb2273b519bef4a08fc006abd50b0e1b8ac8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h109afaf9692ca634753529965ecd77332430;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a118cdd192941861792263fc3e13b15f59c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b7c7d2102762ba7588768e6e355eed77781;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24a9a292f4adf0961638e40c7a74290011;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fd626ca9156703acc5c9f5c9efaa348a0ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedf0784c96e4886a1f1eca6e00eb02db21cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43f852769807f8426d8cc57e63b5be40276a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe8076990bf031ce634fd42177335ce93b38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57418d208589c94000b7b53d7160221ec858;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44ff994df497cdce3a24fe454e74faca6cb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc34943e306fca606c02bb8bb35052409972e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea8546c737859e439fc000ca29a09c6a407c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h308de133240884c16518e328e689896ca52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bd18edc4118aa90e9261fdc6aa14c0a2921;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h523386a5b28f2beb9da820aa28c98ec8d645;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h606c8ce22aad36315feaf9a1b5e5e9cafaca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e2b1dffe0c8bbe7db52774e64b3c323ff36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcb6a2f96684a089ae6e78982efea513b30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e33df3ce63574819467e798f77597c913de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5125364308667dfbf0353c07d355e8401c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6f9ed8de9f61381cb00d12f34308d12452b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4f504deebae0c1e026a227977897a8f28bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb47ef3c58a29822330a620acac4f89b20a4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba2a3a3f961fa6695e25efc65352d28f86e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5b3517fa81d27f3a734c5d749e77e002b2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdff38b0e7d727fded89bcd07606b39f09a5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66b4708d867cda2779348b09bef7cad64863;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfd3a3e3327dea558fae0b95034ec90f0d78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97135a103c0d950264aa18231d60ee6c658e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha20fdf29a02c94b942ee31777bbbc59766a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aef9586fec0b7868120cbb9933f70925cd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70af3b413ae0b06f69da975951c69c05c19f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44d9c8e372a00c79f2ea0937447fdc0783e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he661946406c4641dcd53296062f4ae9672b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h814f49c2a62f9dfddc11ad7fba536b18dc81;
        #1
        $finish();
    end
endmodule
