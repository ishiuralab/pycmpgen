module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    compressor_CLA256_32 compressor_CLA256_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
        src16 <= 256'h0;
        src17 <= 256'h0;
        src18 <= 256'h0;
        src19 <= 256'h0;
        src20 <= 256'h0;
        src21 <= 256'h0;
        src22 <= 256'h0;
        src23 <= 256'h0;
        src24 <= 256'h0;
        src25 <= 256'h0;
        src26 <= 256'h0;
        src27 <= 256'h0;
        src28 <= 256'h0;
        src29 <= 256'h0;
        src30 <= 256'h0;
        src31 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA256_32(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    input [255:0]src16,
    input [255:0]src17,
    input [255:0]src18,
    input [255:0]src19,
    input [255:0]src20,
    input [255:0]src21,
    input [255:0]src22,
    input [255:0]src23,
    input [255:0]src24,
    input [255:0]src25,
    input [255:0]src26,
    input [255:0]src27,
    input [255:0]src28,
    input [255:0]src29,
    input [255:0]src30,
    input [255:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [0:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [0:0] comp_out38;
    wire [0:0] comp_out39;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], 1'h0, comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      input wire [255:0] src16,
      input wire [255:0] src17,
      input wire [255:0] src18,
      input wire [255:0] src19,
      input wire [255:0] src20,
      input wire [255:0] src21,
      input wire [255:0] src22,
      input wire [255:0] src23,
      input wire [255:0] src24,
      input wire [255:0] src25,
      input wire [255:0] src26,
      input wire [255:0] src27,
      input wire [255:0] src28,
      input wire [255:0] src29,
      input wire [255:0] src30,
      input wire [255:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [0:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [0:0] dst38,
      output wire [0:0] dst39);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [255:0] stage0_16;
   wire [255:0] stage0_17;
   wire [255:0] stage0_18;
   wire [255:0] stage0_19;
   wire [255:0] stage0_20;
   wire [255:0] stage0_21;
   wire [255:0] stage0_22;
   wire [255:0] stage0_23;
   wire [255:0] stage0_24;
   wire [255:0] stage0_25;
   wire [255:0] stage0_26;
   wire [255:0] stage0_27;
   wire [255:0] stage0_28;
   wire [255:0] stage0_29;
   wire [255:0] stage0_30;
   wire [255:0] stage0_31;
   wire [49:0] stage1_0;
   wire [97:0] stage1_1;
   wire [91:0] stage1_2;
   wire [90:0] stage1_3;
   wire [148:0] stage1_4;
   wire [125:0] stage1_5;
   wire [95:0] stage1_6;
   wire [100:0] stage1_7;
   wire [119:0] stage1_8;
   wire [131:0] stage1_9;
   wire [96:0] stage1_10;
   wire [139:0] stage1_11;
   wire [197:0] stage1_12;
   wire [92:0] stage1_13;
   wire [113:0] stage1_14;
   wire [92:0] stage1_15;
   wire [95:0] stage1_16;
   wire [126:0] stage1_17;
   wire [150:0] stage1_18;
   wire [93:0] stage1_19;
   wire [115:0] stage1_20;
   wire [138:0] stage1_21;
   wire [93:0] stage1_22;
   wire [93:0] stage1_23;
   wire [253:0] stage1_24;
   wire [117:0] stage1_25;
   wire [236:0] stage1_26;
   wire [107:0] stage1_27;
   wire [101:0] stage1_28;
   wire [117:0] stage1_29;
   wire [96:0] stage1_30;
   wire [132:0] stage1_31;
   wire [73:0] stage1_32;
   wire [33:0] stage1_33;
   wire [23:0] stage2_0;
   wire [32:0] stage2_1;
   wire [34:0] stage2_2;
   wire [42:0] stage2_3;
   wire [73:0] stage2_4;
   wire [41:0] stage2_5;
   wire [52:0] stage2_6;
   wire [53:0] stage2_7;
   wire [55:0] stage2_8;
   wire [65:0] stage2_9;
   wire [48:0] stage2_10;
   wire [57:0] stage2_11;
   wire [74:0] stage2_12;
   wire [56:0] stage2_13;
   wire [89:0] stage2_14;
   wire [46:0] stage2_15;
   wire [40:0] stage2_16;
   wire [54:0] stage2_17;
   wire [90:0] stage2_18;
   wire [45:0] stage2_19;
   wire [125:0] stage2_20;
   wire [71:0] stage2_21;
   wire [46:0] stage2_22;
   wire [56:0] stage2_23;
   wire [63:0] stage2_24;
   wire [65:0] stage2_25;
   wire [67:0] stage2_26;
   wire [95:0] stage2_27;
   wire [71:0] stage2_28;
   wire [39:0] stage2_29;
   wire [44:0] stage2_30;
   wire [47:0] stage2_31;
   wire [43:0] stage2_32;
   wire [30:0] stage2_33;
   wire [16:0] stage2_34;
   wire [5:0] stage2_35;
   wire [5:0] stage3_0;
   wire [27:0] stage3_1;
   wire [24:0] stage3_2;
   wire [34:0] stage3_3;
   wire [35:0] stage3_4;
   wire [15:0] stage3_5;
   wire [19:0] stage3_6;
   wire [23:0] stage3_7;
   wire [26:0] stage3_8;
   wire [21:0] stage3_9;
   wire [18:0] stage3_10;
   wire [25:0] stage3_11;
   wire [31:0] stage3_12;
   wire [36:0] stage3_13;
   wire [25:0] stage3_14;
   wire [32:0] stage3_15;
   wire [26:0] stage3_16;
   wire [19:0] stage3_17;
   wire [37:0] stage3_18;
   wire [34:0] stage3_19;
   wire [36:0] stage3_20;
   wire [32:0] stage3_21;
   wire [34:0] stage3_22;
   wire [20:0] stage3_23;
   wire [23:0] stage3_24;
   wire [35:0] stage3_25;
   wire [23:0] stage3_26;
   wire [38:0] stage3_27;
   wire [44:0] stage3_28;
   wire [27:0] stage3_29;
   wire [17:0] stage3_30;
   wire [36:0] stage3_31;
   wire [19:0] stage3_32;
   wire [17:0] stage3_33;
   wire [9:0] stage3_34;
   wire [12:0] stage3_35;
   wire [2:0] stage3_36;
   wire [5:0] stage4_0;
   wire [12:0] stage4_1;
   wire [7:0] stage4_2;
   wire [11:0] stage4_3;
   wire [15:0] stage4_4;
   wire [11:0] stage4_5;
   wire [14:0] stage4_6;
   wire [14:0] stage4_7;
   wire [7:0] stage4_8;
   wire [9:0] stage4_9;
   wire [14:0] stage4_10;
   wire [10:0] stage4_11;
   wire [11:0] stage4_12;
   wire [20:0] stage4_13;
   wire [11:0] stage4_14;
   wire [16:0] stage4_15;
   wire [18:0] stage4_16;
   wire [7:0] stage4_17;
   wire [13:0] stage4_18;
   wire [13:0] stage4_19;
   wire [18:0] stage4_20;
   wire [11:0] stage4_21;
   wire [24:0] stage4_22;
   wire [10:0] stage4_23;
   wire [7:0] stage4_24;
   wire [11:0] stage4_25;
   wire [15:0] stage4_26;
   wire [16:0] stage4_27;
   wire [19:0] stage4_28;
   wire [23:0] stage4_29;
   wire [9:0] stage4_30;
   wire [16:0] stage4_31;
   wire [9:0] stage4_32;
   wire [8:0] stage4_33;
   wire [5:0] stage4_34;
   wire [11:0] stage4_35;
   wire [5:0] stage4_36;
   wire [0:0] stage4_37;
   wire [0:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [2:0] stage5_3;
   wire [8:0] stage5_4;
   wire [5:0] stage5_5;
   wire [6:0] stage5_6;
   wire [6:0] stage5_7;
   wire [6:0] stage5_8;
   wire [12:0] stage5_9;
   wire [5:0] stage5_10;
   wire [6:0] stage5_11;
   wire [3:0] stage5_12;
   wire [7:0] stage5_13;
   wire [6:0] stage5_14;
   wire [8:0] stage5_15;
   wire [5:0] stage5_16;
   wire [7:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [9:0] stage5_20;
   wire [5:0] stage5_21;
   wire [7:0] stage5_22;
   wire [6:0] stage5_23;
   wire [5:0] stage5_24;
   wire [2:0] stage5_25;
   wire [5:0] stage5_26;
   wire [7:0] stage5_27;
   wire [5:0] stage5_28;
   wire [6:0] stage5_29;
   wire [12:0] stage5_30;
   wire [5:0] stage5_31;
   wire [5:0] stage5_32;
   wire [5:0] stage5_33;
   wire [3:0] stage5_34;
   wire [7:0] stage5_35;
   wire [7:0] stage5_36;
   wire [1:0] stage5_37;
   wire [0:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [0:0] stage6_3;
   wire [3:0] stage6_4;
   wire [2:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [4:0] stage6_8;
   wire [3:0] stage6_9;
   wire [5:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [2:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [1:0] stage6_16;
   wire [2:0] stage6_17;
   wire [4:0] stage6_18;
   wire [1:0] stage6_19;
   wire [5:0] stage6_20;
   wire [2:0] stage6_21;
   wire [5:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [2:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [2:0] stage6_31;
   wire [2:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [2:0] stage6_35;
   wire [3:0] stage6_36;
   wire [3:0] stage6_37;
   wire [0:0] stage6_38;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [0:0] stage7_25;
   wire [1:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [0:0] stage7_38;
   wire [0:0] stage7_39;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc135_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc135_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1406_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[7]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[8]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[3],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[4],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[5],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[6],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[7],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[8],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[9],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[10],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[11],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[12],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[13],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[14],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[15],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[16],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[17],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[18],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[19],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[20],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[21],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[22],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[23],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[24],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[25],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[26],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[27],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[28],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[29],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[30],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[31],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[32],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[33],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[34],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[35],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[36],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[37],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[38],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[39],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[40],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[41],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[42],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[43],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[44],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[45],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[46],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[47],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[48],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[49],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[50],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[51],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[52],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[53],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[54],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[55],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[56],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[57],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[18],stage1_4[58],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[19],stage1_4[59],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[20],stage1_4[60],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[21],stage1_4[61],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[22],stage1_4[62],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[23],stage1_4[63],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[24],stage1_4[64],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[25],stage1_4[65],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[26],stage1_4[66],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[27],stage1_4[67],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[28],stage1_4[68],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[29],stage1_4[69],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[30],stage1_4[70],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[31],stage1_4[71],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[32],stage1_4[72],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[33],stage1_4[73],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[34],stage1_4[74],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[35],stage1_4[75],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[36],stage1_4[76],stage1_3[79],stage1_2[79]}
   );
   gpc606_5 gpc80 (
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[37],stage1_4[77],stage1_3[80],stage1_2[80]}
   );
   gpc623_5 gpc81 (
      {stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage0_3[219], stage0_3[220]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[38],stage1_4[78],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage0_4[18]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[39],stage1_4[79],stage1_3[82]}
   );
   gpc615_5 gpc83 (
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage0_4[19]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[40],stage1_4[80],stage1_3[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235]},
      {stage0_4[20]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[5],stage1_5[41],stage1_4[81],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage0_4[21]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[6],stage1_5[42],stage1_4[82],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245]},
      {stage0_4[22]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[7],stage1_5[43],stage1_4[83],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage0_4[23]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[8],stage1_5[44],stage1_4[84],stage1_3[87]}
   );
   gpc623_5 gpc88 (
      {stage0_3[251], stage0_3[252], stage0_3[253]},
      {stage0_4[24], stage0_4[25]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[9],stage1_5[45],stage1_4[85],stage1_3[88]}
   );
   gpc1163_5 gpc89 (
      {stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[7],stage1_6[10],stage1_5[46],stage1_4[86]}
   );
   gpc1163_5 gpc90 (
      {stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[1]},
      {stage0_7[1]},
      {stage1_8[1],stage1_7[8],stage1_6[11],stage1_5[47],stage1_4[87]}
   );
   gpc1163_5 gpc91 (
      {stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_6[2]},
      {stage0_7[2]},
      {stage1_8[2],stage1_7[9],stage1_6[12],stage1_5[48],stage1_4[88]}
   );
   gpc1163_5 gpc92 (
      {stage0_4[35], stage0_4[36], stage0_4[37]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_6[3]},
      {stage0_7[3]},
      {stage1_8[3],stage1_7[10],stage1_6[13],stage1_5[49],stage1_4[89]}
   );
   gpc1163_5 gpc93 (
      {stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_6[4]},
      {stage0_7[4]},
      {stage1_8[4],stage1_7[11],stage1_6[14],stage1_5[50],stage1_4[90]}
   );
   gpc1163_5 gpc94 (
      {stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_6[5]},
      {stage0_7[5]},
      {stage1_8[5],stage1_7[12],stage1_6[15],stage1_5[51],stage1_4[91]}
   );
   gpc606_5 gpc95 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[6],stage1_7[13],stage1_6[16],stage1_5[52],stage1_4[92]}
   );
   gpc606_5 gpc96 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[7],stage1_7[14],stage1_6[17],stage1_5[53],stage1_4[93]}
   );
   gpc606_5 gpc97 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[8],stage1_7[15],stage1_6[18],stage1_5[54],stage1_4[94]}
   );
   gpc606_5 gpc98 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[9],stage1_7[16],stage1_6[19],stage1_5[55],stage1_4[95]}
   );
   gpc606_5 gpc99 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[10],stage1_7[17],stage1_6[20],stage1_5[56],stage1_4[96]}
   );
   gpc606_5 gpc100 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[11],stage1_7[18],stage1_6[21],stage1_5[57],stage1_4[97]}
   );
   gpc606_5 gpc101 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[12],stage1_7[19],stage1_6[22],stage1_5[58],stage1_4[98]}
   );
   gpc606_5 gpc102 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[13],stage1_7[20],stage1_6[23],stage1_5[59],stage1_4[99]}
   );
   gpc606_5 gpc103 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[14],stage1_7[21],stage1_6[24],stage1_5[60],stage1_4[100]}
   );
   gpc606_5 gpc104 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[15],stage1_7[22],stage1_6[25],stage1_5[61],stage1_4[101]}
   );
   gpc606_5 gpc105 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[16],stage1_7[23],stage1_6[26],stage1_5[62],stage1_4[102]}
   );
   gpc606_5 gpc106 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[17],stage1_7[24],stage1_6[27],stage1_5[63],stage1_4[103]}
   );
   gpc606_5 gpc107 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[18],stage1_7[25],stage1_6[28],stage1_5[64],stage1_4[104]}
   );
   gpc606_5 gpc108 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[19],stage1_7[26],stage1_6[29],stage1_5[65],stage1_4[105]}
   );
   gpc606_5 gpc109 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[20],stage1_7[27],stage1_6[30],stage1_5[66],stage1_4[106]}
   );
   gpc606_5 gpc110 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[21],stage1_7[28],stage1_6[31],stage1_5[67],stage1_4[107]}
   );
   gpc606_5 gpc111 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[22],stage1_7[29],stage1_6[32],stage1_5[68],stage1_4[108]}
   );
   gpc606_5 gpc112 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[23],stage1_7[30],stage1_6[33],stage1_5[69],stage1_4[109]}
   );
   gpc606_5 gpc113 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[24],stage1_7[31],stage1_6[34],stage1_5[70],stage1_4[110]}
   );
   gpc606_5 gpc114 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[25],stage1_7[32],stage1_6[35],stage1_5[71],stage1_4[111]}
   );
   gpc606_5 gpc115 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[26],stage1_7[33],stage1_6[36],stage1_5[72],stage1_4[112]}
   );
   gpc606_5 gpc116 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[27],stage1_7[34],stage1_6[37],stage1_5[73],stage1_4[113]}
   );
   gpc606_5 gpc117 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[28],stage1_7[35],stage1_6[38],stage1_5[74],stage1_4[114]}
   );
   gpc606_5 gpc118 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[29],stage1_7[36],stage1_6[39],stage1_5[75],stage1_4[115]}
   );
   gpc606_5 gpc119 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[30],stage1_7[37],stage1_6[40],stage1_5[76],stage1_4[116]}
   );
   gpc606_5 gpc120 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[31],stage1_7[38],stage1_6[41],stage1_5[77],stage1_4[117]}
   );
   gpc606_5 gpc121 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[32],stage1_7[39],stage1_6[42],stage1_5[78],stage1_4[118]}
   );
   gpc606_5 gpc122 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[33],stage1_7[40],stage1_6[43],stage1_5[79],stage1_4[119]}
   );
   gpc606_5 gpc123 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[34],stage1_7[41],stage1_6[44],stage1_5[80],stage1_4[120]}
   );
   gpc606_5 gpc124 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[35],stage1_7[42],stage1_6[45],stage1_5[81],stage1_4[121]}
   );
   gpc606_5 gpc125 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[36],stage1_7[43],stage1_6[46],stage1_5[82],stage1_4[122]}
   );
   gpc606_5 gpc126 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[0],stage1_8[37],stage1_7[44],stage1_6[47],stage1_5[83]}
   );
   gpc606_5 gpc127 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[1],stage1_8[38],stage1_7[45],stage1_6[48],stage1_5[84]}
   );
   gpc606_5 gpc128 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[2],stage1_8[39],stage1_7[46],stage1_6[49],stage1_5[85]}
   );
   gpc606_5 gpc129 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[3],stage1_8[40],stage1_7[47],stage1_6[50],stage1_5[86]}
   );
   gpc606_5 gpc130 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[4],stage1_8[41],stage1_7[48],stage1_6[51],stage1_5[87]}
   );
   gpc606_5 gpc131 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[5],stage1_8[42],stage1_7[49],stage1_6[52],stage1_5[88]}
   );
   gpc606_5 gpc132 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[6],stage1_8[43],stage1_7[50],stage1_6[53],stage1_5[89]}
   );
   gpc606_5 gpc133 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[7],stage1_8[44],stage1_7[51],stage1_6[54],stage1_5[90]}
   );
   gpc606_5 gpc134 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[8],stage1_8[45],stage1_7[52],stage1_6[55],stage1_5[91]}
   );
   gpc606_5 gpc135 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[9],stage1_8[46],stage1_7[53],stage1_6[56],stage1_5[92]}
   );
   gpc606_5 gpc136 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[10],stage1_8[47],stage1_7[54],stage1_6[57],stage1_5[93]}
   );
   gpc606_5 gpc137 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[11],stage1_8[48],stage1_7[55],stage1_6[58],stage1_5[94]}
   );
   gpc606_5 gpc138 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[12],stage1_8[49],stage1_7[56],stage1_6[59],stage1_5[95]}
   );
   gpc606_5 gpc139 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[13],stage1_8[50],stage1_7[57],stage1_6[60],stage1_5[96]}
   );
   gpc606_5 gpc140 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[14],stage1_8[51],stage1_7[58],stage1_6[61],stage1_5[97]}
   );
   gpc606_5 gpc141 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[15],stage1_8[52],stage1_7[59],stage1_6[62],stage1_5[98]}
   );
   gpc606_5 gpc142 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[16],stage1_8[53],stage1_7[60],stage1_6[63],stage1_5[99]}
   );
   gpc606_5 gpc143 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[17],stage1_8[54],stage1_7[61],stage1_6[64],stage1_5[100]}
   );
   gpc606_5 gpc144 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[18],stage1_8[55],stage1_7[62],stage1_6[65],stage1_5[101]}
   );
   gpc606_5 gpc145 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[19],stage1_8[56],stage1_7[63],stage1_6[66],stage1_5[102]}
   );
   gpc606_5 gpc146 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[20],stage1_8[57],stage1_7[64],stage1_6[67],stage1_5[103]}
   );
   gpc606_5 gpc147 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[21],stage1_8[58],stage1_7[65],stage1_6[68],stage1_5[104]}
   );
   gpc606_5 gpc148 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[22],stage1_8[59],stage1_7[66],stage1_6[69],stage1_5[105]}
   );
   gpc606_5 gpc149 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[23],stage1_8[60],stage1_7[67],stage1_6[70],stage1_5[106]}
   );
   gpc606_5 gpc150 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[24],stage1_8[61],stage1_7[68],stage1_6[71],stage1_5[107]}
   );
   gpc606_5 gpc151 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[25],stage1_8[62],stage1_7[69],stage1_6[72],stage1_5[108]}
   );
   gpc606_5 gpc152 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[26],stage1_8[63],stage1_7[70],stage1_6[73],stage1_5[109]}
   );
   gpc606_5 gpc153 (
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[64],stage1_7[71],stage1_6[74]}
   );
   gpc606_5 gpc154 (
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[65],stage1_7[72],stage1_6[75]}
   );
   gpc606_5 gpc155 (
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[66],stage1_7[73],stage1_6[76]}
   );
   gpc606_5 gpc156 (
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[67],stage1_7[74],stage1_6[77]}
   );
   gpc606_5 gpc157 (
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[68],stage1_7[75],stage1_6[78]}
   );
   gpc606_5 gpc158 (
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[69],stage1_7[76],stage1_6[79]}
   );
   gpc615_5 gpc159 (
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232]},
      {stage0_7[168]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[33],stage1_8[70],stage1_7[77],stage1_6[80]}
   );
   gpc615_5 gpc160 (
      {stage0_6[233], stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237]},
      {stage0_7[169]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[34],stage1_8[71],stage1_7[78],stage1_6[81]}
   );
   gpc615_5 gpc161 (
      {stage0_6[238], stage0_6[239], stage0_6[240], stage0_6[241], stage0_6[242]},
      {stage0_7[170]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[35],stage1_8[72],stage1_7[79],stage1_6[82]}
   );
   gpc615_5 gpc162 (
      {stage0_7[171], stage0_7[172], stage0_7[173], stage0_7[174], stage0_7[175]},
      {stage0_8[54]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[9],stage1_9[36],stage1_8[73],stage1_7[80]}
   );
   gpc615_5 gpc163 (
      {stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179], stage0_7[180]},
      {stage0_8[55]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[10],stage1_9[37],stage1_8[74],stage1_7[81]}
   );
   gpc615_5 gpc164 (
      {stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage0_8[56]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[11],stage1_9[38],stage1_8[75],stage1_7[82]}
   );
   gpc615_5 gpc165 (
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190]},
      {stage0_8[57]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[12],stage1_9[39],stage1_8[76],stage1_7[83]}
   );
   gpc615_5 gpc166 (
      {stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_8[58]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[13],stage1_9[40],stage1_8[77],stage1_7[84]}
   );
   gpc615_5 gpc167 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[59]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[14],stage1_9[41],stage1_8[78],stage1_7[85]}
   );
   gpc615_5 gpc168 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[60]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[15],stage1_9[42],stage1_8[79],stage1_7[86]}
   );
   gpc615_5 gpc169 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[61]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[16],stage1_9[43],stage1_8[80],stage1_7[87]}
   );
   gpc615_5 gpc170 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[62]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[17],stage1_9[44],stage1_8[81],stage1_7[88]}
   );
   gpc615_5 gpc171 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[63]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[18],stage1_9[45],stage1_8[82],stage1_7[89]}
   );
   gpc615_5 gpc172 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[64]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[19],stage1_9[46],stage1_8[83],stage1_7[90]}
   );
   gpc615_5 gpc173 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[65]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[20],stage1_9[47],stage1_8[84],stage1_7[91]}
   );
   gpc615_5 gpc174 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[66]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[21],stage1_9[48],stage1_8[85],stage1_7[92]}
   );
   gpc615_5 gpc175 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[67]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[22],stage1_9[49],stage1_8[86],stage1_7[93]}
   );
   gpc615_5 gpc176 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[68]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[23],stage1_9[50],stage1_8[87],stage1_7[94]}
   );
   gpc615_5 gpc177 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[69]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[24],stage1_9[51],stage1_8[88],stage1_7[95]}
   );
   gpc606_5 gpc178 (
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[16],stage1_10[25],stage1_9[52],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[17],stage1_10[26],stage1_9[53],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[18],stage1_10[27],stage1_9[54],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[19],stage1_10[28],stage1_9[55],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[20],stage1_10[29],stage1_9[56],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[21],stage1_10[30],stage1_9[57],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[22],stage1_10[31],stage1_9[58],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[23],stage1_10[32],stage1_9[59],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[24],stage1_10[33],stage1_9[60],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[25],stage1_10[34],stage1_9[61],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[26],stage1_10[35],stage1_9[62],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[27],stage1_10[36],stage1_9[63],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[28],stage1_10[37],stage1_9[64],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[29],stage1_10[38],stage1_9[65],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[30],stage1_10[39],stage1_9[66],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[31],stage1_10[40],stage1_9[67],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[32],stage1_10[41],stage1_9[68],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[33],stage1_10[42],stage1_9[69],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[34],stage1_10[43],stage1_9[70],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[35],stage1_10[44],stage1_9[71],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[36],stage1_10[45],stage1_9[72],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[37],stage1_10[46],stage1_9[73],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[38],stage1_10[47],stage1_9[74],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[39],stage1_10[48],stage1_9[75],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[40],stage1_10[49],stage1_9[76],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[41],stage1_10[50],stage1_9[77],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[42],stage1_10[51],stage1_9[78],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[43],stage1_10[52],stage1_9[79],stage1_8[116]}
   );
   gpc606_5 gpc206 (
      {stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[44],stage1_10[53],stage1_9[80],stage1_8[117]}
   );
   gpc606_5 gpc207 (
      {stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[45],stage1_10[54],stage1_9[81],stage1_8[118]}
   );
   gpc606_5 gpc208 (
      {stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[46],stage1_10[55],stage1_9[82],stage1_8[119]}
   );
   gpc606_5 gpc209 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[31],stage1_11[47],stage1_10[56],stage1_9[83]}
   );
   gpc606_5 gpc210 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[32],stage1_11[48],stage1_10[57],stage1_9[84]}
   );
   gpc606_5 gpc211 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[33],stage1_11[49],stage1_10[58],stage1_9[85]}
   );
   gpc606_5 gpc212 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[34],stage1_11[50],stage1_10[59],stage1_9[86]}
   );
   gpc606_5 gpc213 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[35],stage1_11[51],stage1_10[60],stage1_9[87]}
   );
   gpc606_5 gpc214 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[36],stage1_11[52],stage1_10[61],stage1_9[88]}
   );
   gpc606_5 gpc215 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[37],stage1_11[53],stage1_10[62],stage1_9[89]}
   );
   gpc606_5 gpc216 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[38],stage1_11[54],stage1_10[63],stage1_9[90]}
   );
   gpc606_5 gpc217 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[39],stage1_11[55],stage1_10[64],stage1_9[91]}
   );
   gpc606_5 gpc218 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[40],stage1_11[56],stage1_10[65],stage1_9[92]}
   );
   gpc606_5 gpc219 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[41],stage1_11[57],stage1_10[66],stage1_9[93]}
   );
   gpc606_5 gpc220 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[42],stage1_11[58],stage1_10[67],stage1_9[94]}
   );
   gpc606_5 gpc221 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[43],stage1_11[59],stage1_10[68],stage1_9[95]}
   );
   gpc606_5 gpc222 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[44],stage1_11[60],stage1_10[69],stage1_9[96]}
   );
   gpc606_5 gpc223 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[45],stage1_11[61],stage1_10[70],stage1_9[97]}
   );
   gpc606_5 gpc224 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[46],stage1_11[62],stage1_10[71],stage1_9[98]}
   );
   gpc606_5 gpc225 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[47],stage1_11[63],stage1_10[72],stage1_9[99]}
   );
   gpc606_5 gpc226 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[48],stage1_11[64],stage1_10[73],stage1_9[100]}
   );
   gpc606_5 gpc227 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[49],stage1_11[65],stage1_10[74],stage1_9[101]}
   );
   gpc615_5 gpc228 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214]},
      {stage0_10[186]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[50],stage1_11[66],stage1_10[75],stage1_9[102]}
   );
   gpc615_5 gpc229 (
      {stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_10[187]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[51],stage1_11[67],stage1_10[76],stage1_9[103]}
   );
   gpc615_5 gpc230 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_10[188]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[52],stage1_11[68],stage1_10[77],stage1_9[104]}
   );
   gpc615_5 gpc231 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229]},
      {stage0_10[189]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[53],stage1_11[69],stage1_10[78],stage1_9[105]}
   );
   gpc615_5 gpc232 (
      {stage0_10[190], stage0_10[191], stage0_10[192], stage0_10[193], stage0_10[194]},
      {stage0_11[138]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[23],stage1_12[54],stage1_11[70],stage1_10[79]}
   );
   gpc615_5 gpc233 (
      {stage0_10[195], stage0_10[196], stage0_10[197], stage0_10[198], stage0_10[199]},
      {stage0_11[139]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[24],stage1_12[55],stage1_11[71],stage1_10[80]}
   );
   gpc615_5 gpc234 (
      {stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203], stage0_10[204]},
      {stage0_11[140]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[25],stage1_12[56],stage1_11[72],stage1_10[81]}
   );
   gpc615_5 gpc235 (
      {stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage0_11[141]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[26],stage1_12[57],stage1_11[73],stage1_10[82]}
   );
   gpc615_5 gpc236 (
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214]},
      {stage0_11[142]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[27],stage1_12[58],stage1_11[74],stage1_10[83]}
   );
   gpc615_5 gpc237 (
      {stage0_10[215], stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219]},
      {stage0_11[143]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[28],stage1_12[59],stage1_11[75],stage1_10[84]}
   );
   gpc615_5 gpc238 (
      {stage0_10[220], stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224]},
      {stage0_11[144]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[29],stage1_12[60],stage1_11[76],stage1_10[85]}
   );
   gpc615_5 gpc239 (
      {stage0_10[225], stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229]},
      {stage0_11[145]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[30],stage1_12[61],stage1_11[77],stage1_10[86]}
   );
   gpc615_5 gpc240 (
      {stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234]},
      {stage0_11[146]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[31],stage1_12[62],stage1_11[78],stage1_10[87]}
   );
   gpc615_5 gpc241 (
      {stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage0_11[147]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[32],stage1_12[63],stage1_11[79],stage1_10[88]}
   );
   gpc615_5 gpc242 (
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244]},
      {stage0_11[148]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[33],stage1_12[64],stage1_11[80],stage1_10[89]}
   );
   gpc615_5 gpc243 (
      {stage0_10[245], stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249]},
      {stage0_11[149]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[34],stage1_12[65],stage1_11[81],stage1_10[90]}
   );
   gpc615_5 gpc244 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[72]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[12],stage1_13[35],stage1_12[66],stage1_11[82]}
   );
   gpc615_5 gpc245 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[13],stage1_13[36],stage1_12[67],stage1_11[83]}
   );
   gpc615_5 gpc246 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[74]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[14],stage1_13[37],stage1_12[68],stage1_11[84]}
   );
   gpc615_5 gpc247 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[75]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[15],stage1_13[38],stage1_12[69],stage1_11[85]}
   );
   gpc615_5 gpc248 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[76]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[16],stage1_13[39],stage1_12[70],stage1_11[86]}
   );
   gpc615_5 gpc249 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[77]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[17],stage1_13[40],stage1_12[71],stage1_11[87]}
   );
   gpc615_5 gpc250 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[78]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[18],stage1_13[41],stage1_12[72],stage1_11[88]}
   );
   gpc615_5 gpc251 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[79]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[19],stage1_13[42],stage1_12[73],stage1_11[89]}
   );
   gpc615_5 gpc252 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[80]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[20],stage1_13[43],stage1_12[74],stage1_11[90]}
   );
   gpc615_5 gpc253 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[81]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[21],stage1_13[44],stage1_12[75],stage1_11[91]}
   );
   gpc615_5 gpc254 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[82]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[22],stage1_13[45],stage1_12[76],stage1_11[92]}
   );
   gpc615_5 gpc255 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[83]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[23],stage1_13[46],stage1_12[77],stage1_11[93]}
   );
   gpc117_4 gpc256 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90]},
      {stage0_13[72]},
      {stage0_14[0]},
      {stage1_15[12],stage1_14[24],stage1_13[47],stage1_12[78]}
   );
   gpc606_5 gpc257 (
      {stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96]},
      {stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6]},
      {stage1_16[0],stage1_15[13],stage1_14[25],stage1_13[48],stage1_12[79]}
   );
   gpc606_5 gpc258 (
      {stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102]},
      {stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage1_16[1],stage1_15[14],stage1_14[26],stage1_13[49],stage1_12[80]}
   );
   gpc615_5 gpc259 (
      {stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_13[73]},
      {stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18]},
      {stage1_16[2],stage1_15[15],stage1_14[27],stage1_13[50],stage1_12[81]}
   );
   gpc615_5 gpc260 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112]},
      {stage0_13[74]},
      {stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24]},
      {stage1_16[3],stage1_15[16],stage1_14[28],stage1_13[51],stage1_12[82]}
   );
   gpc615_5 gpc261 (
      {stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage0_13[75]},
      {stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30]},
      {stage1_16[4],stage1_15[17],stage1_14[29],stage1_13[52],stage1_12[83]}
   );
   gpc615_5 gpc262 (
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_13[76]},
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36]},
      {stage1_16[5],stage1_15[18],stage1_14[30],stage1_13[53],stage1_12[84]}
   );
   gpc615_5 gpc263 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_13[77]},
      {stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42]},
      {stage1_16[6],stage1_15[19],stage1_14[31],stage1_13[54],stage1_12[85]}
   );
   gpc615_5 gpc264 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132]},
      {stage0_13[78]},
      {stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48]},
      {stage1_16[7],stage1_15[20],stage1_14[32],stage1_13[55],stage1_12[86]}
   );
   gpc615_5 gpc265 (
      {stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_13[79]},
      {stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54]},
      {stage1_16[8],stage1_15[21],stage1_14[33],stage1_13[56],stage1_12[87]}
   );
   gpc615_5 gpc266 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142]},
      {stage0_13[80]},
      {stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage1_16[9],stage1_15[22],stage1_14[34],stage1_13[57],stage1_12[88]}
   );
   gpc615_5 gpc267 (
      {stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_13[81]},
      {stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66]},
      {stage1_16[10],stage1_15[23],stage1_14[35],stage1_13[58],stage1_12[89]}
   );
   gpc606_5 gpc268 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[11],stage1_15[24],stage1_14[36],stage1_13[59]}
   );
   gpc606_5 gpc269 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[12],stage1_15[25],stage1_14[37],stage1_13[60]}
   );
   gpc606_5 gpc270 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[13],stage1_15[26],stage1_14[38],stage1_13[61]}
   );
   gpc606_5 gpc271 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[14],stage1_15[27],stage1_14[39],stage1_13[62]}
   );
   gpc615_5 gpc272 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110]},
      {stage0_14[67]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[15],stage1_15[28],stage1_14[40],stage1_13[63]}
   );
   gpc615_5 gpc273 (
      {stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115]},
      {stage0_14[68]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[16],stage1_15[29],stage1_14[41],stage1_13[64]}
   );
   gpc615_5 gpc274 (
      {stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119], stage0_13[120]},
      {stage0_14[69]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[17],stage1_15[30],stage1_14[42],stage1_13[65]}
   );
   gpc615_5 gpc275 (
      {stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_14[70]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[18],stage1_15[31],stage1_14[43],stage1_13[66]}
   );
   gpc615_5 gpc276 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130]},
      {stage0_14[71]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[19],stage1_15[32],stage1_14[44],stage1_13[67]}
   );
   gpc615_5 gpc277 (
      {stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_14[72]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[20],stage1_15[33],stage1_14[45],stage1_13[68]}
   );
   gpc615_5 gpc278 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140]},
      {stage0_14[73]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[21],stage1_15[34],stage1_14[46],stage1_13[69]}
   );
   gpc615_5 gpc279 (
      {stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145]},
      {stage0_14[74]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[22],stage1_15[35],stage1_14[47],stage1_13[70]}
   );
   gpc615_5 gpc280 (
      {stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150]},
      {stage0_14[75]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[23],stage1_15[36],stage1_14[48],stage1_13[71]}
   );
   gpc615_5 gpc281 (
      {stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_14[76]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[24],stage1_15[37],stage1_14[49],stage1_13[72]}
   );
   gpc615_5 gpc282 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160]},
      {stage0_14[77]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[25],stage1_15[38],stage1_14[50],stage1_13[73]}
   );
   gpc615_5 gpc283 (
      {stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_14[78]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[26],stage1_15[39],stage1_14[51],stage1_13[74]}
   );
   gpc615_5 gpc284 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_14[79]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[27],stage1_15[40],stage1_14[52],stage1_13[75]}
   );
   gpc615_5 gpc285 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175]},
      {stage0_14[80]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[28],stage1_15[41],stage1_14[53],stage1_13[76]}
   );
   gpc615_5 gpc286 (
      {stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180]},
      {stage0_14[81]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[29],stage1_15[42],stage1_14[54],stage1_13[77]}
   );
   gpc615_5 gpc287 (
      {stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_14[82]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[30],stage1_15[43],stage1_14[55],stage1_13[78]}
   );
   gpc615_5 gpc288 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190]},
      {stage0_14[83]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[31],stage1_15[44],stage1_14[56],stage1_13[79]}
   );
   gpc615_5 gpc289 (
      {stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_14[84]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[32],stage1_15[45],stage1_14[57],stage1_13[80]}
   );
   gpc615_5 gpc290 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_14[85]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[33],stage1_15[46],stage1_14[58],stage1_13[81]}
   );
   gpc615_5 gpc291 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[86]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[34],stage1_15[47],stage1_14[59],stage1_13[82]}
   );
   gpc615_5 gpc292 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[87]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[35],stage1_15[48],stage1_14[60],stage1_13[83]}
   );
   gpc615_5 gpc293 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[88]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[36],stage1_15[49],stage1_14[61],stage1_13[84]}
   );
   gpc615_5 gpc294 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[89]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[37],stage1_15[50],stage1_14[62],stage1_13[85]}
   );
   gpc615_5 gpc295 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[90]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[38],stage1_15[51],stage1_14[63],stage1_13[86]}
   );
   gpc615_5 gpc296 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[91]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[39],stage1_15[52],stage1_14[64],stage1_13[87]}
   );
   gpc615_5 gpc297 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[92]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[40],stage1_15[53],stage1_14[65],stage1_13[88]}
   );
   gpc615_5 gpc298 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[93]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[41],stage1_15[54],stage1_14[66],stage1_13[89]}
   );
   gpc615_5 gpc299 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[94]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[42],stage1_15[55],stage1_14[67],stage1_13[90]}
   );
   gpc615_5 gpc300 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[95]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[43],stage1_15[56],stage1_14[68],stage1_13[91]}
   );
   gpc615_5 gpc301 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[96]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[44],stage1_15[57],stage1_14[69],stage1_13[92]}
   );
   gpc606_5 gpc302 (
      {stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[34],stage1_16[45],stage1_15[58],stage1_14[70]}
   );
   gpc606_5 gpc303 (
      {stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[35],stage1_16[46],stage1_15[59],stage1_14[71]}
   );
   gpc606_5 gpc304 (
      {stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[36],stage1_16[47],stage1_15[60],stage1_14[72]}
   );
   gpc606_5 gpc305 (
      {stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[37],stage1_16[48],stage1_15[61],stage1_14[73]}
   );
   gpc606_5 gpc306 (
      {stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[38],stage1_16[49],stage1_15[62],stage1_14[74]}
   );
   gpc606_5 gpc307 (
      {stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[39],stage1_16[50],stage1_15[63],stage1_14[75]}
   );
   gpc606_5 gpc308 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[40],stage1_16[51],stage1_15[64],stage1_14[76]}
   );
   gpc606_5 gpc309 (
      {stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[41],stage1_16[52],stage1_15[65],stage1_14[77]}
   );
   gpc606_5 gpc310 (
      {stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[42],stage1_16[53],stage1_15[66],stage1_14[78]}
   );
   gpc606_5 gpc311 (
      {stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[43],stage1_16[54],stage1_15[67],stage1_14[79]}
   );
   gpc606_5 gpc312 (
      {stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[44],stage1_16[55],stage1_15[68],stage1_14[80]}
   );
   gpc606_5 gpc313 (
      {stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[45],stage1_16[56],stage1_15[69],stage1_14[81]}
   );
   gpc606_5 gpc314 (
      {stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[46],stage1_16[57],stage1_15[70],stage1_14[82]}
   );
   gpc606_5 gpc315 (
      {stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[47],stage1_16[58],stage1_15[71],stage1_14[83]}
   );
   gpc606_5 gpc316 (
      {stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[48],stage1_16[59],stage1_15[72],stage1_14[84]}
   );
   gpc606_5 gpc317 (
      {stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[49],stage1_16[60],stage1_15[73],stage1_14[85]}
   );
   gpc606_5 gpc318 (
      {stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[50],stage1_16[61],stage1_15[74],stage1_14[86]}
   );
   gpc606_5 gpc319 (
      {stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[51],stage1_16[62],stage1_15[75],stage1_14[87]}
   );
   gpc606_5 gpc320 (
      {stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[52],stage1_16[63],stage1_15[76],stage1_14[88]}
   );
   gpc606_5 gpc321 (
      {stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[53],stage1_16[64],stage1_15[77],stage1_14[89]}
   );
   gpc606_5 gpc322 (
      {stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[54],stage1_16[65],stage1_15[78],stage1_14[90]}
   );
   gpc606_5 gpc323 (
      {stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[55],stage1_16[66],stage1_15[79],stage1_14[91]}
   );
   gpc606_5 gpc324 (
      {stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[56],stage1_16[67],stage1_15[80],stage1_14[92]}
   );
   gpc615_5 gpc325 (
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208]},
      {stage0_16[138]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[23],stage1_17[57],stage1_16[68],stage1_15[81]}
   );
   gpc615_5 gpc326 (
      {stage0_15[209], stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213]},
      {stage0_16[139]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[24],stage1_17[58],stage1_16[69],stage1_15[82]}
   );
   gpc615_5 gpc327 (
      {stage0_15[214], stage0_15[215], stage0_15[216], stage0_15[217], stage0_15[218]},
      {stage0_16[140]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[25],stage1_17[59],stage1_16[70],stage1_15[83]}
   );
   gpc615_5 gpc328 (
      {stage0_15[219], stage0_15[220], stage0_15[221], stage0_15[222], stage0_15[223]},
      {stage0_16[141]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[26],stage1_17[60],stage1_16[71],stage1_15[84]}
   );
   gpc615_5 gpc329 (
      {stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227], stage0_15[228]},
      {stage0_16[142]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[27],stage1_17[61],stage1_16[72],stage1_15[85]}
   );
   gpc615_5 gpc330 (
      {stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage0_16[143]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[28],stage1_17[62],stage1_16[73],stage1_15[86]}
   );
   gpc615_5 gpc331 (
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238]},
      {stage0_16[144]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[29],stage1_17[63],stage1_16[74],stage1_15[87]}
   );
   gpc615_5 gpc332 (
      {stage0_15[239], stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243]},
      {stage0_16[145]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[30],stage1_17[64],stage1_16[75],stage1_15[88]}
   );
   gpc615_5 gpc333 (
      {stage0_15[244], stage0_15[245], stage0_15[246], stage0_15[247], stage0_15[248]},
      {stage0_16[146]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[31],stage1_17[65],stage1_16[76],stage1_15[89]}
   );
   gpc615_5 gpc334 (
      {stage0_15[249], stage0_15[250], stage0_15[251], stage0_15[252], stage0_15[253]},
      {stage0_16[147]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[32],stage1_17[66],stage1_16[77],stage1_15[90]}
   );
   gpc606_5 gpc335 (
      {stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[10],stage1_18[33],stage1_17[67],stage1_16[78]}
   );
   gpc606_5 gpc336 (
      {stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158], stage0_16[159]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[11],stage1_18[34],stage1_17[68],stage1_16[79]}
   );
   gpc606_5 gpc337 (
      {stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164], stage0_16[165]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[12],stage1_18[35],stage1_17[69],stage1_16[80]}
   );
   gpc606_5 gpc338 (
      {stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170], stage0_16[171]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[13],stage1_18[36],stage1_17[70],stage1_16[81]}
   );
   gpc606_5 gpc339 (
      {stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176], stage0_16[177]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[14],stage1_18[37],stage1_17[71],stage1_16[82]}
   );
   gpc606_5 gpc340 (
      {stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182], stage0_16[183]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[15],stage1_18[38],stage1_17[72],stage1_16[83]}
   );
   gpc606_5 gpc341 (
      {stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188], stage0_16[189]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[16],stage1_18[39],stage1_17[73],stage1_16[84]}
   );
   gpc606_5 gpc342 (
      {stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194], stage0_16[195]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[17],stage1_18[40],stage1_17[74],stage1_16[85]}
   );
   gpc606_5 gpc343 (
      {stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200], stage0_16[201]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[18],stage1_18[41],stage1_17[75],stage1_16[86]}
   );
   gpc606_5 gpc344 (
      {stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206], stage0_16[207]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[19],stage1_18[42],stage1_17[76],stage1_16[87]}
   );
   gpc606_5 gpc345 (
      {stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212], stage0_16[213]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[20],stage1_18[43],stage1_17[77],stage1_16[88]}
   );
   gpc606_5 gpc346 (
      {stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218], stage0_16[219]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[21],stage1_18[44],stage1_17[78],stage1_16[89]}
   );
   gpc606_5 gpc347 (
      {stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224], stage0_16[225]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[22],stage1_18[45],stage1_17[79],stage1_16[90]}
   );
   gpc606_5 gpc348 (
      {stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230], stage0_16[231]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[23],stage1_18[46],stage1_17[80],stage1_16[91]}
   );
   gpc606_5 gpc349 (
      {stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236], stage0_16[237]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[24],stage1_18[47],stage1_17[81],stage1_16[92]}
   );
   gpc606_5 gpc350 (
      {stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242], stage0_16[243]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[25],stage1_18[48],stage1_17[82],stage1_16[93]}
   );
   gpc606_5 gpc351 (
      {stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248], stage0_16[249]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[26],stage1_18[49],stage1_17[83],stage1_16[94]}
   );
   gpc606_5 gpc352 (
      {stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254], stage0_16[255]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[27],stage1_18[50],stage1_17[84],stage1_16[95]}
   );
   gpc606_5 gpc353 (
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[18],stage1_19[28],stage1_18[51],stage1_17[85]}
   );
   gpc606_5 gpc354 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[19],stage1_19[29],stage1_18[52],stage1_17[86]}
   );
   gpc615_5 gpc355 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76]},
      {stage0_18[108]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[20],stage1_19[30],stage1_18[53],stage1_17[87]}
   );
   gpc615_5 gpc356 (
      {stage0_17[77], stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81]},
      {stage0_18[109]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[21],stage1_19[31],stage1_18[54],stage1_17[88]}
   );
   gpc615_5 gpc357 (
      {stage0_17[82], stage0_17[83], stage0_17[84], stage0_17[85], stage0_17[86]},
      {stage0_18[110]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[22],stage1_19[32],stage1_18[55],stage1_17[89]}
   );
   gpc615_5 gpc358 (
      {stage0_17[87], stage0_17[88], stage0_17[89], stage0_17[90], stage0_17[91]},
      {stage0_18[111]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[23],stage1_19[33],stage1_18[56],stage1_17[90]}
   );
   gpc615_5 gpc359 (
      {stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95], stage0_17[96]},
      {stage0_18[112]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[24],stage1_19[34],stage1_18[57],stage1_17[91]}
   );
   gpc615_5 gpc360 (
      {stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_18[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[25],stage1_19[35],stage1_18[58],stage1_17[92]}
   );
   gpc615_5 gpc361 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106]},
      {stage0_18[114]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[26],stage1_19[36],stage1_18[59],stage1_17[93]}
   );
   gpc615_5 gpc362 (
      {stage0_17[107], stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111]},
      {stage0_18[115]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[27],stage1_19[37],stage1_18[60],stage1_17[94]}
   );
   gpc615_5 gpc363 (
      {stage0_17[112], stage0_17[113], stage0_17[114], stage0_17[115], stage0_17[116]},
      {stage0_18[116]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[28],stage1_19[38],stage1_18[61],stage1_17[95]}
   );
   gpc615_5 gpc364 (
      {stage0_17[117], stage0_17[118], stage0_17[119], stage0_17[120], stage0_17[121]},
      {stage0_18[117]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[29],stage1_19[39],stage1_18[62],stage1_17[96]}
   );
   gpc615_5 gpc365 (
      {stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125], stage0_17[126]},
      {stage0_18[118]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[30],stage1_19[40],stage1_18[63],stage1_17[97]}
   );
   gpc615_5 gpc366 (
      {stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_18[119]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[31],stage1_19[41],stage1_18[64],stage1_17[98]}
   );
   gpc615_5 gpc367 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136]},
      {stage0_18[120]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[32],stage1_19[42],stage1_18[65],stage1_17[99]}
   );
   gpc615_5 gpc368 (
      {stage0_17[137], stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141]},
      {stage0_18[121]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[33],stage1_19[43],stage1_18[66],stage1_17[100]}
   );
   gpc615_5 gpc369 (
      {stage0_17[142], stage0_17[143], stage0_17[144], stage0_17[145], stage0_17[146]},
      {stage0_18[122]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[34],stage1_19[44],stage1_18[67],stage1_17[101]}
   );
   gpc615_5 gpc370 (
      {stage0_17[147], stage0_17[148], stage0_17[149], stage0_17[150], stage0_17[151]},
      {stage0_18[123]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[35],stage1_19[45],stage1_18[68],stage1_17[102]}
   );
   gpc615_5 gpc371 (
      {stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155], stage0_17[156]},
      {stage0_18[124]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[36],stage1_19[46],stage1_18[69],stage1_17[103]}
   );
   gpc615_5 gpc372 (
      {stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_18[125]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[37],stage1_19[47],stage1_18[70],stage1_17[104]}
   );
   gpc615_5 gpc373 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166]},
      {stage0_18[126]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[38],stage1_19[48],stage1_18[71],stage1_17[105]}
   );
   gpc615_5 gpc374 (
      {stage0_17[167], stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171]},
      {stage0_18[127]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[39],stage1_19[49],stage1_18[72],stage1_17[106]}
   );
   gpc615_5 gpc375 (
      {stage0_17[172], stage0_17[173], stage0_17[174], stage0_17[175], stage0_17[176]},
      {stage0_18[128]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[40],stage1_19[50],stage1_18[73],stage1_17[107]}
   );
   gpc615_5 gpc376 (
      {stage0_17[177], stage0_17[178], stage0_17[179], stage0_17[180], stage0_17[181]},
      {stage0_18[129]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[41],stage1_19[51],stage1_18[74],stage1_17[108]}
   );
   gpc615_5 gpc377 (
      {stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185], stage0_17[186]},
      {stage0_18[130]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[42],stage1_19[52],stage1_18[75],stage1_17[109]}
   );
   gpc615_5 gpc378 (
      {stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_18[131]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[43],stage1_19[53],stage1_18[76],stage1_17[110]}
   );
   gpc615_5 gpc379 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196]},
      {stage0_18[132]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[44],stage1_19[54],stage1_18[77],stage1_17[111]}
   );
   gpc615_5 gpc380 (
      {stage0_17[197], stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201]},
      {stage0_18[133]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[45],stage1_19[55],stage1_18[78],stage1_17[112]}
   );
   gpc615_5 gpc381 (
      {stage0_17[202], stage0_17[203], stage0_17[204], stage0_17[205], stage0_17[206]},
      {stage0_18[134]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[46],stage1_19[56],stage1_18[79],stage1_17[113]}
   );
   gpc615_5 gpc382 (
      {stage0_17[207], stage0_17[208], stage0_17[209], stage0_17[210], stage0_17[211]},
      {stage0_18[135]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[47],stage1_19[57],stage1_18[80],stage1_17[114]}
   );
   gpc615_5 gpc383 (
      {stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215], stage0_17[216]},
      {stage0_18[136]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[48],stage1_19[58],stage1_18[81],stage1_17[115]}
   );
   gpc615_5 gpc384 (
      {stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_18[137]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[49],stage1_19[59],stage1_18[82],stage1_17[116]}
   );
   gpc615_5 gpc385 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226]},
      {stage0_18[138]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[50],stage1_19[60],stage1_18[83],stage1_17[117]}
   );
   gpc615_5 gpc386 (
      {stage0_17[227], stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231]},
      {stage0_18[139]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[51],stage1_19[61],stage1_18[84],stage1_17[118]}
   );
   gpc615_5 gpc387 (
      {stage0_17[232], stage0_17[233], stage0_17[234], stage0_17[235], stage0_17[236]},
      {stage0_18[140]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[52],stage1_19[62],stage1_18[85],stage1_17[119]}
   );
   gpc615_5 gpc388 (
      {stage0_17[237], stage0_17[238], stage0_17[239], stage0_17[240], stage0_17[241]},
      {stage0_18[141]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[53],stage1_19[63],stage1_18[86],stage1_17[120]}
   );
   gpc615_5 gpc389 (
      {stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245], stage0_17[246]},
      {stage0_18[142]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[54],stage1_19[64],stage1_18[87],stage1_17[121]}
   );
   gpc615_5 gpc390 (
      {stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_18[143]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[55],stage1_19[65],stage1_18[88],stage1_17[122]}
   );
   gpc606_5 gpc391 (
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[56],stage1_19[66],stage1_18[89]}
   );
   gpc606_5 gpc392 (
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[57],stage1_19[67],stage1_18[90]}
   );
   gpc606_5 gpc393 (
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[58],stage1_19[68],stage1_18[91]}
   );
   gpc606_5 gpc394 (
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[59],stage1_19[69],stage1_18[92]}
   );
   gpc606_5 gpc395 (
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[42],stage1_20[60],stage1_19[70],stage1_18[93]}
   );
   gpc606_5 gpc396 (
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[43],stage1_20[61],stage1_19[71],stage1_18[94]}
   );
   gpc606_5 gpc397 (
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[44],stage1_20[62],stage1_19[72],stage1_18[95]}
   );
   gpc606_5 gpc398 (
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[45],stage1_20[63],stage1_19[73],stage1_18[96]}
   );
   gpc606_5 gpc399 (
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[46],stage1_20[64],stage1_19[74],stage1_18[97]}
   );
   gpc606_5 gpc400 (
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[47],stage1_20[65],stage1_19[75],stage1_18[98]}
   );
   gpc606_5 gpc401 (
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[10],stage1_21[48],stage1_20[66],stage1_19[76]}
   );
   gpc606_5 gpc402 (
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[11],stage1_21[49],stage1_20[67],stage1_19[77]}
   );
   gpc615_5 gpc403 (
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[12],stage1_21[50],stage1_20[68]}
   );
   gpc615_5 gpc404 (
      {stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[13],stage1_21[51],stage1_20[69]}
   );
   gpc615_5 gpc405 (
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[14],stage1_21[52],stage1_20[70]}
   );
   gpc615_5 gpc406 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[15],stage1_21[53],stage1_20[71]}
   );
   gpc615_5 gpc407 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[16],stage1_21[54],stage1_20[72]}
   );
   gpc615_5 gpc408 (
      {stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[17],stage1_21[55],stage1_20[73]}
   );
   gpc615_5 gpc409 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[18],stage1_21[56],stage1_20[74]}
   );
   gpc615_5 gpc410 (
      {stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_21[19]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[19],stage1_21[57],stage1_20[75]}
   );
   gpc615_5 gpc411 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_21[20]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[10],stage1_22[20],stage1_21[58],stage1_20[76]}
   );
   gpc615_5 gpc412 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_21[21]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[11],stage1_22[21],stage1_21[59],stage1_20[77]}
   );
   gpc615_5 gpc413 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114]},
      {stage0_21[22]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[12],stage1_22[22],stage1_21[60],stage1_20[78]}
   );
   gpc615_5 gpc414 (
      {stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_21[23]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[13],stage1_22[23],stage1_21[61],stage1_20[79]}
   );
   gpc615_5 gpc415 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124]},
      {stage0_21[24]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[14],stage1_22[24],stage1_21[62],stage1_20[80]}
   );
   gpc615_5 gpc416 (
      {stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129]},
      {stage0_21[25]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[15],stage1_22[25],stage1_21[63],stage1_20[81]}
   );
   gpc615_5 gpc417 (
      {stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_21[26]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[16],stage1_22[26],stage1_21[64],stage1_20[82]}
   );
   gpc615_5 gpc418 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_21[27]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[17],stage1_22[27],stage1_21[65],stage1_20[83]}
   );
   gpc615_5 gpc419 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144]},
      {stage0_21[28]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[18],stage1_22[28],stage1_21[66],stage1_20[84]}
   );
   gpc615_5 gpc420 (
      {stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_21[29]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[19],stage1_22[29],stage1_21[67],stage1_20[85]}
   );
   gpc615_5 gpc421 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154]},
      {stage0_21[30]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[20],stage1_22[30],stage1_21[68],stage1_20[86]}
   );
   gpc615_5 gpc422 (
      {stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159]},
      {stage0_21[31]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[21],stage1_22[31],stage1_21[69],stage1_20[87]}
   );
   gpc615_5 gpc423 (
      {stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163], stage0_20[164]},
      {stage0_21[32]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[22],stage1_22[32],stage1_21[70],stage1_20[88]}
   );
   gpc615_5 gpc424 (
      {stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_21[33]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[23],stage1_22[33],stage1_21[71],stage1_20[89]}
   );
   gpc615_5 gpc425 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174]},
      {stage0_21[34]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[24],stage1_22[34],stage1_21[72],stage1_20[90]}
   );
   gpc615_5 gpc426 (
      {stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_21[35]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[25],stage1_22[35],stage1_21[73],stage1_20[91]}
   );
   gpc615_5 gpc427 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184]},
      {stage0_21[36]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[26],stage1_22[36],stage1_21[74],stage1_20[92]}
   );
   gpc615_5 gpc428 (
      {stage0_20[185], stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189]},
      {stage0_21[37]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[27],stage1_22[37],stage1_21[75],stage1_20[93]}
   );
   gpc615_5 gpc429 (
      {stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193], stage0_20[194]},
      {stage0_21[38]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[28],stage1_22[38],stage1_21[76],stage1_20[94]}
   );
   gpc615_5 gpc430 (
      {stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_21[39]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[29],stage1_22[39],stage1_21[77],stage1_20[95]}
   );
   gpc615_5 gpc431 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204]},
      {stage0_21[40]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[30],stage1_22[40],stage1_21[78],stage1_20[96]}
   );
   gpc615_5 gpc432 (
      {stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_21[41]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[31],stage1_22[41],stage1_21[79],stage1_20[97]}
   );
   gpc615_5 gpc433 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214]},
      {stage0_21[42]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[32],stage1_22[42],stage1_21[80],stage1_20[98]}
   );
   gpc615_5 gpc434 (
      {stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_21[43]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[33],stage1_22[43],stage1_21[81],stage1_20[99]}
   );
   gpc615_5 gpc435 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224]},
      {stage0_21[44]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[34],stage1_22[44],stage1_21[82],stage1_20[100]}
   );
   gpc615_5 gpc436 (
      {stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_21[45]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[35],stage1_22[45],stage1_21[83],stage1_20[101]}
   );
   gpc615_5 gpc437 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234]},
      {stage0_21[46]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[36],stage1_22[46],stage1_21[84],stage1_20[102]}
   );
   gpc615_5 gpc438 (
      {stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_21[47]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[37],stage1_22[47],stage1_21[85],stage1_20[103]}
   );
   gpc615_5 gpc439 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244]},
      {stage0_21[48]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[38],stage1_22[48],stage1_21[86],stage1_20[104]}
   );
   gpc606_5 gpc440 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[37],stage1_23[39],stage1_22[49],stage1_21[87]}
   );
   gpc606_5 gpc441 (
      {stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[38],stage1_23[40],stage1_22[50],stage1_21[88]}
   );
   gpc606_5 gpc442 (
      {stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[39],stage1_23[41],stage1_22[51],stage1_21[89]}
   );
   gpc606_5 gpc443 (
      {stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[40],stage1_23[42],stage1_22[52],stage1_21[90]}
   );
   gpc606_5 gpc444 (
      {stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[41],stage1_23[43],stage1_22[53],stage1_21[91]}
   );
   gpc606_5 gpc445 (
      {stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[42],stage1_23[44],stage1_22[54],stage1_21[92]}
   );
   gpc606_5 gpc446 (
      {stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[43],stage1_23[45],stage1_22[55],stage1_21[93]}
   );
   gpc606_5 gpc447 (
      {stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[44],stage1_23[46],stage1_22[56],stage1_21[94]}
   );
   gpc606_5 gpc448 (
      {stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[45],stage1_23[47],stage1_22[57],stage1_21[95]}
   );
   gpc606_5 gpc449 (
      {stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[46],stage1_23[48],stage1_22[58],stage1_21[96]}
   );
   gpc606_5 gpc450 (
      {stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[47],stage1_23[49],stage1_22[59],stage1_21[97]}
   );
   gpc606_5 gpc451 (
      {stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[48],stage1_23[50],stage1_22[60],stage1_21[98]}
   );
   gpc606_5 gpc452 (
      {stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[49],stage1_23[51],stage1_22[61],stage1_21[99]}
   );
   gpc606_5 gpc453 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131], stage0_21[132]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[50],stage1_23[52],stage1_22[62],stage1_21[100]}
   );
   gpc606_5 gpc454 (
      {stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137], stage0_21[138]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[51],stage1_23[53],stage1_22[63],stage1_21[101]}
   );
   gpc606_5 gpc455 (
      {stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143], stage0_21[144]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[52],stage1_23[54],stage1_22[64],stage1_21[102]}
   );
   gpc606_5 gpc456 (
      {stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149], stage0_21[150]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[53],stage1_23[55],stage1_22[65],stage1_21[103]}
   );
   gpc606_5 gpc457 (
      {stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155], stage0_21[156]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[54],stage1_23[56],stage1_22[66],stage1_21[104]}
   );
   gpc606_5 gpc458 (
      {stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161], stage0_21[162]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[55],stage1_23[57],stage1_22[67],stage1_21[105]}
   );
   gpc606_5 gpc459 (
      {stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167], stage0_21[168]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[56],stage1_23[58],stage1_22[68],stage1_21[106]}
   );
   gpc606_5 gpc460 (
      {stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173], stage0_21[174]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[57],stage1_23[59],stage1_22[69],stage1_21[107]}
   );
   gpc606_5 gpc461 (
      {stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179], stage0_21[180]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[58],stage1_23[60],stage1_22[70],stage1_21[108]}
   );
   gpc606_5 gpc462 (
      {stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185], stage0_21[186]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[59],stage1_23[61],stage1_22[71],stage1_21[109]}
   );
   gpc606_5 gpc463 (
      {stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191], stage0_21[192]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[60],stage1_23[62],stage1_22[72],stage1_21[110]}
   );
   gpc606_5 gpc464 (
      {stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197], stage0_21[198]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[61],stage1_23[63],stage1_22[73],stage1_21[111]}
   );
   gpc606_5 gpc465 (
      {stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203], stage0_21[204]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[62],stage1_23[64],stage1_22[74],stage1_21[112]}
   );
   gpc606_5 gpc466 (
      {stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209], stage0_21[210]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[63],stage1_23[65],stage1_22[75],stage1_21[113]}
   );
   gpc606_5 gpc467 (
      {stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215], stage0_21[216]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[64],stage1_23[66],stage1_22[76],stage1_21[114]}
   );
   gpc606_5 gpc468 (
      {stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221], stage0_21[222]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[65],stage1_23[67],stage1_22[77],stage1_21[115]}
   );
   gpc606_5 gpc469 (
      {stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227], stage0_21[228]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[66],stage1_23[68],stage1_22[78],stage1_21[116]}
   );
   gpc606_5 gpc470 (
      {stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233], stage0_21[234]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[67],stage1_23[69],stage1_22[79],stage1_21[117]}
   );
   gpc606_5 gpc471 (
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[31],stage1_24[68],stage1_23[70],stage1_22[80]}
   );
   gpc606_5 gpc472 (
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[32],stage1_24[69],stage1_23[71],stage1_22[81]}
   );
   gpc606_5 gpc473 (
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[33],stage1_24[70],stage1_23[72],stage1_22[82]}
   );
   gpc606_5 gpc474 (
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[34],stage1_24[71],stage1_23[73],stage1_22[83]}
   );
   gpc606_5 gpc475 (
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[4],stage1_25[35],stage1_24[72],stage1_23[74]}
   );
   gpc606_5 gpc476 (
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[5],stage1_25[36],stage1_24[73],stage1_23[75]}
   );
   gpc606_5 gpc477 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[6],stage1_25[37],stage1_24[74],stage1_23[76]}
   );
   gpc606_5 gpc478 (
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[7],stage1_25[38],stage1_24[75],stage1_23[77]}
   );
   gpc606_5 gpc479 (
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[8],stage1_25[39],stage1_24[76],stage1_23[78]}
   );
   gpc606_5 gpc480 (
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[9],stage1_25[40],stage1_24[77],stage1_23[79]}
   );
   gpc606_5 gpc481 (
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[10],stage1_25[41],stage1_24[78],stage1_23[80]}
   );
   gpc606_5 gpc482 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[11],stage1_25[42],stage1_24[79],stage1_23[81]}
   );
   gpc606_5 gpc483 (
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[12],stage1_25[43],stage1_24[80],stage1_23[82]}
   );
   gpc606_5 gpc484 (
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[13],stage1_25[44],stage1_24[81],stage1_23[83]}
   );
   gpc606_5 gpc485 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[14],stage1_25[45],stage1_24[82]}
   );
   gpc606_5 gpc486 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[15],stage1_25[46],stage1_24[83]}
   );
   gpc606_5 gpc487 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[16],stage1_25[47],stage1_24[84]}
   );
   gpc606_5 gpc488 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[17],stage1_25[48],stage1_24[85]}
   );
   gpc606_5 gpc489 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[18],stage1_25[49],stage1_24[86]}
   );
   gpc606_5 gpc490 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[19],stage1_25[50],stage1_24[87]}
   );
   gpc606_5 gpc491 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[20],stage1_25[51],stage1_24[88]}
   );
   gpc606_5 gpc492 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[21],stage1_25[52],stage1_24[89]}
   );
   gpc606_5 gpc493 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[22],stage1_25[53],stage1_24[90]}
   );
   gpc606_5 gpc494 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[23],stage1_25[54],stage1_24[91]}
   );
   gpc606_5 gpc495 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[24],stage1_25[55],stage1_24[92]}
   );
   gpc606_5 gpc496 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[25],stage1_25[56],stage1_24[93]}
   );
   gpc606_5 gpc497 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[12],stage1_27[22],stage1_26[26],stage1_25[57]}
   );
   gpc606_5 gpc498 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[13],stage1_27[23],stage1_26[27],stage1_25[58]}
   );
   gpc606_5 gpc499 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[14],stage1_27[24],stage1_26[28],stage1_25[59]}
   );
   gpc606_5 gpc500 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[15],stage1_27[25],stage1_26[29],stage1_25[60]}
   );
   gpc606_5 gpc501 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[16],stage1_27[26],stage1_26[30],stage1_25[61]}
   );
   gpc606_5 gpc502 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[17],stage1_27[27],stage1_26[31],stage1_25[62]}
   );
   gpc606_5 gpc503 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[18],stage1_27[28],stage1_26[32],stage1_25[63]}
   );
   gpc606_5 gpc504 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[19],stage1_27[29],stage1_26[33],stage1_25[64]}
   );
   gpc606_5 gpc505 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[20],stage1_27[30],stage1_26[34],stage1_25[65]}
   );
   gpc606_5 gpc506 (
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[21],stage1_27[31],stage1_26[35],stage1_25[66]}
   );
   gpc606_5 gpc507 (
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[22],stage1_27[32],stage1_26[36],stage1_25[67]}
   );
   gpc606_5 gpc508 (
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[23],stage1_27[33],stage1_26[37],stage1_25[68]}
   );
   gpc606_5 gpc509 (
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[24],stage1_27[34],stage1_26[38],stage1_25[69]}
   );
   gpc606_5 gpc510 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[25],stage1_27[35],stage1_26[39],stage1_25[70]}
   );
   gpc606_5 gpc511 (
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[26],stage1_27[36],stage1_26[40],stage1_25[71]}
   );
   gpc606_5 gpc512 (
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[27],stage1_27[37],stage1_26[41],stage1_25[72]}
   );
   gpc606_5 gpc513 (
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[28],stage1_27[38],stage1_26[42],stage1_25[73]}
   );
   gpc606_5 gpc514 (
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[29],stage1_27[39],stage1_26[43],stage1_25[74]}
   );
   gpc606_5 gpc515 (
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[30],stage1_27[40],stage1_26[44],stage1_25[75]}
   );
   gpc606_5 gpc516 (
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[31],stage1_27[41],stage1_26[45],stage1_25[76]}
   );
   gpc606_5 gpc517 (
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[32],stage1_27[42],stage1_26[46],stage1_25[77]}
   );
   gpc606_5 gpc518 (
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[33],stage1_27[43],stage1_26[47],stage1_25[78]}
   );
   gpc606_5 gpc519 (
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[34],stage1_27[44],stage1_26[48],stage1_25[79]}
   );
   gpc606_5 gpc520 (
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[35],stage1_27[45],stage1_26[49],stage1_25[80]}
   );
   gpc606_5 gpc521 (
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[36],stage1_27[46],stage1_26[50],stage1_25[81]}
   );
   gpc606_5 gpc522 (
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[37],stage1_27[47],stage1_26[51],stage1_25[82]}
   );
   gpc606_5 gpc523 (
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[38],stage1_27[48],stage1_26[52],stage1_25[83]}
   );
   gpc606_5 gpc524 (
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[27],stage1_28[39],stage1_27[49]}
   );
   gpc606_5 gpc525 (
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[28],stage1_28[40],stage1_27[50]}
   );
   gpc606_5 gpc526 (
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[29],stage1_28[41],stage1_27[51]}
   );
   gpc606_5 gpc527 (
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[30],stage1_28[42],stage1_27[52]}
   );
   gpc606_5 gpc528 (
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[31],stage1_28[43],stage1_27[53]}
   );
   gpc606_5 gpc529 (
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[32],stage1_28[44],stage1_27[54]}
   );
   gpc606_5 gpc530 (
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[33],stage1_28[45],stage1_27[55]}
   );
   gpc606_5 gpc531 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[34],stage1_28[46]}
   );
   gpc606_5 gpc532 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[35],stage1_28[47]}
   );
   gpc606_5 gpc533 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[36],stage1_28[48]}
   );
   gpc606_5 gpc534 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[37],stage1_28[49]}
   );
   gpc606_5 gpc535 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[38],stage1_28[50]}
   );
   gpc606_5 gpc536 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[39],stage1_28[51]}
   );
   gpc606_5 gpc537 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[40],stage1_28[52]}
   );
   gpc606_5 gpc538 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[41],stage1_28[53]}
   );
   gpc606_5 gpc539 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[42],stage1_28[54]}
   );
   gpc606_5 gpc540 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[43],stage1_28[55]}
   );
   gpc606_5 gpc541 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[44],stage1_28[56]}
   );
   gpc606_5 gpc542 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[45],stage1_28[57]}
   );
   gpc606_5 gpc543 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[46],stage1_28[58]}
   );
   gpc606_5 gpc544 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[47],stage1_28[59]}
   );
   gpc606_5 gpc545 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[48],stage1_28[60]}
   );
   gpc606_5 gpc546 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[49],stage1_28[61]}
   );
   gpc606_5 gpc547 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[50],stage1_28[62]}
   );
   gpc606_5 gpc548 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[51],stage1_28[63]}
   );
   gpc606_5 gpc549 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[52],stage1_28[64]}
   );
   gpc606_5 gpc550 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[53],stage1_28[65]}
   );
   gpc606_5 gpc551 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[54],stage1_28[66]}
   );
   gpc606_5 gpc552 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[55],stage1_28[67]}
   );
   gpc606_5 gpc553 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[56],stage1_28[68]}
   );
   gpc606_5 gpc554 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[57],stage1_28[69]}
   );
   gpc606_5 gpc555 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[58],stage1_28[70]}
   );
   gpc606_5 gpc556 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[59],stage1_28[71]}
   );
   gpc606_5 gpc557 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[60],stage1_28[72]}
   );
   gpc606_5 gpc558 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[61],stage1_28[73]}
   );
   gpc606_5 gpc559 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[62],stage1_28[74]}
   );
   gpc606_5 gpc560 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[63],stage1_28[75]}
   );
   gpc606_5 gpc561 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[64],stage1_28[76]}
   );
   gpc606_5 gpc562 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[65],stage1_28[77]}
   );
   gpc606_5 gpc563 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[66],stage1_28[78]}
   );
   gpc606_5 gpc564 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[67],stage1_28[79]}
   );
   gpc606_5 gpc565 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[68],stage1_28[80]}
   );
   gpc606_5 gpc566 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[69],stage1_28[81]}
   );
   gpc606_5 gpc567 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[70],stage1_28[82]}
   );
   gpc606_5 gpc568 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[71],stage1_28[83]}
   );
   gpc606_5 gpc569 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[72],stage1_28[84]}
   );
   gpc606_5 gpc570 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[73],stage1_28[85]}
   );
   gpc606_5 gpc571 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[74]}
   );
   gpc606_5 gpc572 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[75]}
   );
   gpc606_5 gpc573 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[76]}
   );
   gpc606_5 gpc574 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[77]}
   );
   gpc606_5 gpc575 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[78]}
   );
   gpc606_5 gpc576 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[45],stage1_31[52],stage1_30[52],stage1_29[79]}
   );
   gpc606_5 gpc577 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[46],stage1_31[53],stage1_30[53],stage1_29[80]}
   );
   gpc606_5 gpc578 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[47],stage1_31[54],stage1_30[54],stage1_29[81]}
   );
   gpc606_5 gpc579 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[48],stage1_31[55],stage1_30[55],stage1_29[82]}
   );
   gpc606_5 gpc580 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[49],stage1_31[56],stage1_30[56],stage1_29[83]}
   );
   gpc606_5 gpc581 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[50],stage1_31[57],stage1_30[57],stage1_29[84]}
   );
   gpc606_5 gpc582 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[51],stage1_31[58],stage1_30[58],stage1_29[85]}
   );
   gpc606_5 gpc583 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[52],stage1_31[59],stage1_30[59],stage1_29[86]}
   );
   gpc606_5 gpc584 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[53],stage1_31[60],stage1_30[60],stage1_29[87]}
   );
   gpc606_5 gpc585 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[54],stage1_31[61],stage1_30[61],stage1_29[88]}
   );
   gpc606_5 gpc586 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[55],stage1_31[62],stage1_30[62],stage1_29[89]}
   );
   gpc606_5 gpc587 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[56],stage1_31[63],stage1_30[63],stage1_29[90]}
   );
   gpc606_5 gpc588 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[57],stage1_31[64],stage1_30[64],stage1_29[91]}
   );
   gpc606_5 gpc589 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[58],stage1_31[65],stage1_30[65],stage1_29[92]}
   );
   gpc606_5 gpc590 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[59],stage1_31[66],stage1_30[66],stage1_29[93]}
   );
   gpc606_5 gpc591 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[60],stage1_31[67],stage1_30[67],stage1_29[94]}
   );
   gpc606_5 gpc592 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[61],stage1_31[68],stage1_30[68],stage1_29[95]}
   );
   gpc606_5 gpc593 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[62],stage1_31[69],stage1_30[69],stage1_29[96]}
   );
   gpc606_5 gpc594 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[63],stage1_31[70],stage1_30[70],stage1_29[97]}
   );
   gpc606_5 gpc595 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[64],stage1_31[71],stage1_30[71],stage1_29[98]}
   );
   gpc606_5 gpc596 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[65],stage1_31[72],stage1_30[72],stage1_29[99]}
   );
   gpc606_5 gpc597 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[66],stage1_31[73],stage1_30[73],stage1_29[100]}
   );
   gpc606_5 gpc598 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[67],stage1_31[74],stage1_30[74],stage1_29[101]}
   );
   gpc606_5 gpc599 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[68],stage1_31[75],stage1_30[75],stage1_29[102]}
   );
   gpc606_5 gpc600 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[69],stage1_31[76],stage1_30[76],stage1_29[103]}
   );
   gpc606_5 gpc601 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[70],stage1_31[77],stage1_30[77],stage1_29[104]}
   );
   gpc606_5 gpc602 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[71],stage1_31[78],stage1_30[78],stage1_29[105]}
   );
   gpc606_5 gpc603 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[72],stage1_31[79],stage1_30[79],stage1_29[106]}
   );
   gpc606_5 gpc604 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[73],stage1_31[80],stage1_30[80],stage1_29[107]}
   );
   gpc1_1 gpc605 (
      {stage0_0[249]},
      {stage1_0[43]}
   );
   gpc1_1 gpc606 (
      {stage0_0[250]},
      {stage1_0[44]}
   );
   gpc1_1 gpc607 (
      {stage0_0[251]},
      {stage1_0[45]}
   );
   gpc1_1 gpc608 (
      {stage0_0[252]},
      {stage1_0[46]}
   );
   gpc1_1 gpc609 (
      {stage0_0[253]},
      {stage1_0[47]}
   );
   gpc1_1 gpc610 (
      {stage0_0[254]},
      {stage1_0[48]}
   );
   gpc1_1 gpc611 (
      {stage0_0[255]},
      {stage1_0[49]}
   );
   gpc1_1 gpc612 (
      {stage0_1[237]},
      {stage1_1[79]}
   );
   gpc1_1 gpc613 (
      {stage0_1[238]},
      {stage1_1[80]}
   );
   gpc1_1 gpc614 (
      {stage0_1[239]},
      {stage1_1[81]}
   );
   gpc1_1 gpc615 (
      {stage0_1[240]},
      {stage1_1[82]}
   );
   gpc1_1 gpc616 (
      {stage0_1[241]},
      {stage1_1[83]}
   );
   gpc1_1 gpc617 (
      {stage0_1[242]},
      {stage1_1[84]}
   );
   gpc1_1 gpc618 (
      {stage0_1[243]},
      {stage1_1[85]}
   );
   gpc1_1 gpc619 (
      {stage0_1[244]},
      {stage1_1[86]}
   );
   gpc1_1 gpc620 (
      {stage0_1[245]},
      {stage1_1[87]}
   );
   gpc1_1 gpc621 (
      {stage0_1[246]},
      {stage1_1[88]}
   );
   gpc1_1 gpc622 (
      {stage0_1[247]},
      {stage1_1[89]}
   );
   gpc1_1 gpc623 (
      {stage0_1[248]},
      {stage1_1[90]}
   );
   gpc1_1 gpc624 (
      {stage0_1[249]},
      {stage1_1[91]}
   );
   gpc1_1 gpc625 (
      {stage0_1[250]},
      {stage1_1[92]}
   );
   gpc1_1 gpc626 (
      {stage0_1[251]},
      {stage1_1[93]}
   );
   gpc1_1 gpc627 (
      {stage0_1[252]},
      {stage1_1[94]}
   );
   gpc1_1 gpc628 (
      {stage0_1[253]},
      {stage1_1[95]}
   );
   gpc1_1 gpc629 (
      {stage0_1[254]},
      {stage1_1[96]}
   );
   gpc1_1 gpc630 (
      {stage0_1[255]},
      {stage1_1[97]}
   );
   gpc1_1 gpc631 (
      {stage0_2[246]},
      {stage1_2[82]}
   );
   gpc1_1 gpc632 (
      {stage0_2[247]},
      {stage1_2[83]}
   );
   gpc1_1 gpc633 (
      {stage0_2[248]},
      {stage1_2[84]}
   );
   gpc1_1 gpc634 (
      {stage0_2[249]},
      {stage1_2[85]}
   );
   gpc1_1 gpc635 (
      {stage0_2[250]},
      {stage1_2[86]}
   );
   gpc1_1 gpc636 (
      {stage0_2[251]},
      {stage1_2[87]}
   );
   gpc1_1 gpc637 (
      {stage0_2[252]},
      {stage1_2[88]}
   );
   gpc1_1 gpc638 (
      {stage0_2[253]},
      {stage1_2[89]}
   );
   gpc1_1 gpc639 (
      {stage0_2[254]},
      {stage1_2[90]}
   );
   gpc1_1 gpc640 (
      {stage0_2[255]},
      {stage1_2[91]}
   );
   gpc1_1 gpc641 (
      {stage0_3[254]},
      {stage1_3[89]}
   );
   gpc1_1 gpc642 (
      {stage0_3[255]},
      {stage1_3[90]}
   );
   gpc1_1 gpc643 (
      {stage0_4[230]},
      {stage1_4[123]}
   );
   gpc1_1 gpc644 (
      {stage0_4[231]},
      {stage1_4[124]}
   );
   gpc1_1 gpc645 (
      {stage0_4[232]},
      {stage1_4[125]}
   );
   gpc1_1 gpc646 (
      {stage0_4[233]},
      {stage1_4[126]}
   );
   gpc1_1 gpc647 (
      {stage0_4[234]},
      {stage1_4[127]}
   );
   gpc1_1 gpc648 (
      {stage0_4[235]},
      {stage1_4[128]}
   );
   gpc1_1 gpc649 (
      {stage0_4[236]},
      {stage1_4[129]}
   );
   gpc1_1 gpc650 (
      {stage0_4[237]},
      {stage1_4[130]}
   );
   gpc1_1 gpc651 (
      {stage0_4[238]},
      {stage1_4[131]}
   );
   gpc1_1 gpc652 (
      {stage0_4[239]},
      {stage1_4[132]}
   );
   gpc1_1 gpc653 (
      {stage0_4[240]},
      {stage1_4[133]}
   );
   gpc1_1 gpc654 (
      {stage0_4[241]},
      {stage1_4[134]}
   );
   gpc1_1 gpc655 (
      {stage0_4[242]},
      {stage1_4[135]}
   );
   gpc1_1 gpc656 (
      {stage0_4[243]},
      {stage1_4[136]}
   );
   gpc1_1 gpc657 (
      {stage0_4[244]},
      {stage1_4[137]}
   );
   gpc1_1 gpc658 (
      {stage0_4[245]},
      {stage1_4[138]}
   );
   gpc1_1 gpc659 (
      {stage0_4[246]},
      {stage1_4[139]}
   );
   gpc1_1 gpc660 (
      {stage0_4[247]},
      {stage1_4[140]}
   );
   gpc1_1 gpc661 (
      {stage0_4[248]},
      {stage1_4[141]}
   );
   gpc1_1 gpc662 (
      {stage0_4[249]},
      {stage1_4[142]}
   );
   gpc1_1 gpc663 (
      {stage0_4[250]},
      {stage1_4[143]}
   );
   gpc1_1 gpc664 (
      {stage0_4[251]},
      {stage1_4[144]}
   );
   gpc1_1 gpc665 (
      {stage0_4[252]},
      {stage1_4[145]}
   );
   gpc1_1 gpc666 (
      {stage0_4[253]},
      {stage1_4[146]}
   );
   gpc1_1 gpc667 (
      {stage0_4[254]},
      {stage1_4[147]}
   );
   gpc1_1 gpc668 (
      {stage0_4[255]},
      {stage1_4[148]}
   );
   gpc1_1 gpc669 (
      {stage0_5[240]},
      {stage1_5[110]}
   );
   gpc1_1 gpc670 (
      {stage0_5[241]},
      {stage1_5[111]}
   );
   gpc1_1 gpc671 (
      {stage0_5[242]},
      {stage1_5[112]}
   );
   gpc1_1 gpc672 (
      {stage0_5[243]},
      {stage1_5[113]}
   );
   gpc1_1 gpc673 (
      {stage0_5[244]},
      {stage1_5[114]}
   );
   gpc1_1 gpc674 (
      {stage0_5[245]},
      {stage1_5[115]}
   );
   gpc1_1 gpc675 (
      {stage0_5[246]},
      {stage1_5[116]}
   );
   gpc1_1 gpc676 (
      {stage0_5[247]},
      {stage1_5[117]}
   );
   gpc1_1 gpc677 (
      {stage0_5[248]},
      {stage1_5[118]}
   );
   gpc1_1 gpc678 (
      {stage0_5[249]},
      {stage1_5[119]}
   );
   gpc1_1 gpc679 (
      {stage0_5[250]},
      {stage1_5[120]}
   );
   gpc1_1 gpc680 (
      {stage0_5[251]},
      {stage1_5[121]}
   );
   gpc1_1 gpc681 (
      {stage0_5[252]},
      {stage1_5[122]}
   );
   gpc1_1 gpc682 (
      {stage0_5[253]},
      {stage1_5[123]}
   );
   gpc1_1 gpc683 (
      {stage0_5[254]},
      {stage1_5[124]}
   );
   gpc1_1 gpc684 (
      {stage0_5[255]},
      {stage1_5[125]}
   );
   gpc1_1 gpc685 (
      {stage0_6[243]},
      {stage1_6[83]}
   );
   gpc1_1 gpc686 (
      {stage0_6[244]},
      {stage1_6[84]}
   );
   gpc1_1 gpc687 (
      {stage0_6[245]},
      {stage1_6[85]}
   );
   gpc1_1 gpc688 (
      {stage0_6[246]},
      {stage1_6[86]}
   );
   gpc1_1 gpc689 (
      {stage0_6[247]},
      {stage1_6[87]}
   );
   gpc1_1 gpc690 (
      {stage0_6[248]},
      {stage1_6[88]}
   );
   gpc1_1 gpc691 (
      {stage0_6[249]},
      {stage1_6[89]}
   );
   gpc1_1 gpc692 (
      {stage0_6[250]},
      {stage1_6[90]}
   );
   gpc1_1 gpc693 (
      {stage0_6[251]},
      {stage1_6[91]}
   );
   gpc1_1 gpc694 (
      {stage0_6[252]},
      {stage1_6[92]}
   );
   gpc1_1 gpc695 (
      {stage0_6[253]},
      {stage1_6[93]}
   );
   gpc1_1 gpc696 (
      {stage0_6[254]},
      {stage1_6[94]}
   );
   gpc1_1 gpc697 (
      {stage0_6[255]},
      {stage1_6[95]}
   );
   gpc1_1 gpc698 (
      {stage0_7[251]},
      {stage1_7[96]}
   );
   gpc1_1 gpc699 (
      {stage0_7[252]},
      {stage1_7[97]}
   );
   gpc1_1 gpc700 (
      {stage0_7[253]},
      {stage1_7[98]}
   );
   gpc1_1 gpc701 (
      {stage0_7[254]},
      {stage1_7[99]}
   );
   gpc1_1 gpc702 (
      {stage0_7[255]},
      {stage1_7[100]}
   );
   gpc1_1 gpc703 (
      {stage0_9[230]},
      {stage1_9[106]}
   );
   gpc1_1 gpc704 (
      {stage0_9[231]},
      {stage1_9[107]}
   );
   gpc1_1 gpc705 (
      {stage0_9[232]},
      {stage1_9[108]}
   );
   gpc1_1 gpc706 (
      {stage0_9[233]},
      {stage1_9[109]}
   );
   gpc1_1 gpc707 (
      {stage0_9[234]},
      {stage1_9[110]}
   );
   gpc1_1 gpc708 (
      {stage0_9[235]},
      {stage1_9[111]}
   );
   gpc1_1 gpc709 (
      {stage0_9[236]},
      {stage1_9[112]}
   );
   gpc1_1 gpc710 (
      {stage0_9[237]},
      {stage1_9[113]}
   );
   gpc1_1 gpc711 (
      {stage0_9[238]},
      {stage1_9[114]}
   );
   gpc1_1 gpc712 (
      {stage0_9[239]},
      {stage1_9[115]}
   );
   gpc1_1 gpc713 (
      {stage0_9[240]},
      {stage1_9[116]}
   );
   gpc1_1 gpc714 (
      {stage0_9[241]},
      {stage1_9[117]}
   );
   gpc1_1 gpc715 (
      {stage0_9[242]},
      {stage1_9[118]}
   );
   gpc1_1 gpc716 (
      {stage0_9[243]},
      {stage1_9[119]}
   );
   gpc1_1 gpc717 (
      {stage0_9[244]},
      {stage1_9[120]}
   );
   gpc1_1 gpc718 (
      {stage0_9[245]},
      {stage1_9[121]}
   );
   gpc1_1 gpc719 (
      {stage0_9[246]},
      {stage1_9[122]}
   );
   gpc1_1 gpc720 (
      {stage0_9[247]},
      {stage1_9[123]}
   );
   gpc1_1 gpc721 (
      {stage0_9[248]},
      {stage1_9[124]}
   );
   gpc1_1 gpc722 (
      {stage0_9[249]},
      {stage1_9[125]}
   );
   gpc1_1 gpc723 (
      {stage0_9[250]},
      {stage1_9[126]}
   );
   gpc1_1 gpc724 (
      {stage0_9[251]},
      {stage1_9[127]}
   );
   gpc1_1 gpc725 (
      {stage0_9[252]},
      {stage1_9[128]}
   );
   gpc1_1 gpc726 (
      {stage0_9[253]},
      {stage1_9[129]}
   );
   gpc1_1 gpc727 (
      {stage0_9[254]},
      {stage1_9[130]}
   );
   gpc1_1 gpc728 (
      {stage0_9[255]},
      {stage1_9[131]}
   );
   gpc1_1 gpc729 (
      {stage0_10[250]},
      {stage1_10[91]}
   );
   gpc1_1 gpc730 (
      {stage0_10[251]},
      {stage1_10[92]}
   );
   gpc1_1 gpc731 (
      {stage0_10[252]},
      {stage1_10[93]}
   );
   gpc1_1 gpc732 (
      {stage0_10[253]},
      {stage1_10[94]}
   );
   gpc1_1 gpc733 (
      {stage0_10[254]},
      {stage1_10[95]}
   );
   gpc1_1 gpc734 (
      {stage0_10[255]},
      {stage1_10[96]}
   );
   gpc1_1 gpc735 (
      {stage0_11[210]},
      {stage1_11[94]}
   );
   gpc1_1 gpc736 (
      {stage0_11[211]},
      {stage1_11[95]}
   );
   gpc1_1 gpc737 (
      {stage0_11[212]},
      {stage1_11[96]}
   );
   gpc1_1 gpc738 (
      {stage0_11[213]},
      {stage1_11[97]}
   );
   gpc1_1 gpc739 (
      {stage0_11[214]},
      {stage1_11[98]}
   );
   gpc1_1 gpc740 (
      {stage0_11[215]},
      {stage1_11[99]}
   );
   gpc1_1 gpc741 (
      {stage0_11[216]},
      {stage1_11[100]}
   );
   gpc1_1 gpc742 (
      {stage0_11[217]},
      {stage1_11[101]}
   );
   gpc1_1 gpc743 (
      {stage0_11[218]},
      {stage1_11[102]}
   );
   gpc1_1 gpc744 (
      {stage0_11[219]},
      {stage1_11[103]}
   );
   gpc1_1 gpc745 (
      {stage0_11[220]},
      {stage1_11[104]}
   );
   gpc1_1 gpc746 (
      {stage0_11[221]},
      {stage1_11[105]}
   );
   gpc1_1 gpc747 (
      {stage0_11[222]},
      {stage1_11[106]}
   );
   gpc1_1 gpc748 (
      {stage0_11[223]},
      {stage1_11[107]}
   );
   gpc1_1 gpc749 (
      {stage0_11[224]},
      {stage1_11[108]}
   );
   gpc1_1 gpc750 (
      {stage0_11[225]},
      {stage1_11[109]}
   );
   gpc1_1 gpc751 (
      {stage0_11[226]},
      {stage1_11[110]}
   );
   gpc1_1 gpc752 (
      {stage0_11[227]},
      {stage1_11[111]}
   );
   gpc1_1 gpc753 (
      {stage0_11[228]},
      {stage1_11[112]}
   );
   gpc1_1 gpc754 (
      {stage0_11[229]},
      {stage1_11[113]}
   );
   gpc1_1 gpc755 (
      {stage0_11[230]},
      {stage1_11[114]}
   );
   gpc1_1 gpc756 (
      {stage0_11[231]},
      {stage1_11[115]}
   );
   gpc1_1 gpc757 (
      {stage0_11[232]},
      {stage1_11[116]}
   );
   gpc1_1 gpc758 (
      {stage0_11[233]},
      {stage1_11[117]}
   );
   gpc1_1 gpc759 (
      {stage0_11[234]},
      {stage1_11[118]}
   );
   gpc1_1 gpc760 (
      {stage0_11[235]},
      {stage1_11[119]}
   );
   gpc1_1 gpc761 (
      {stage0_11[236]},
      {stage1_11[120]}
   );
   gpc1_1 gpc762 (
      {stage0_11[237]},
      {stage1_11[121]}
   );
   gpc1_1 gpc763 (
      {stage0_11[238]},
      {stage1_11[122]}
   );
   gpc1_1 gpc764 (
      {stage0_11[239]},
      {stage1_11[123]}
   );
   gpc1_1 gpc765 (
      {stage0_11[240]},
      {stage1_11[124]}
   );
   gpc1_1 gpc766 (
      {stage0_11[241]},
      {stage1_11[125]}
   );
   gpc1_1 gpc767 (
      {stage0_11[242]},
      {stage1_11[126]}
   );
   gpc1_1 gpc768 (
      {stage0_11[243]},
      {stage1_11[127]}
   );
   gpc1_1 gpc769 (
      {stage0_11[244]},
      {stage1_11[128]}
   );
   gpc1_1 gpc770 (
      {stage0_11[245]},
      {stage1_11[129]}
   );
   gpc1_1 gpc771 (
      {stage0_11[246]},
      {stage1_11[130]}
   );
   gpc1_1 gpc772 (
      {stage0_11[247]},
      {stage1_11[131]}
   );
   gpc1_1 gpc773 (
      {stage0_11[248]},
      {stage1_11[132]}
   );
   gpc1_1 gpc774 (
      {stage0_11[249]},
      {stage1_11[133]}
   );
   gpc1_1 gpc775 (
      {stage0_11[250]},
      {stage1_11[134]}
   );
   gpc1_1 gpc776 (
      {stage0_11[251]},
      {stage1_11[135]}
   );
   gpc1_1 gpc777 (
      {stage0_11[252]},
      {stage1_11[136]}
   );
   gpc1_1 gpc778 (
      {stage0_11[253]},
      {stage1_11[137]}
   );
   gpc1_1 gpc779 (
      {stage0_11[254]},
      {stage1_11[138]}
   );
   gpc1_1 gpc780 (
      {stage0_11[255]},
      {stage1_11[139]}
   );
   gpc1_1 gpc781 (
      {stage0_12[148]},
      {stage1_12[90]}
   );
   gpc1_1 gpc782 (
      {stage0_12[149]},
      {stage1_12[91]}
   );
   gpc1_1 gpc783 (
      {stage0_12[150]},
      {stage1_12[92]}
   );
   gpc1_1 gpc784 (
      {stage0_12[151]},
      {stage1_12[93]}
   );
   gpc1_1 gpc785 (
      {stage0_12[152]},
      {stage1_12[94]}
   );
   gpc1_1 gpc786 (
      {stage0_12[153]},
      {stage1_12[95]}
   );
   gpc1_1 gpc787 (
      {stage0_12[154]},
      {stage1_12[96]}
   );
   gpc1_1 gpc788 (
      {stage0_12[155]},
      {stage1_12[97]}
   );
   gpc1_1 gpc789 (
      {stage0_12[156]},
      {stage1_12[98]}
   );
   gpc1_1 gpc790 (
      {stage0_12[157]},
      {stage1_12[99]}
   );
   gpc1_1 gpc791 (
      {stage0_12[158]},
      {stage1_12[100]}
   );
   gpc1_1 gpc792 (
      {stage0_12[159]},
      {stage1_12[101]}
   );
   gpc1_1 gpc793 (
      {stage0_12[160]},
      {stage1_12[102]}
   );
   gpc1_1 gpc794 (
      {stage0_12[161]},
      {stage1_12[103]}
   );
   gpc1_1 gpc795 (
      {stage0_12[162]},
      {stage1_12[104]}
   );
   gpc1_1 gpc796 (
      {stage0_12[163]},
      {stage1_12[105]}
   );
   gpc1_1 gpc797 (
      {stage0_12[164]},
      {stage1_12[106]}
   );
   gpc1_1 gpc798 (
      {stage0_12[165]},
      {stage1_12[107]}
   );
   gpc1_1 gpc799 (
      {stage0_12[166]},
      {stage1_12[108]}
   );
   gpc1_1 gpc800 (
      {stage0_12[167]},
      {stage1_12[109]}
   );
   gpc1_1 gpc801 (
      {stage0_12[168]},
      {stage1_12[110]}
   );
   gpc1_1 gpc802 (
      {stage0_12[169]},
      {stage1_12[111]}
   );
   gpc1_1 gpc803 (
      {stage0_12[170]},
      {stage1_12[112]}
   );
   gpc1_1 gpc804 (
      {stage0_12[171]},
      {stage1_12[113]}
   );
   gpc1_1 gpc805 (
      {stage0_12[172]},
      {stage1_12[114]}
   );
   gpc1_1 gpc806 (
      {stage0_12[173]},
      {stage1_12[115]}
   );
   gpc1_1 gpc807 (
      {stage0_12[174]},
      {stage1_12[116]}
   );
   gpc1_1 gpc808 (
      {stage0_12[175]},
      {stage1_12[117]}
   );
   gpc1_1 gpc809 (
      {stage0_12[176]},
      {stage1_12[118]}
   );
   gpc1_1 gpc810 (
      {stage0_12[177]},
      {stage1_12[119]}
   );
   gpc1_1 gpc811 (
      {stage0_12[178]},
      {stage1_12[120]}
   );
   gpc1_1 gpc812 (
      {stage0_12[179]},
      {stage1_12[121]}
   );
   gpc1_1 gpc813 (
      {stage0_12[180]},
      {stage1_12[122]}
   );
   gpc1_1 gpc814 (
      {stage0_12[181]},
      {stage1_12[123]}
   );
   gpc1_1 gpc815 (
      {stage0_12[182]},
      {stage1_12[124]}
   );
   gpc1_1 gpc816 (
      {stage0_12[183]},
      {stage1_12[125]}
   );
   gpc1_1 gpc817 (
      {stage0_12[184]},
      {stage1_12[126]}
   );
   gpc1_1 gpc818 (
      {stage0_12[185]},
      {stage1_12[127]}
   );
   gpc1_1 gpc819 (
      {stage0_12[186]},
      {stage1_12[128]}
   );
   gpc1_1 gpc820 (
      {stage0_12[187]},
      {stage1_12[129]}
   );
   gpc1_1 gpc821 (
      {stage0_12[188]},
      {stage1_12[130]}
   );
   gpc1_1 gpc822 (
      {stage0_12[189]},
      {stage1_12[131]}
   );
   gpc1_1 gpc823 (
      {stage0_12[190]},
      {stage1_12[132]}
   );
   gpc1_1 gpc824 (
      {stage0_12[191]},
      {stage1_12[133]}
   );
   gpc1_1 gpc825 (
      {stage0_12[192]},
      {stage1_12[134]}
   );
   gpc1_1 gpc826 (
      {stage0_12[193]},
      {stage1_12[135]}
   );
   gpc1_1 gpc827 (
      {stage0_12[194]},
      {stage1_12[136]}
   );
   gpc1_1 gpc828 (
      {stage0_12[195]},
      {stage1_12[137]}
   );
   gpc1_1 gpc829 (
      {stage0_12[196]},
      {stage1_12[138]}
   );
   gpc1_1 gpc830 (
      {stage0_12[197]},
      {stage1_12[139]}
   );
   gpc1_1 gpc831 (
      {stage0_12[198]},
      {stage1_12[140]}
   );
   gpc1_1 gpc832 (
      {stage0_12[199]},
      {stage1_12[141]}
   );
   gpc1_1 gpc833 (
      {stage0_12[200]},
      {stage1_12[142]}
   );
   gpc1_1 gpc834 (
      {stage0_12[201]},
      {stage1_12[143]}
   );
   gpc1_1 gpc835 (
      {stage0_12[202]},
      {stage1_12[144]}
   );
   gpc1_1 gpc836 (
      {stage0_12[203]},
      {stage1_12[145]}
   );
   gpc1_1 gpc837 (
      {stage0_12[204]},
      {stage1_12[146]}
   );
   gpc1_1 gpc838 (
      {stage0_12[205]},
      {stage1_12[147]}
   );
   gpc1_1 gpc839 (
      {stage0_12[206]},
      {stage1_12[148]}
   );
   gpc1_1 gpc840 (
      {stage0_12[207]},
      {stage1_12[149]}
   );
   gpc1_1 gpc841 (
      {stage0_12[208]},
      {stage1_12[150]}
   );
   gpc1_1 gpc842 (
      {stage0_12[209]},
      {stage1_12[151]}
   );
   gpc1_1 gpc843 (
      {stage0_12[210]},
      {stage1_12[152]}
   );
   gpc1_1 gpc844 (
      {stage0_12[211]},
      {stage1_12[153]}
   );
   gpc1_1 gpc845 (
      {stage0_12[212]},
      {stage1_12[154]}
   );
   gpc1_1 gpc846 (
      {stage0_12[213]},
      {stage1_12[155]}
   );
   gpc1_1 gpc847 (
      {stage0_12[214]},
      {stage1_12[156]}
   );
   gpc1_1 gpc848 (
      {stage0_12[215]},
      {stage1_12[157]}
   );
   gpc1_1 gpc849 (
      {stage0_12[216]},
      {stage1_12[158]}
   );
   gpc1_1 gpc850 (
      {stage0_12[217]},
      {stage1_12[159]}
   );
   gpc1_1 gpc851 (
      {stage0_12[218]},
      {stage1_12[160]}
   );
   gpc1_1 gpc852 (
      {stage0_12[219]},
      {stage1_12[161]}
   );
   gpc1_1 gpc853 (
      {stage0_12[220]},
      {stage1_12[162]}
   );
   gpc1_1 gpc854 (
      {stage0_12[221]},
      {stage1_12[163]}
   );
   gpc1_1 gpc855 (
      {stage0_12[222]},
      {stage1_12[164]}
   );
   gpc1_1 gpc856 (
      {stage0_12[223]},
      {stage1_12[165]}
   );
   gpc1_1 gpc857 (
      {stage0_12[224]},
      {stage1_12[166]}
   );
   gpc1_1 gpc858 (
      {stage0_12[225]},
      {stage1_12[167]}
   );
   gpc1_1 gpc859 (
      {stage0_12[226]},
      {stage1_12[168]}
   );
   gpc1_1 gpc860 (
      {stage0_12[227]},
      {stage1_12[169]}
   );
   gpc1_1 gpc861 (
      {stage0_12[228]},
      {stage1_12[170]}
   );
   gpc1_1 gpc862 (
      {stage0_12[229]},
      {stage1_12[171]}
   );
   gpc1_1 gpc863 (
      {stage0_12[230]},
      {stage1_12[172]}
   );
   gpc1_1 gpc864 (
      {stage0_12[231]},
      {stage1_12[173]}
   );
   gpc1_1 gpc865 (
      {stage0_12[232]},
      {stage1_12[174]}
   );
   gpc1_1 gpc866 (
      {stage0_12[233]},
      {stage1_12[175]}
   );
   gpc1_1 gpc867 (
      {stage0_12[234]},
      {stage1_12[176]}
   );
   gpc1_1 gpc868 (
      {stage0_12[235]},
      {stage1_12[177]}
   );
   gpc1_1 gpc869 (
      {stage0_12[236]},
      {stage1_12[178]}
   );
   gpc1_1 gpc870 (
      {stage0_12[237]},
      {stage1_12[179]}
   );
   gpc1_1 gpc871 (
      {stage0_12[238]},
      {stage1_12[180]}
   );
   gpc1_1 gpc872 (
      {stage0_12[239]},
      {stage1_12[181]}
   );
   gpc1_1 gpc873 (
      {stage0_12[240]},
      {stage1_12[182]}
   );
   gpc1_1 gpc874 (
      {stage0_12[241]},
      {stage1_12[183]}
   );
   gpc1_1 gpc875 (
      {stage0_12[242]},
      {stage1_12[184]}
   );
   gpc1_1 gpc876 (
      {stage0_12[243]},
      {stage1_12[185]}
   );
   gpc1_1 gpc877 (
      {stage0_12[244]},
      {stage1_12[186]}
   );
   gpc1_1 gpc878 (
      {stage0_12[245]},
      {stage1_12[187]}
   );
   gpc1_1 gpc879 (
      {stage0_12[246]},
      {stage1_12[188]}
   );
   gpc1_1 gpc880 (
      {stage0_12[247]},
      {stage1_12[189]}
   );
   gpc1_1 gpc881 (
      {stage0_12[248]},
      {stage1_12[190]}
   );
   gpc1_1 gpc882 (
      {stage0_12[249]},
      {stage1_12[191]}
   );
   gpc1_1 gpc883 (
      {stage0_12[250]},
      {stage1_12[192]}
   );
   gpc1_1 gpc884 (
      {stage0_12[251]},
      {stage1_12[193]}
   );
   gpc1_1 gpc885 (
      {stage0_12[252]},
      {stage1_12[194]}
   );
   gpc1_1 gpc886 (
      {stage0_12[253]},
      {stage1_12[195]}
   );
   gpc1_1 gpc887 (
      {stage0_12[254]},
      {stage1_12[196]}
   );
   gpc1_1 gpc888 (
      {stage0_12[255]},
      {stage1_12[197]}
   );
   gpc1_1 gpc889 (
      {stage0_14[235]},
      {stage1_14[93]}
   );
   gpc1_1 gpc890 (
      {stage0_14[236]},
      {stage1_14[94]}
   );
   gpc1_1 gpc891 (
      {stage0_14[237]},
      {stage1_14[95]}
   );
   gpc1_1 gpc892 (
      {stage0_14[238]},
      {stage1_14[96]}
   );
   gpc1_1 gpc893 (
      {stage0_14[239]},
      {stage1_14[97]}
   );
   gpc1_1 gpc894 (
      {stage0_14[240]},
      {stage1_14[98]}
   );
   gpc1_1 gpc895 (
      {stage0_14[241]},
      {stage1_14[99]}
   );
   gpc1_1 gpc896 (
      {stage0_14[242]},
      {stage1_14[100]}
   );
   gpc1_1 gpc897 (
      {stage0_14[243]},
      {stage1_14[101]}
   );
   gpc1_1 gpc898 (
      {stage0_14[244]},
      {stage1_14[102]}
   );
   gpc1_1 gpc899 (
      {stage0_14[245]},
      {stage1_14[103]}
   );
   gpc1_1 gpc900 (
      {stage0_14[246]},
      {stage1_14[104]}
   );
   gpc1_1 gpc901 (
      {stage0_14[247]},
      {stage1_14[105]}
   );
   gpc1_1 gpc902 (
      {stage0_14[248]},
      {stage1_14[106]}
   );
   gpc1_1 gpc903 (
      {stage0_14[249]},
      {stage1_14[107]}
   );
   gpc1_1 gpc904 (
      {stage0_14[250]},
      {stage1_14[108]}
   );
   gpc1_1 gpc905 (
      {stage0_14[251]},
      {stage1_14[109]}
   );
   gpc1_1 gpc906 (
      {stage0_14[252]},
      {stage1_14[110]}
   );
   gpc1_1 gpc907 (
      {stage0_14[253]},
      {stage1_14[111]}
   );
   gpc1_1 gpc908 (
      {stage0_14[254]},
      {stage1_14[112]}
   );
   gpc1_1 gpc909 (
      {stage0_14[255]},
      {stage1_14[113]}
   );
   gpc1_1 gpc910 (
      {stage0_15[254]},
      {stage1_15[91]}
   );
   gpc1_1 gpc911 (
      {stage0_15[255]},
      {stage1_15[92]}
   );
   gpc1_1 gpc912 (
      {stage0_17[252]},
      {stage1_17[123]}
   );
   gpc1_1 gpc913 (
      {stage0_17[253]},
      {stage1_17[124]}
   );
   gpc1_1 gpc914 (
      {stage0_17[254]},
      {stage1_17[125]}
   );
   gpc1_1 gpc915 (
      {stage0_17[255]},
      {stage1_17[126]}
   );
   gpc1_1 gpc916 (
      {stage0_18[204]},
      {stage1_18[99]}
   );
   gpc1_1 gpc917 (
      {stage0_18[205]},
      {stage1_18[100]}
   );
   gpc1_1 gpc918 (
      {stage0_18[206]},
      {stage1_18[101]}
   );
   gpc1_1 gpc919 (
      {stage0_18[207]},
      {stage1_18[102]}
   );
   gpc1_1 gpc920 (
      {stage0_18[208]},
      {stage1_18[103]}
   );
   gpc1_1 gpc921 (
      {stage0_18[209]},
      {stage1_18[104]}
   );
   gpc1_1 gpc922 (
      {stage0_18[210]},
      {stage1_18[105]}
   );
   gpc1_1 gpc923 (
      {stage0_18[211]},
      {stage1_18[106]}
   );
   gpc1_1 gpc924 (
      {stage0_18[212]},
      {stage1_18[107]}
   );
   gpc1_1 gpc925 (
      {stage0_18[213]},
      {stage1_18[108]}
   );
   gpc1_1 gpc926 (
      {stage0_18[214]},
      {stage1_18[109]}
   );
   gpc1_1 gpc927 (
      {stage0_18[215]},
      {stage1_18[110]}
   );
   gpc1_1 gpc928 (
      {stage0_18[216]},
      {stage1_18[111]}
   );
   gpc1_1 gpc929 (
      {stage0_18[217]},
      {stage1_18[112]}
   );
   gpc1_1 gpc930 (
      {stage0_18[218]},
      {stage1_18[113]}
   );
   gpc1_1 gpc931 (
      {stage0_18[219]},
      {stage1_18[114]}
   );
   gpc1_1 gpc932 (
      {stage0_18[220]},
      {stage1_18[115]}
   );
   gpc1_1 gpc933 (
      {stage0_18[221]},
      {stage1_18[116]}
   );
   gpc1_1 gpc934 (
      {stage0_18[222]},
      {stage1_18[117]}
   );
   gpc1_1 gpc935 (
      {stage0_18[223]},
      {stage1_18[118]}
   );
   gpc1_1 gpc936 (
      {stage0_18[224]},
      {stage1_18[119]}
   );
   gpc1_1 gpc937 (
      {stage0_18[225]},
      {stage1_18[120]}
   );
   gpc1_1 gpc938 (
      {stage0_18[226]},
      {stage1_18[121]}
   );
   gpc1_1 gpc939 (
      {stage0_18[227]},
      {stage1_18[122]}
   );
   gpc1_1 gpc940 (
      {stage0_18[228]},
      {stage1_18[123]}
   );
   gpc1_1 gpc941 (
      {stage0_18[229]},
      {stage1_18[124]}
   );
   gpc1_1 gpc942 (
      {stage0_18[230]},
      {stage1_18[125]}
   );
   gpc1_1 gpc943 (
      {stage0_18[231]},
      {stage1_18[126]}
   );
   gpc1_1 gpc944 (
      {stage0_18[232]},
      {stage1_18[127]}
   );
   gpc1_1 gpc945 (
      {stage0_18[233]},
      {stage1_18[128]}
   );
   gpc1_1 gpc946 (
      {stage0_18[234]},
      {stage1_18[129]}
   );
   gpc1_1 gpc947 (
      {stage0_18[235]},
      {stage1_18[130]}
   );
   gpc1_1 gpc948 (
      {stage0_18[236]},
      {stage1_18[131]}
   );
   gpc1_1 gpc949 (
      {stage0_18[237]},
      {stage1_18[132]}
   );
   gpc1_1 gpc950 (
      {stage0_18[238]},
      {stage1_18[133]}
   );
   gpc1_1 gpc951 (
      {stage0_18[239]},
      {stage1_18[134]}
   );
   gpc1_1 gpc952 (
      {stage0_18[240]},
      {stage1_18[135]}
   );
   gpc1_1 gpc953 (
      {stage0_18[241]},
      {stage1_18[136]}
   );
   gpc1_1 gpc954 (
      {stage0_18[242]},
      {stage1_18[137]}
   );
   gpc1_1 gpc955 (
      {stage0_18[243]},
      {stage1_18[138]}
   );
   gpc1_1 gpc956 (
      {stage0_18[244]},
      {stage1_18[139]}
   );
   gpc1_1 gpc957 (
      {stage0_18[245]},
      {stage1_18[140]}
   );
   gpc1_1 gpc958 (
      {stage0_18[246]},
      {stage1_18[141]}
   );
   gpc1_1 gpc959 (
      {stage0_18[247]},
      {stage1_18[142]}
   );
   gpc1_1 gpc960 (
      {stage0_18[248]},
      {stage1_18[143]}
   );
   gpc1_1 gpc961 (
      {stage0_18[249]},
      {stage1_18[144]}
   );
   gpc1_1 gpc962 (
      {stage0_18[250]},
      {stage1_18[145]}
   );
   gpc1_1 gpc963 (
      {stage0_18[251]},
      {stage1_18[146]}
   );
   gpc1_1 gpc964 (
      {stage0_18[252]},
      {stage1_18[147]}
   );
   gpc1_1 gpc965 (
      {stage0_18[253]},
      {stage1_18[148]}
   );
   gpc1_1 gpc966 (
      {stage0_18[254]},
      {stage1_18[149]}
   );
   gpc1_1 gpc967 (
      {stage0_18[255]},
      {stage1_18[150]}
   );
   gpc1_1 gpc968 (
      {stage0_19[240]},
      {stage1_19[78]}
   );
   gpc1_1 gpc969 (
      {stage0_19[241]},
      {stage1_19[79]}
   );
   gpc1_1 gpc970 (
      {stage0_19[242]},
      {stage1_19[80]}
   );
   gpc1_1 gpc971 (
      {stage0_19[243]},
      {stage1_19[81]}
   );
   gpc1_1 gpc972 (
      {stage0_19[244]},
      {stage1_19[82]}
   );
   gpc1_1 gpc973 (
      {stage0_19[245]},
      {stage1_19[83]}
   );
   gpc1_1 gpc974 (
      {stage0_19[246]},
      {stage1_19[84]}
   );
   gpc1_1 gpc975 (
      {stage0_19[247]},
      {stage1_19[85]}
   );
   gpc1_1 gpc976 (
      {stage0_19[248]},
      {stage1_19[86]}
   );
   gpc1_1 gpc977 (
      {stage0_19[249]},
      {stage1_19[87]}
   );
   gpc1_1 gpc978 (
      {stage0_19[250]},
      {stage1_19[88]}
   );
   gpc1_1 gpc979 (
      {stage0_19[251]},
      {stage1_19[89]}
   );
   gpc1_1 gpc980 (
      {stage0_19[252]},
      {stage1_19[90]}
   );
   gpc1_1 gpc981 (
      {stage0_19[253]},
      {stage1_19[91]}
   );
   gpc1_1 gpc982 (
      {stage0_19[254]},
      {stage1_19[92]}
   );
   gpc1_1 gpc983 (
      {stage0_19[255]},
      {stage1_19[93]}
   );
   gpc1_1 gpc984 (
      {stage0_20[245]},
      {stage1_20[105]}
   );
   gpc1_1 gpc985 (
      {stage0_20[246]},
      {stage1_20[106]}
   );
   gpc1_1 gpc986 (
      {stage0_20[247]},
      {stage1_20[107]}
   );
   gpc1_1 gpc987 (
      {stage0_20[248]},
      {stage1_20[108]}
   );
   gpc1_1 gpc988 (
      {stage0_20[249]},
      {stage1_20[109]}
   );
   gpc1_1 gpc989 (
      {stage0_20[250]},
      {stage1_20[110]}
   );
   gpc1_1 gpc990 (
      {stage0_20[251]},
      {stage1_20[111]}
   );
   gpc1_1 gpc991 (
      {stage0_20[252]},
      {stage1_20[112]}
   );
   gpc1_1 gpc992 (
      {stage0_20[253]},
      {stage1_20[113]}
   );
   gpc1_1 gpc993 (
      {stage0_20[254]},
      {stage1_20[114]}
   );
   gpc1_1 gpc994 (
      {stage0_20[255]},
      {stage1_20[115]}
   );
   gpc1_1 gpc995 (
      {stage0_21[235]},
      {stage1_21[118]}
   );
   gpc1_1 gpc996 (
      {stage0_21[236]},
      {stage1_21[119]}
   );
   gpc1_1 gpc997 (
      {stage0_21[237]},
      {stage1_21[120]}
   );
   gpc1_1 gpc998 (
      {stage0_21[238]},
      {stage1_21[121]}
   );
   gpc1_1 gpc999 (
      {stage0_21[239]},
      {stage1_21[122]}
   );
   gpc1_1 gpc1000 (
      {stage0_21[240]},
      {stage1_21[123]}
   );
   gpc1_1 gpc1001 (
      {stage0_21[241]},
      {stage1_21[124]}
   );
   gpc1_1 gpc1002 (
      {stage0_21[242]},
      {stage1_21[125]}
   );
   gpc1_1 gpc1003 (
      {stage0_21[243]},
      {stage1_21[126]}
   );
   gpc1_1 gpc1004 (
      {stage0_21[244]},
      {stage1_21[127]}
   );
   gpc1_1 gpc1005 (
      {stage0_21[245]},
      {stage1_21[128]}
   );
   gpc1_1 gpc1006 (
      {stage0_21[246]},
      {stage1_21[129]}
   );
   gpc1_1 gpc1007 (
      {stage0_21[247]},
      {stage1_21[130]}
   );
   gpc1_1 gpc1008 (
      {stage0_21[248]},
      {stage1_21[131]}
   );
   gpc1_1 gpc1009 (
      {stage0_21[249]},
      {stage1_21[132]}
   );
   gpc1_1 gpc1010 (
      {stage0_21[250]},
      {stage1_21[133]}
   );
   gpc1_1 gpc1011 (
      {stage0_21[251]},
      {stage1_21[134]}
   );
   gpc1_1 gpc1012 (
      {stage0_21[252]},
      {stage1_21[135]}
   );
   gpc1_1 gpc1013 (
      {stage0_21[253]},
      {stage1_21[136]}
   );
   gpc1_1 gpc1014 (
      {stage0_21[254]},
      {stage1_21[137]}
   );
   gpc1_1 gpc1015 (
      {stage0_21[255]},
      {stage1_21[138]}
   );
   gpc1_1 gpc1016 (
      {stage0_22[246]},
      {stage1_22[84]}
   );
   gpc1_1 gpc1017 (
      {stage0_22[247]},
      {stage1_22[85]}
   );
   gpc1_1 gpc1018 (
      {stage0_22[248]},
      {stage1_22[86]}
   );
   gpc1_1 gpc1019 (
      {stage0_22[249]},
      {stage1_22[87]}
   );
   gpc1_1 gpc1020 (
      {stage0_22[250]},
      {stage1_22[88]}
   );
   gpc1_1 gpc1021 (
      {stage0_22[251]},
      {stage1_22[89]}
   );
   gpc1_1 gpc1022 (
      {stage0_22[252]},
      {stage1_22[90]}
   );
   gpc1_1 gpc1023 (
      {stage0_22[253]},
      {stage1_22[91]}
   );
   gpc1_1 gpc1024 (
      {stage0_22[254]},
      {stage1_22[92]}
   );
   gpc1_1 gpc1025 (
      {stage0_22[255]},
      {stage1_22[93]}
   );
   gpc1_1 gpc1026 (
      {stage0_23[246]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1027 (
      {stage0_23[247]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1028 (
      {stage0_23[248]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1029 (
      {stage0_23[249]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1030 (
      {stage0_23[250]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1031 (
      {stage0_23[251]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1032 (
      {stage0_23[252]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1033 (
      {stage0_23[253]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1034 (
      {stage0_23[254]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1035 (
      {stage0_23[255]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1036 (
      {stage0_24[96]},
      {stage1_24[94]}
   );
   gpc1_1 gpc1037 (
      {stage0_24[97]},
      {stage1_24[95]}
   );
   gpc1_1 gpc1038 (
      {stage0_24[98]},
      {stage1_24[96]}
   );
   gpc1_1 gpc1039 (
      {stage0_24[99]},
      {stage1_24[97]}
   );
   gpc1_1 gpc1040 (
      {stage0_24[100]},
      {stage1_24[98]}
   );
   gpc1_1 gpc1041 (
      {stage0_24[101]},
      {stage1_24[99]}
   );
   gpc1_1 gpc1042 (
      {stage0_24[102]},
      {stage1_24[100]}
   );
   gpc1_1 gpc1043 (
      {stage0_24[103]},
      {stage1_24[101]}
   );
   gpc1_1 gpc1044 (
      {stage0_24[104]},
      {stage1_24[102]}
   );
   gpc1_1 gpc1045 (
      {stage0_24[105]},
      {stage1_24[103]}
   );
   gpc1_1 gpc1046 (
      {stage0_24[106]},
      {stage1_24[104]}
   );
   gpc1_1 gpc1047 (
      {stage0_24[107]},
      {stage1_24[105]}
   );
   gpc1_1 gpc1048 (
      {stage0_24[108]},
      {stage1_24[106]}
   );
   gpc1_1 gpc1049 (
      {stage0_24[109]},
      {stage1_24[107]}
   );
   gpc1_1 gpc1050 (
      {stage0_24[110]},
      {stage1_24[108]}
   );
   gpc1_1 gpc1051 (
      {stage0_24[111]},
      {stage1_24[109]}
   );
   gpc1_1 gpc1052 (
      {stage0_24[112]},
      {stage1_24[110]}
   );
   gpc1_1 gpc1053 (
      {stage0_24[113]},
      {stage1_24[111]}
   );
   gpc1_1 gpc1054 (
      {stage0_24[114]},
      {stage1_24[112]}
   );
   gpc1_1 gpc1055 (
      {stage0_24[115]},
      {stage1_24[113]}
   );
   gpc1_1 gpc1056 (
      {stage0_24[116]},
      {stage1_24[114]}
   );
   gpc1_1 gpc1057 (
      {stage0_24[117]},
      {stage1_24[115]}
   );
   gpc1_1 gpc1058 (
      {stage0_24[118]},
      {stage1_24[116]}
   );
   gpc1_1 gpc1059 (
      {stage0_24[119]},
      {stage1_24[117]}
   );
   gpc1_1 gpc1060 (
      {stage0_24[120]},
      {stage1_24[118]}
   );
   gpc1_1 gpc1061 (
      {stage0_24[121]},
      {stage1_24[119]}
   );
   gpc1_1 gpc1062 (
      {stage0_24[122]},
      {stage1_24[120]}
   );
   gpc1_1 gpc1063 (
      {stage0_24[123]},
      {stage1_24[121]}
   );
   gpc1_1 gpc1064 (
      {stage0_24[124]},
      {stage1_24[122]}
   );
   gpc1_1 gpc1065 (
      {stage0_24[125]},
      {stage1_24[123]}
   );
   gpc1_1 gpc1066 (
      {stage0_24[126]},
      {stage1_24[124]}
   );
   gpc1_1 gpc1067 (
      {stage0_24[127]},
      {stage1_24[125]}
   );
   gpc1_1 gpc1068 (
      {stage0_24[128]},
      {stage1_24[126]}
   );
   gpc1_1 gpc1069 (
      {stage0_24[129]},
      {stage1_24[127]}
   );
   gpc1_1 gpc1070 (
      {stage0_24[130]},
      {stage1_24[128]}
   );
   gpc1_1 gpc1071 (
      {stage0_24[131]},
      {stage1_24[129]}
   );
   gpc1_1 gpc1072 (
      {stage0_24[132]},
      {stage1_24[130]}
   );
   gpc1_1 gpc1073 (
      {stage0_24[133]},
      {stage1_24[131]}
   );
   gpc1_1 gpc1074 (
      {stage0_24[134]},
      {stage1_24[132]}
   );
   gpc1_1 gpc1075 (
      {stage0_24[135]},
      {stage1_24[133]}
   );
   gpc1_1 gpc1076 (
      {stage0_24[136]},
      {stage1_24[134]}
   );
   gpc1_1 gpc1077 (
      {stage0_24[137]},
      {stage1_24[135]}
   );
   gpc1_1 gpc1078 (
      {stage0_24[138]},
      {stage1_24[136]}
   );
   gpc1_1 gpc1079 (
      {stage0_24[139]},
      {stage1_24[137]}
   );
   gpc1_1 gpc1080 (
      {stage0_24[140]},
      {stage1_24[138]}
   );
   gpc1_1 gpc1081 (
      {stage0_24[141]},
      {stage1_24[139]}
   );
   gpc1_1 gpc1082 (
      {stage0_24[142]},
      {stage1_24[140]}
   );
   gpc1_1 gpc1083 (
      {stage0_24[143]},
      {stage1_24[141]}
   );
   gpc1_1 gpc1084 (
      {stage0_24[144]},
      {stage1_24[142]}
   );
   gpc1_1 gpc1085 (
      {stage0_24[145]},
      {stage1_24[143]}
   );
   gpc1_1 gpc1086 (
      {stage0_24[146]},
      {stage1_24[144]}
   );
   gpc1_1 gpc1087 (
      {stage0_24[147]},
      {stage1_24[145]}
   );
   gpc1_1 gpc1088 (
      {stage0_24[148]},
      {stage1_24[146]}
   );
   gpc1_1 gpc1089 (
      {stage0_24[149]},
      {stage1_24[147]}
   );
   gpc1_1 gpc1090 (
      {stage0_24[150]},
      {stage1_24[148]}
   );
   gpc1_1 gpc1091 (
      {stage0_24[151]},
      {stage1_24[149]}
   );
   gpc1_1 gpc1092 (
      {stage0_24[152]},
      {stage1_24[150]}
   );
   gpc1_1 gpc1093 (
      {stage0_24[153]},
      {stage1_24[151]}
   );
   gpc1_1 gpc1094 (
      {stage0_24[154]},
      {stage1_24[152]}
   );
   gpc1_1 gpc1095 (
      {stage0_24[155]},
      {stage1_24[153]}
   );
   gpc1_1 gpc1096 (
      {stage0_24[156]},
      {stage1_24[154]}
   );
   gpc1_1 gpc1097 (
      {stage0_24[157]},
      {stage1_24[155]}
   );
   gpc1_1 gpc1098 (
      {stage0_24[158]},
      {stage1_24[156]}
   );
   gpc1_1 gpc1099 (
      {stage0_24[159]},
      {stage1_24[157]}
   );
   gpc1_1 gpc1100 (
      {stage0_24[160]},
      {stage1_24[158]}
   );
   gpc1_1 gpc1101 (
      {stage0_24[161]},
      {stage1_24[159]}
   );
   gpc1_1 gpc1102 (
      {stage0_24[162]},
      {stage1_24[160]}
   );
   gpc1_1 gpc1103 (
      {stage0_24[163]},
      {stage1_24[161]}
   );
   gpc1_1 gpc1104 (
      {stage0_24[164]},
      {stage1_24[162]}
   );
   gpc1_1 gpc1105 (
      {stage0_24[165]},
      {stage1_24[163]}
   );
   gpc1_1 gpc1106 (
      {stage0_24[166]},
      {stage1_24[164]}
   );
   gpc1_1 gpc1107 (
      {stage0_24[167]},
      {stage1_24[165]}
   );
   gpc1_1 gpc1108 (
      {stage0_24[168]},
      {stage1_24[166]}
   );
   gpc1_1 gpc1109 (
      {stage0_24[169]},
      {stage1_24[167]}
   );
   gpc1_1 gpc1110 (
      {stage0_24[170]},
      {stage1_24[168]}
   );
   gpc1_1 gpc1111 (
      {stage0_24[171]},
      {stage1_24[169]}
   );
   gpc1_1 gpc1112 (
      {stage0_24[172]},
      {stage1_24[170]}
   );
   gpc1_1 gpc1113 (
      {stage0_24[173]},
      {stage1_24[171]}
   );
   gpc1_1 gpc1114 (
      {stage0_24[174]},
      {stage1_24[172]}
   );
   gpc1_1 gpc1115 (
      {stage0_24[175]},
      {stage1_24[173]}
   );
   gpc1_1 gpc1116 (
      {stage0_24[176]},
      {stage1_24[174]}
   );
   gpc1_1 gpc1117 (
      {stage0_24[177]},
      {stage1_24[175]}
   );
   gpc1_1 gpc1118 (
      {stage0_24[178]},
      {stage1_24[176]}
   );
   gpc1_1 gpc1119 (
      {stage0_24[179]},
      {stage1_24[177]}
   );
   gpc1_1 gpc1120 (
      {stage0_24[180]},
      {stage1_24[178]}
   );
   gpc1_1 gpc1121 (
      {stage0_24[181]},
      {stage1_24[179]}
   );
   gpc1_1 gpc1122 (
      {stage0_24[182]},
      {stage1_24[180]}
   );
   gpc1_1 gpc1123 (
      {stage0_24[183]},
      {stage1_24[181]}
   );
   gpc1_1 gpc1124 (
      {stage0_24[184]},
      {stage1_24[182]}
   );
   gpc1_1 gpc1125 (
      {stage0_24[185]},
      {stage1_24[183]}
   );
   gpc1_1 gpc1126 (
      {stage0_24[186]},
      {stage1_24[184]}
   );
   gpc1_1 gpc1127 (
      {stage0_24[187]},
      {stage1_24[185]}
   );
   gpc1_1 gpc1128 (
      {stage0_24[188]},
      {stage1_24[186]}
   );
   gpc1_1 gpc1129 (
      {stage0_24[189]},
      {stage1_24[187]}
   );
   gpc1_1 gpc1130 (
      {stage0_24[190]},
      {stage1_24[188]}
   );
   gpc1_1 gpc1131 (
      {stage0_24[191]},
      {stage1_24[189]}
   );
   gpc1_1 gpc1132 (
      {stage0_24[192]},
      {stage1_24[190]}
   );
   gpc1_1 gpc1133 (
      {stage0_24[193]},
      {stage1_24[191]}
   );
   gpc1_1 gpc1134 (
      {stage0_24[194]},
      {stage1_24[192]}
   );
   gpc1_1 gpc1135 (
      {stage0_24[195]},
      {stage1_24[193]}
   );
   gpc1_1 gpc1136 (
      {stage0_24[196]},
      {stage1_24[194]}
   );
   gpc1_1 gpc1137 (
      {stage0_24[197]},
      {stage1_24[195]}
   );
   gpc1_1 gpc1138 (
      {stage0_24[198]},
      {stage1_24[196]}
   );
   gpc1_1 gpc1139 (
      {stage0_24[199]},
      {stage1_24[197]}
   );
   gpc1_1 gpc1140 (
      {stage0_24[200]},
      {stage1_24[198]}
   );
   gpc1_1 gpc1141 (
      {stage0_24[201]},
      {stage1_24[199]}
   );
   gpc1_1 gpc1142 (
      {stage0_24[202]},
      {stage1_24[200]}
   );
   gpc1_1 gpc1143 (
      {stage0_24[203]},
      {stage1_24[201]}
   );
   gpc1_1 gpc1144 (
      {stage0_24[204]},
      {stage1_24[202]}
   );
   gpc1_1 gpc1145 (
      {stage0_24[205]},
      {stage1_24[203]}
   );
   gpc1_1 gpc1146 (
      {stage0_24[206]},
      {stage1_24[204]}
   );
   gpc1_1 gpc1147 (
      {stage0_24[207]},
      {stage1_24[205]}
   );
   gpc1_1 gpc1148 (
      {stage0_24[208]},
      {stage1_24[206]}
   );
   gpc1_1 gpc1149 (
      {stage0_24[209]},
      {stage1_24[207]}
   );
   gpc1_1 gpc1150 (
      {stage0_24[210]},
      {stage1_24[208]}
   );
   gpc1_1 gpc1151 (
      {stage0_24[211]},
      {stage1_24[209]}
   );
   gpc1_1 gpc1152 (
      {stage0_24[212]},
      {stage1_24[210]}
   );
   gpc1_1 gpc1153 (
      {stage0_24[213]},
      {stage1_24[211]}
   );
   gpc1_1 gpc1154 (
      {stage0_24[214]},
      {stage1_24[212]}
   );
   gpc1_1 gpc1155 (
      {stage0_24[215]},
      {stage1_24[213]}
   );
   gpc1_1 gpc1156 (
      {stage0_24[216]},
      {stage1_24[214]}
   );
   gpc1_1 gpc1157 (
      {stage0_24[217]},
      {stage1_24[215]}
   );
   gpc1_1 gpc1158 (
      {stage0_24[218]},
      {stage1_24[216]}
   );
   gpc1_1 gpc1159 (
      {stage0_24[219]},
      {stage1_24[217]}
   );
   gpc1_1 gpc1160 (
      {stage0_24[220]},
      {stage1_24[218]}
   );
   gpc1_1 gpc1161 (
      {stage0_24[221]},
      {stage1_24[219]}
   );
   gpc1_1 gpc1162 (
      {stage0_24[222]},
      {stage1_24[220]}
   );
   gpc1_1 gpc1163 (
      {stage0_24[223]},
      {stage1_24[221]}
   );
   gpc1_1 gpc1164 (
      {stage0_24[224]},
      {stage1_24[222]}
   );
   gpc1_1 gpc1165 (
      {stage0_24[225]},
      {stage1_24[223]}
   );
   gpc1_1 gpc1166 (
      {stage0_24[226]},
      {stage1_24[224]}
   );
   gpc1_1 gpc1167 (
      {stage0_24[227]},
      {stage1_24[225]}
   );
   gpc1_1 gpc1168 (
      {stage0_24[228]},
      {stage1_24[226]}
   );
   gpc1_1 gpc1169 (
      {stage0_24[229]},
      {stage1_24[227]}
   );
   gpc1_1 gpc1170 (
      {stage0_24[230]},
      {stage1_24[228]}
   );
   gpc1_1 gpc1171 (
      {stage0_24[231]},
      {stage1_24[229]}
   );
   gpc1_1 gpc1172 (
      {stage0_24[232]},
      {stage1_24[230]}
   );
   gpc1_1 gpc1173 (
      {stage0_24[233]},
      {stage1_24[231]}
   );
   gpc1_1 gpc1174 (
      {stage0_24[234]},
      {stage1_24[232]}
   );
   gpc1_1 gpc1175 (
      {stage0_24[235]},
      {stage1_24[233]}
   );
   gpc1_1 gpc1176 (
      {stage0_24[236]},
      {stage1_24[234]}
   );
   gpc1_1 gpc1177 (
      {stage0_24[237]},
      {stage1_24[235]}
   );
   gpc1_1 gpc1178 (
      {stage0_24[238]},
      {stage1_24[236]}
   );
   gpc1_1 gpc1179 (
      {stage0_24[239]},
      {stage1_24[237]}
   );
   gpc1_1 gpc1180 (
      {stage0_24[240]},
      {stage1_24[238]}
   );
   gpc1_1 gpc1181 (
      {stage0_24[241]},
      {stage1_24[239]}
   );
   gpc1_1 gpc1182 (
      {stage0_24[242]},
      {stage1_24[240]}
   );
   gpc1_1 gpc1183 (
      {stage0_24[243]},
      {stage1_24[241]}
   );
   gpc1_1 gpc1184 (
      {stage0_24[244]},
      {stage1_24[242]}
   );
   gpc1_1 gpc1185 (
      {stage0_24[245]},
      {stage1_24[243]}
   );
   gpc1_1 gpc1186 (
      {stage0_24[246]},
      {stage1_24[244]}
   );
   gpc1_1 gpc1187 (
      {stage0_24[247]},
      {stage1_24[245]}
   );
   gpc1_1 gpc1188 (
      {stage0_24[248]},
      {stage1_24[246]}
   );
   gpc1_1 gpc1189 (
      {stage0_24[249]},
      {stage1_24[247]}
   );
   gpc1_1 gpc1190 (
      {stage0_24[250]},
      {stage1_24[248]}
   );
   gpc1_1 gpc1191 (
      {stage0_24[251]},
      {stage1_24[249]}
   );
   gpc1_1 gpc1192 (
      {stage0_24[252]},
      {stage1_24[250]}
   );
   gpc1_1 gpc1193 (
      {stage0_24[253]},
      {stage1_24[251]}
   );
   gpc1_1 gpc1194 (
      {stage0_24[254]},
      {stage1_24[252]}
   );
   gpc1_1 gpc1195 (
      {stage0_24[255]},
      {stage1_24[253]}
   );
   gpc1_1 gpc1196 (
      {stage0_25[222]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1197 (
      {stage0_25[223]},
      {stage1_25[85]}
   );
   gpc1_1 gpc1198 (
      {stage0_25[224]},
      {stage1_25[86]}
   );
   gpc1_1 gpc1199 (
      {stage0_25[225]},
      {stage1_25[87]}
   );
   gpc1_1 gpc1200 (
      {stage0_25[226]},
      {stage1_25[88]}
   );
   gpc1_1 gpc1201 (
      {stage0_25[227]},
      {stage1_25[89]}
   );
   gpc1_1 gpc1202 (
      {stage0_25[228]},
      {stage1_25[90]}
   );
   gpc1_1 gpc1203 (
      {stage0_25[229]},
      {stage1_25[91]}
   );
   gpc1_1 gpc1204 (
      {stage0_25[230]},
      {stage1_25[92]}
   );
   gpc1_1 gpc1205 (
      {stage0_25[231]},
      {stage1_25[93]}
   );
   gpc1_1 gpc1206 (
      {stage0_25[232]},
      {stage1_25[94]}
   );
   gpc1_1 gpc1207 (
      {stage0_25[233]},
      {stage1_25[95]}
   );
   gpc1_1 gpc1208 (
      {stage0_25[234]},
      {stage1_25[96]}
   );
   gpc1_1 gpc1209 (
      {stage0_25[235]},
      {stage1_25[97]}
   );
   gpc1_1 gpc1210 (
      {stage0_25[236]},
      {stage1_25[98]}
   );
   gpc1_1 gpc1211 (
      {stage0_25[237]},
      {stage1_25[99]}
   );
   gpc1_1 gpc1212 (
      {stage0_25[238]},
      {stage1_25[100]}
   );
   gpc1_1 gpc1213 (
      {stage0_25[239]},
      {stage1_25[101]}
   );
   gpc1_1 gpc1214 (
      {stage0_25[240]},
      {stage1_25[102]}
   );
   gpc1_1 gpc1215 (
      {stage0_25[241]},
      {stage1_25[103]}
   );
   gpc1_1 gpc1216 (
      {stage0_25[242]},
      {stage1_25[104]}
   );
   gpc1_1 gpc1217 (
      {stage0_25[243]},
      {stage1_25[105]}
   );
   gpc1_1 gpc1218 (
      {stage0_25[244]},
      {stage1_25[106]}
   );
   gpc1_1 gpc1219 (
      {stage0_25[245]},
      {stage1_25[107]}
   );
   gpc1_1 gpc1220 (
      {stage0_25[246]},
      {stage1_25[108]}
   );
   gpc1_1 gpc1221 (
      {stage0_25[247]},
      {stage1_25[109]}
   );
   gpc1_1 gpc1222 (
      {stage0_25[248]},
      {stage1_25[110]}
   );
   gpc1_1 gpc1223 (
      {stage0_25[249]},
      {stage1_25[111]}
   );
   gpc1_1 gpc1224 (
      {stage0_25[250]},
      {stage1_25[112]}
   );
   gpc1_1 gpc1225 (
      {stage0_25[251]},
      {stage1_25[113]}
   );
   gpc1_1 gpc1226 (
      {stage0_25[252]},
      {stage1_25[114]}
   );
   gpc1_1 gpc1227 (
      {stage0_25[253]},
      {stage1_25[115]}
   );
   gpc1_1 gpc1228 (
      {stage0_25[254]},
      {stage1_25[116]}
   );
   gpc1_1 gpc1229 (
      {stage0_25[255]},
      {stage1_25[117]}
   );
   gpc1_1 gpc1230 (
      {stage0_26[72]},
      {stage1_26[53]}
   );
   gpc1_1 gpc1231 (
      {stage0_26[73]},
      {stage1_26[54]}
   );
   gpc1_1 gpc1232 (
      {stage0_26[74]},
      {stage1_26[55]}
   );
   gpc1_1 gpc1233 (
      {stage0_26[75]},
      {stage1_26[56]}
   );
   gpc1_1 gpc1234 (
      {stage0_26[76]},
      {stage1_26[57]}
   );
   gpc1_1 gpc1235 (
      {stage0_26[77]},
      {stage1_26[58]}
   );
   gpc1_1 gpc1236 (
      {stage0_26[78]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1237 (
      {stage0_26[79]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1238 (
      {stage0_26[80]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1239 (
      {stage0_26[81]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1240 (
      {stage0_26[82]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1241 (
      {stage0_26[83]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1242 (
      {stage0_26[84]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1243 (
      {stage0_26[85]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1244 (
      {stage0_26[86]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1245 (
      {stage0_26[87]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1246 (
      {stage0_26[88]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1247 (
      {stage0_26[89]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1248 (
      {stage0_26[90]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1249 (
      {stage0_26[91]},
      {stage1_26[72]}
   );
   gpc1_1 gpc1250 (
      {stage0_26[92]},
      {stage1_26[73]}
   );
   gpc1_1 gpc1251 (
      {stage0_26[93]},
      {stage1_26[74]}
   );
   gpc1_1 gpc1252 (
      {stage0_26[94]},
      {stage1_26[75]}
   );
   gpc1_1 gpc1253 (
      {stage0_26[95]},
      {stage1_26[76]}
   );
   gpc1_1 gpc1254 (
      {stage0_26[96]},
      {stage1_26[77]}
   );
   gpc1_1 gpc1255 (
      {stage0_26[97]},
      {stage1_26[78]}
   );
   gpc1_1 gpc1256 (
      {stage0_26[98]},
      {stage1_26[79]}
   );
   gpc1_1 gpc1257 (
      {stage0_26[99]},
      {stage1_26[80]}
   );
   gpc1_1 gpc1258 (
      {stage0_26[100]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1259 (
      {stage0_26[101]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1260 (
      {stage0_26[102]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1261 (
      {stage0_26[103]},
      {stage1_26[84]}
   );
   gpc1_1 gpc1262 (
      {stage0_26[104]},
      {stage1_26[85]}
   );
   gpc1_1 gpc1263 (
      {stage0_26[105]},
      {stage1_26[86]}
   );
   gpc1_1 gpc1264 (
      {stage0_26[106]},
      {stage1_26[87]}
   );
   gpc1_1 gpc1265 (
      {stage0_26[107]},
      {stage1_26[88]}
   );
   gpc1_1 gpc1266 (
      {stage0_26[108]},
      {stage1_26[89]}
   );
   gpc1_1 gpc1267 (
      {stage0_26[109]},
      {stage1_26[90]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[110]},
      {stage1_26[91]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[111]},
      {stage1_26[92]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[112]},
      {stage1_26[93]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[113]},
      {stage1_26[94]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[114]},
      {stage1_26[95]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[115]},
      {stage1_26[96]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[116]},
      {stage1_26[97]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[117]},
      {stage1_26[98]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[118]},
      {stage1_26[99]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[119]},
      {stage1_26[100]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[120]},
      {stage1_26[101]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[121]},
      {stage1_26[102]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[122]},
      {stage1_26[103]}
   );
   gpc1_1 gpc1281 (
      {stage0_26[123]},
      {stage1_26[104]}
   );
   gpc1_1 gpc1282 (
      {stage0_26[124]},
      {stage1_26[105]}
   );
   gpc1_1 gpc1283 (
      {stage0_26[125]},
      {stage1_26[106]}
   );
   gpc1_1 gpc1284 (
      {stage0_26[126]},
      {stage1_26[107]}
   );
   gpc1_1 gpc1285 (
      {stage0_26[127]},
      {stage1_26[108]}
   );
   gpc1_1 gpc1286 (
      {stage0_26[128]},
      {stage1_26[109]}
   );
   gpc1_1 gpc1287 (
      {stage0_26[129]},
      {stage1_26[110]}
   );
   gpc1_1 gpc1288 (
      {stage0_26[130]},
      {stage1_26[111]}
   );
   gpc1_1 gpc1289 (
      {stage0_26[131]},
      {stage1_26[112]}
   );
   gpc1_1 gpc1290 (
      {stage0_26[132]},
      {stage1_26[113]}
   );
   gpc1_1 gpc1291 (
      {stage0_26[133]},
      {stage1_26[114]}
   );
   gpc1_1 gpc1292 (
      {stage0_26[134]},
      {stage1_26[115]}
   );
   gpc1_1 gpc1293 (
      {stage0_26[135]},
      {stage1_26[116]}
   );
   gpc1_1 gpc1294 (
      {stage0_26[136]},
      {stage1_26[117]}
   );
   gpc1_1 gpc1295 (
      {stage0_26[137]},
      {stage1_26[118]}
   );
   gpc1_1 gpc1296 (
      {stage0_26[138]},
      {stage1_26[119]}
   );
   gpc1_1 gpc1297 (
      {stage0_26[139]},
      {stage1_26[120]}
   );
   gpc1_1 gpc1298 (
      {stage0_26[140]},
      {stage1_26[121]}
   );
   gpc1_1 gpc1299 (
      {stage0_26[141]},
      {stage1_26[122]}
   );
   gpc1_1 gpc1300 (
      {stage0_26[142]},
      {stage1_26[123]}
   );
   gpc1_1 gpc1301 (
      {stage0_26[143]},
      {stage1_26[124]}
   );
   gpc1_1 gpc1302 (
      {stage0_26[144]},
      {stage1_26[125]}
   );
   gpc1_1 gpc1303 (
      {stage0_26[145]},
      {stage1_26[126]}
   );
   gpc1_1 gpc1304 (
      {stage0_26[146]},
      {stage1_26[127]}
   );
   gpc1_1 gpc1305 (
      {stage0_26[147]},
      {stage1_26[128]}
   );
   gpc1_1 gpc1306 (
      {stage0_26[148]},
      {stage1_26[129]}
   );
   gpc1_1 gpc1307 (
      {stage0_26[149]},
      {stage1_26[130]}
   );
   gpc1_1 gpc1308 (
      {stage0_26[150]},
      {stage1_26[131]}
   );
   gpc1_1 gpc1309 (
      {stage0_26[151]},
      {stage1_26[132]}
   );
   gpc1_1 gpc1310 (
      {stage0_26[152]},
      {stage1_26[133]}
   );
   gpc1_1 gpc1311 (
      {stage0_26[153]},
      {stage1_26[134]}
   );
   gpc1_1 gpc1312 (
      {stage0_26[154]},
      {stage1_26[135]}
   );
   gpc1_1 gpc1313 (
      {stage0_26[155]},
      {stage1_26[136]}
   );
   gpc1_1 gpc1314 (
      {stage0_26[156]},
      {stage1_26[137]}
   );
   gpc1_1 gpc1315 (
      {stage0_26[157]},
      {stage1_26[138]}
   );
   gpc1_1 gpc1316 (
      {stage0_26[158]},
      {stage1_26[139]}
   );
   gpc1_1 gpc1317 (
      {stage0_26[159]},
      {stage1_26[140]}
   );
   gpc1_1 gpc1318 (
      {stage0_26[160]},
      {stage1_26[141]}
   );
   gpc1_1 gpc1319 (
      {stage0_26[161]},
      {stage1_26[142]}
   );
   gpc1_1 gpc1320 (
      {stage0_26[162]},
      {stage1_26[143]}
   );
   gpc1_1 gpc1321 (
      {stage0_26[163]},
      {stage1_26[144]}
   );
   gpc1_1 gpc1322 (
      {stage0_26[164]},
      {stage1_26[145]}
   );
   gpc1_1 gpc1323 (
      {stage0_26[165]},
      {stage1_26[146]}
   );
   gpc1_1 gpc1324 (
      {stage0_26[166]},
      {stage1_26[147]}
   );
   gpc1_1 gpc1325 (
      {stage0_26[167]},
      {stage1_26[148]}
   );
   gpc1_1 gpc1326 (
      {stage0_26[168]},
      {stage1_26[149]}
   );
   gpc1_1 gpc1327 (
      {stage0_26[169]},
      {stage1_26[150]}
   );
   gpc1_1 gpc1328 (
      {stage0_26[170]},
      {stage1_26[151]}
   );
   gpc1_1 gpc1329 (
      {stage0_26[171]},
      {stage1_26[152]}
   );
   gpc1_1 gpc1330 (
      {stage0_26[172]},
      {stage1_26[153]}
   );
   gpc1_1 gpc1331 (
      {stage0_26[173]},
      {stage1_26[154]}
   );
   gpc1_1 gpc1332 (
      {stage0_26[174]},
      {stage1_26[155]}
   );
   gpc1_1 gpc1333 (
      {stage0_26[175]},
      {stage1_26[156]}
   );
   gpc1_1 gpc1334 (
      {stage0_26[176]},
      {stage1_26[157]}
   );
   gpc1_1 gpc1335 (
      {stage0_26[177]},
      {stage1_26[158]}
   );
   gpc1_1 gpc1336 (
      {stage0_26[178]},
      {stage1_26[159]}
   );
   gpc1_1 gpc1337 (
      {stage0_26[179]},
      {stage1_26[160]}
   );
   gpc1_1 gpc1338 (
      {stage0_26[180]},
      {stage1_26[161]}
   );
   gpc1_1 gpc1339 (
      {stage0_26[181]},
      {stage1_26[162]}
   );
   gpc1_1 gpc1340 (
      {stage0_26[182]},
      {stage1_26[163]}
   );
   gpc1_1 gpc1341 (
      {stage0_26[183]},
      {stage1_26[164]}
   );
   gpc1_1 gpc1342 (
      {stage0_26[184]},
      {stage1_26[165]}
   );
   gpc1_1 gpc1343 (
      {stage0_26[185]},
      {stage1_26[166]}
   );
   gpc1_1 gpc1344 (
      {stage0_26[186]},
      {stage1_26[167]}
   );
   gpc1_1 gpc1345 (
      {stage0_26[187]},
      {stage1_26[168]}
   );
   gpc1_1 gpc1346 (
      {stage0_26[188]},
      {stage1_26[169]}
   );
   gpc1_1 gpc1347 (
      {stage0_26[189]},
      {stage1_26[170]}
   );
   gpc1_1 gpc1348 (
      {stage0_26[190]},
      {stage1_26[171]}
   );
   gpc1_1 gpc1349 (
      {stage0_26[191]},
      {stage1_26[172]}
   );
   gpc1_1 gpc1350 (
      {stage0_26[192]},
      {stage1_26[173]}
   );
   gpc1_1 gpc1351 (
      {stage0_26[193]},
      {stage1_26[174]}
   );
   gpc1_1 gpc1352 (
      {stage0_26[194]},
      {stage1_26[175]}
   );
   gpc1_1 gpc1353 (
      {stage0_26[195]},
      {stage1_26[176]}
   );
   gpc1_1 gpc1354 (
      {stage0_26[196]},
      {stage1_26[177]}
   );
   gpc1_1 gpc1355 (
      {stage0_26[197]},
      {stage1_26[178]}
   );
   gpc1_1 gpc1356 (
      {stage0_26[198]},
      {stage1_26[179]}
   );
   gpc1_1 gpc1357 (
      {stage0_26[199]},
      {stage1_26[180]}
   );
   gpc1_1 gpc1358 (
      {stage0_26[200]},
      {stage1_26[181]}
   );
   gpc1_1 gpc1359 (
      {stage0_26[201]},
      {stage1_26[182]}
   );
   gpc1_1 gpc1360 (
      {stage0_26[202]},
      {stage1_26[183]}
   );
   gpc1_1 gpc1361 (
      {stage0_26[203]},
      {stage1_26[184]}
   );
   gpc1_1 gpc1362 (
      {stage0_26[204]},
      {stage1_26[185]}
   );
   gpc1_1 gpc1363 (
      {stage0_26[205]},
      {stage1_26[186]}
   );
   gpc1_1 gpc1364 (
      {stage0_26[206]},
      {stage1_26[187]}
   );
   gpc1_1 gpc1365 (
      {stage0_26[207]},
      {stage1_26[188]}
   );
   gpc1_1 gpc1366 (
      {stage0_26[208]},
      {stage1_26[189]}
   );
   gpc1_1 gpc1367 (
      {stage0_26[209]},
      {stage1_26[190]}
   );
   gpc1_1 gpc1368 (
      {stage0_26[210]},
      {stage1_26[191]}
   );
   gpc1_1 gpc1369 (
      {stage0_26[211]},
      {stage1_26[192]}
   );
   gpc1_1 gpc1370 (
      {stage0_26[212]},
      {stage1_26[193]}
   );
   gpc1_1 gpc1371 (
      {stage0_26[213]},
      {stage1_26[194]}
   );
   gpc1_1 gpc1372 (
      {stage0_26[214]},
      {stage1_26[195]}
   );
   gpc1_1 gpc1373 (
      {stage0_26[215]},
      {stage1_26[196]}
   );
   gpc1_1 gpc1374 (
      {stage0_26[216]},
      {stage1_26[197]}
   );
   gpc1_1 gpc1375 (
      {stage0_26[217]},
      {stage1_26[198]}
   );
   gpc1_1 gpc1376 (
      {stage0_26[218]},
      {stage1_26[199]}
   );
   gpc1_1 gpc1377 (
      {stage0_26[219]},
      {stage1_26[200]}
   );
   gpc1_1 gpc1378 (
      {stage0_26[220]},
      {stage1_26[201]}
   );
   gpc1_1 gpc1379 (
      {stage0_26[221]},
      {stage1_26[202]}
   );
   gpc1_1 gpc1380 (
      {stage0_26[222]},
      {stage1_26[203]}
   );
   gpc1_1 gpc1381 (
      {stage0_26[223]},
      {stage1_26[204]}
   );
   gpc1_1 gpc1382 (
      {stage0_26[224]},
      {stage1_26[205]}
   );
   gpc1_1 gpc1383 (
      {stage0_26[225]},
      {stage1_26[206]}
   );
   gpc1_1 gpc1384 (
      {stage0_26[226]},
      {stage1_26[207]}
   );
   gpc1_1 gpc1385 (
      {stage0_26[227]},
      {stage1_26[208]}
   );
   gpc1_1 gpc1386 (
      {stage0_26[228]},
      {stage1_26[209]}
   );
   gpc1_1 gpc1387 (
      {stage0_26[229]},
      {stage1_26[210]}
   );
   gpc1_1 gpc1388 (
      {stage0_26[230]},
      {stage1_26[211]}
   );
   gpc1_1 gpc1389 (
      {stage0_26[231]},
      {stage1_26[212]}
   );
   gpc1_1 gpc1390 (
      {stage0_26[232]},
      {stage1_26[213]}
   );
   gpc1_1 gpc1391 (
      {stage0_26[233]},
      {stage1_26[214]}
   );
   gpc1_1 gpc1392 (
      {stage0_26[234]},
      {stage1_26[215]}
   );
   gpc1_1 gpc1393 (
      {stage0_26[235]},
      {stage1_26[216]}
   );
   gpc1_1 gpc1394 (
      {stage0_26[236]},
      {stage1_26[217]}
   );
   gpc1_1 gpc1395 (
      {stage0_26[237]},
      {stage1_26[218]}
   );
   gpc1_1 gpc1396 (
      {stage0_26[238]},
      {stage1_26[219]}
   );
   gpc1_1 gpc1397 (
      {stage0_26[239]},
      {stage1_26[220]}
   );
   gpc1_1 gpc1398 (
      {stage0_26[240]},
      {stage1_26[221]}
   );
   gpc1_1 gpc1399 (
      {stage0_26[241]},
      {stage1_26[222]}
   );
   gpc1_1 gpc1400 (
      {stage0_26[242]},
      {stage1_26[223]}
   );
   gpc1_1 gpc1401 (
      {stage0_26[243]},
      {stage1_26[224]}
   );
   gpc1_1 gpc1402 (
      {stage0_26[244]},
      {stage1_26[225]}
   );
   gpc1_1 gpc1403 (
      {stage0_26[245]},
      {stage1_26[226]}
   );
   gpc1_1 gpc1404 (
      {stage0_26[246]},
      {stage1_26[227]}
   );
   gpc1_1 gpc1405 (
      {stage0_26[247]},
      {stage1_26[228]}
   );
   gpc1_1 gpc1406 (
      {stage0_26[248]},
      {stage1_26[229]}
   );
   gpc1_1 gpc1407 (
      {stage0_26[249]},
      {stage1_26[230]}
   );
   gpc1_1 gpc1408 (
      {stage0_26[250]},
      {stage1_26[231]}
   );
   gpc1_1 gpc1409 (
      {stage0_26[251]},
      {stage1_26[232]}
   );
   gpc1_1 gpc1410 (
      {stage0_26[252]},
      {stage1_26[233]}
   );
   gpc1_1 gpc1411 (
      {stage0_26[253]},
      {stage1_26[234]}
   );
   gpc1_1 gpc1412 (
      {stage0_26[254]},
      {stage1_26[235]}
   );
   gpc1_1 gpc1413 (
      {stage0_26[255]},
      {stage1_26[236]}
   );
   gpc1_1 gpc1414 (
      {stage0_27[204]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1415 (
      {stage0_27[205]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1416 (
      {stage0_27[206]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1417 (
      {stage0_27[207]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1418 (
      {stage0_27[208]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1419 (
      {stage0_27[209]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1420 (
      {stage0_27[210]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1421 (
      {stage0_27[211]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1422 (
      {stage0_27[212]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1423 (
      {stage0_27[213]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1424 (
      {stage0_27[214]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1425 (
      {stage0_27[215]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1426 (
      {stage0_27[216]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1427 (
      {stage0_27[217]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1428 (
      {stage0_27[218]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1429 (
      {stage0_27[219]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1430 (
      {stage0_27[220]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1431 (
      {stage0_27[221]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1432 (
      {stage0_27[222]},
      {stage1_27[74]}
   );
   gpc1_1 gpc1433 (
      {stage0_27[223]},
      {stage1_27[75]}
   );
   gpc1_1 gpc1434 (
      {stage0_27[224]},
      {stage1_27[76]}
   );
   gpc1_1 gpc1435 (
      {stage0_27[225]},
      {stage1_27[77]}
   );
   gpc1_1 gpc1436 (
      {stage0_27[226]},
      {stage1_27[78]}
   );
   gpc1_1 gpc1437 (
      {stage0_27[227]},
      {stage1_27[79]}
   );
   gpc1_1 gpc1438 (
      {stage0_27[228]},
      {stage1_27[80]}
   );
   gpc1_1 gpc1439 (
      {stage0_27[229]},
      {stage1_27[81]}
   );
   gpc1_1 gpc1440 (
      {stage0_27[230]},
      {stage1_27[82]}
   );
   gpc1_1 gpc1441 (
      {stage0_27[231]},
      {stage1_27[83]}
   );
   gpc1_1 gpc1442 (
      {stage0_27[232]},
      {stage1_27[84]}
   );
   gpc1_1 gpc1443 (
      {stage0_27[233]},
      {stage1_27[85]}
   );
   gpc1_1 gpc1444 (
      {stage0_27[234]},
      {stage1_27[86]}
   );
   gpc1_1 gpc1445 (
      {stage0_27[235]},
      {stage1_27[87]}
   );
   gpc1_1 gpc1446 (
      {stage0_27[236]},
      {stage1_27[88]}
   );
   gpc1_1 gpc1447 (
      {stage0_27[237]},
      {stage1_27[89]}
   );
   gpc1_1 gpc1448 (
      {stage0_27[238]},
      {stage1_27[90]}
   );
   gpc1_1 gpc1449 (
      {stage0_27[239]},
      {stage1_27[91]}
   );
   gpc1_1 gpc1450 (
      {stage0_27[240]},
      {stage1_27[92]}
   );
   gpc1_1 gpc1451 (
      {stage0_27[241]},
      {stage1_27[93]}
   );
   gpc1_1 gpc1452 (
      {stage0_27[242]},
      {stage1_27[94]}
   );
   gpc1_1 gpc1453 (
      {stage0_27[243]},
      {stage1_27[95]}
   );
   gpc1_1 gpc1454 (
      {stage0_27[244]},
      {stage1_27[96]}
   );
   gpc1_1 gpc1455 (
      {stage0_27[245]},
      {stage1_27[97]}
   );
   gpc1_1 gpc1456 (
      {stage0_27[246]},
      {stage1_27[98]}
   );
   gpc1_1 gpc1457 (
      {stage0_27[247]},
      {stage1_27[99]}
   );
   gpc1_1 gpc1458 (
      {stage0_27[248]},
      {stage1_27[100]}
   );
   gpc1_1 gpc1459 (
      {stage0_27[249]},
      {stage1_27[101]}
   );
   gpc1_1 gpc1460 (
      {stage0_27[250]},
      {stage1_27[102]}
   );
   gpc1_1 gpc1461 (
      {stage0_27[251]},
      {stage1_27[103]}
   );
   gpc1_1 gpc1462 (
      {stage0_27[252]},
      {stage1_27[104]}
   );
   gpc1_1 gpc1463 (
      {stage0_27[253]},
      {stage1_27[105]}
   );
   gpc1_1 gpc1464 (
      {stage0_27[254]},
      {stage1_27[106]}
   );
   gpc1_1 gpc1465 (
      {stage0_27[255]},
      {stage1_27[107]}
   );
   gpc1_1 gpc1466 (
      {stage0_28[240]},
      {stage1_28[86]}
   );
   gpc1_1 gpc1467 (
      {stage0_28[241]},
      {stage1_28[87]}
   );
   gpc1_1 gpc1468 (
      {stage0_28[242]},
      {stage1_28[88]}
   );
   gpc1_1 gpc1469 (
      {stage0_28[243]},
      {stage1_28[89]}
   );
   gpc1_1 gpc1470 (
      {stage0_28[244]},
      {stage1_28[90]}
   );
   gpc1_1 gpc1471 (
      {stage0_28[245]},
      {stage1_28[91]}
   );
   gpc1_1 gpc1472 (
      {stage0_28[246]},
      {stage1_28[92]}
   );
   gpc1_1 gpc1473 (
      {stage0_28[247]},
      {stage1_28[93]}
   );
   gpc1_1 gpc1474 (
      {stage0_28[248]},
      {stage1_28[94]}
   );
   gpc1_1 gpc1475 (
      {stage0_28[249]},
      {stage1_28[95]}
   );
   gpc1_1 gpc1476 (
      {stage0_28[250]},
      {stage1_28[96]}
   );
   gpc1_1 gpc1477 (
      {stage0_28[251]},
      {stage1_28[97]}
   );
   gpc1_1 gpc1478 (
      {stage0_28[252]},
      {stage1_28[98]}
   );
   gpc1_1 gpc1479 (
      {stage0_28[253]},
      {stage1_28[99]}
   );
   gpc1_1 gpc1480 (
      {stage0_28[254]},
      {stage1_28[100]}
   );
   gpc1_1 gpc1481 (
      {stage0_28[255]},
      {stage1_28[101]}
   );
   gpc1_1 gpc1482 (
      {stage0_29[246]},
      {stage1_29[108]}
   );
   gpc1_1 gpc1483 (
      {stage0_29[247]},
      {stage1_29[109]}
   );
   gpc1_1 gpc1484 (
      {stage0_29[248]},
      {stage1_29[110]}
   );
   gpc1_1 gpc1485 (
      {stage0_29[249]},
      {stage1_29[111]}
   );
   gpc1_1 gpc1486 (
      {stage0_29[250]},
      {stage1_29[112]}
   );
   gpc1_1 gpc1487 (
      {stage0_29[251]},
      {stage1_29[113]}
   );
   gpc1_1 gpc1488 (
      {stage0_29[252]},
      {stage1_29[114]}
   );
   gpc1_1 gpc1489 (
      {stage0_29[253]},
      {stage1_29[115]}
   );
   gpc1_1 gpc1490 (
      {stage0_29[254]},
      {stage1_29[116]}
   );
   gpc1_1 gpc1491 (
      {stage0_29[255]},
      {stage1_29[117]}
   );
   gpc1_1 gpc1492 (
      {stage0_30[240]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1493 (
      {stage0_30[241]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1494 (
      {stage0_30[242]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1495 (
      {stage0_30[243]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1496 (
      {stage0_30[244]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1497 (
      {stage0_30[245]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1498 (
      {stage0_30[246]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1499 (
      {stage0_30[247]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1500 (
      {stage0_30[248]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1501 (
      {stage0_30[249]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1502 (
      {stage0_30[250]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1503 (
      {stage0_30[251]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1504 (
      {stage0_30[252]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1505 (
      {stage0_30[253]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1506 (
      {stage0_30[254]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1507 (
      {stage0_30[255]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1508 (
      {stage0_31[204]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1509 (
      {stage0_31[205]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1510 (
      {stage0_31[206]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1511 (
      {stage0_31[207]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1512 (
      {stage0_31[208]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1513 (
      {stage0_31[209]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1514 (
      {stage0_31[210]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1515 (
      {stage0_31[211]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1516 (
      {stage0_31[212]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1517 (
      {stage0_31[213]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1518 (
      {stage0_31[214]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1519 (
      {stage0_31[215]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1520 (
      {stage0_31[216]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1521 (
      {stage0_31[217]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1522 (
      {stage0_31[218]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1523 (
      {stage0_31[219]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1524 (
      {stage0_31[220]},
      {stage1_31[97]}
   );
   gpc1_1 gpc1525 (
      {stage0_31[221]},
      {stage1_31[98]}
   );
   gpc1_1 gpc1526 (
      {stage0_31[222]},
      {stage1_31[99]}
   );
   gpc1_1 gpc1527 (
      {stage0_31[223]},
      {stage1_31[100]}
   );
   gpc1_1 gpc1528 (
      {stage0_31[224]},
      {stage1_31[101]}
   );
   gpc1_1 gpc1529 (
      {stage0_31[225]},
      {stage1_31[102]}
   );
   gpc1_1 gpc1530 (
      {stage0_31[226]},
      {stage1_31[103]}
   );
   gpc1_1 gpc1531 (
      {stage0_31[227]},
      {stage1_31[104]}
   );
   gpc1_1 gpc1532 (
      {stage0_31[228]},
      {stage1_31[105]}
   );
   gpc1_1 gpc1533 (
      {stage0_31[229]},
      {stage1_31[106]}
   );
   gpc1_1 gpc1534 (
      {stage0_31[230]},
      {stage1_31[107]}
   );
   gpc1_1 gpc1535 (
      {stage0_31[231]},
      {stage1_31[108]}
   );
   gpc1_1 gpc1536 (
      {stage0_31[232]},
      {stage1_31[109]}
   );
   gpc1_1 gpc1537 (
      {stage0_31[233]},
      {stage1_31[110]}
   );
   gpc1_1 gpc1538 (
      {stage0_31[234]},
      {stage1_31[111]}
   );
   gpc1_1 gpc1539 (
      {stage0_31[235]},
      {stage1_31[112]}
   );
   gpc1_1 gpc1540 (
      {stage0_31[236]},
      {stage1_31[113]}
   );
   gpc1_1 gpc1541 (
      {stage0_31[237]},
      {stage1_31[114]}
   );
   gpc1_1 gpc1542 (
      {stage0_31[238]},
      {stage1_31[115]}
   );
   gpc1_1 gpc1543 (
      {stage0_31[239]},
      {stage1_31[116]}
   );
   gpc1_1 gpc1544 (
      {stage0_31[240]},
      {stage1_31[117]}
   );
   gpc1_1 gpc1545 (
      {stage0_31[241]},
      {stage1_31[118]}
   );
   gpc1_1 gpc1546 (
      {stage0_31[242]},
      {stage1_31[119]}
   );
   gpc1_1 gpc1547 (
      {stage0_31[243]},
      {stage1_31[120]}
   );
   gpc1_1 gpc1548 (
      {stage0_31[244]},
      {stage1_31[121]}
   );
   gpc1_1 gpc1549 (
      {stage0_31[245]},
      {stage1_31[122]}
   );
   gpc1_1 gpc1550 (
      {stage0_31[246]},
      {stage1_31[123]}
   );
   gpc1_1 gpc1551 (
      {stage0_31[247]},
      {stage1_31[124]}
   );
   gpc1_1 gpc1552 (
      {stage0_31[248]},
      {stage1_31[125]}
   );
   gpc1_1 gpc1553 (
      {stage0_31[249]},
      {stage1_31[126]}
   );
   gpc1_1 gpc1554 (
      {stage0_31[250]},
      {stage1_31[127]}
   );
   gpc1_1 gpc1555 (
      {stage0_31[251]},
      {stage1_31[128]}
   );
   gpc1_1 gpc1556 (
      {stage0_31[252]},
      {stage1_31[129]}
   );
   gpc1_1 gpc1557 (
      {stage0_31[253]},
      {stage1_31[130]}
   );
   gpc1_1 gpc1558 (
      {stage0_31[254]},
      {stage1_31[131]}
   );
   gpc1_1 gpc1559 (
      {stage0_31[255]},
      {stage1_31[132]}
   );
   gpc1163_5 gpc1560 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1561 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1562 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1563 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1564 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1565 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1566 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1567 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1568 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1569 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1570 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1571 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc1572 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1573 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc1574 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[13]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc1575 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28]},
      {stage1_3[14]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc1576 (
      {stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_3[15]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc1577 (
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage1_3[16]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[17],stage2_2[17]}
   );
   gpc615_5 gpc1578 (
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_3[17]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[18],stage2_2[18]}
   );
   gpc615_5 gpc1579 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage1_3[18]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[19],stage2_2[19]}
   );
   gpc615_5 gpc1580 (
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_3[19]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[20],stage2_2[20]}
   );
   gpc615_5 gpc1581 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58]},
      {stage1_3[20]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[21],stage2_2[21]}
   );
   gpc615_5 gpc1582 (
      {stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage1_3[21]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[22],stage2_2[22]}
   );
   gpc615_5 gpc1583 (
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68]},
      {stage1_3[22]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc1584 (
      {stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73]},
      {stage1_3[23]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc1585 (
      {stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage1_3[24]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc615_5 gpc1586 (
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_3[25]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc1587 (
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[27]}
   );
   gpc615_5 gpc1588 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[84]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[28]}
   );
   gpc615_5 gpc1589 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[85]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[29]}
   );
   gpc615_5 gpc1590 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[86]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[30]}
   );
   gpc615_5 gpc1591 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[87]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[31]}
   );
   gpc615_5 gpc1592 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[88]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[32]}
   );
   gpc615_5 gpc1593 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[89]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[33]}
   );
   gpc615_5 gpc1594 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[90]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[34]}
   );
   gpc615_5 gpc1595 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[91]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[35]}
   );
   gpc615_5 gpc1596 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[92]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[36]}
   );
   gpc615_5 gpc1597 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[93]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[37]}
   );
   gpc615_5 gpc1598 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[94]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[38]}
   );
   gpc207_4 gpc1599 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[12],stage2_6[26],stage2_5[26],stage2_4[39]}
   );
   gpc606_5 gpc1600 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[13],stage2_6[27],stage2_5[27],stage2_4[40]}
   );
   gpc615_5 gpc1601 (
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_5[72]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[14],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc615_5 gpc1602 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117]},
      {stage1_5[73]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[15],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc1603 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[3],stage2_7[16],stage2_6[30],stage2_5[30]}
   );
   gpc606_5 gpc1604 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[4],stage2_7[17],stage2_6[31],stage2_5[31]}
   );
   gpc606_5 gpc1605 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[5],stage2_7[18],stage2_6[32],stage2_5[32]}
   );
   gpc606_5 gpc1606 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[6],stage2_7[19],stage2_6[33],stage2_5[33]}
   );
   gpc606_5 gpc1607 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[7],stage2_7[20],stage2_6[34],stage2_5[34]}
   );
   gpc606_5 gpc1608 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[8],stage2_7[21],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc1609 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[9],stage2_7[22],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc1610 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[10],stage2_7[23],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc1611 (
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[11],stage2_7[24],stage2_6[38]}
   );
   gpc615_5 gpc1612 (
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage1_7[48]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[12],stage2_7[25],stage2_6[39]}
   );
   gpc615_5 gpc1613 (
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_7[49]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[13],stage2_7[26],stage2_6[40]}
   );
   gpc615_5 gpc1614 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[50]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[14],stage2_7[27],stage2_6[41]}
   );
   gpc615_5 gpc1615 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[51]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[15],stage2_7[28],stage2_6[42]}
   );
   gpc615_5 gpc1616 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[52]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[16],stage2_7[29],stage2_6[43]}
   );
   gpc615_5 gpc1617 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[53]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[17],stage2_7[30],stage2_6[44]}
   );
   gpc615_5 gpc1618 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[54]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[18],stage2_7[31],stage2_6[45]}
   );
   gpc615_5 gpc1619 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[55]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[19],stage2_7[32],stage2_6[46]}
   );
   gpc615_5 gpc1620 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[56]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[20],stage2_7[33],stage2_6[47]}
   );
   gpc615_5 gpc1621 (
      {stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75]},
      {stage1_7[57]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[21],stage2_7[34],stage2_6[48]}
   );
   gpc615_5 gpc1622 (
      {stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80]},
      {stage1_7[58]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[22],stage2_7[35],stage2_6[49]}
   );
   gpc615_5 gpc1623 (
      {stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage1_7[59]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[23],stage2_7[36],stage2_6[50]}
   );
   gpc615_5 gpc1624 (
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_7[60]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[24],stage2_7[37],stage2_6[51]}
   );
   gpc615_5 gpc1625 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_7[61]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[25],stage2_7[38],stage2_6[52]}
   );
   gpc615_5 gpc1626 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[90]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[15],stage2_9[23],stage2_8[26],stage2_7[39]}
   );
   gpc615_5 gpc1627 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[91]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[16],stage2_9[24],stage2_8[27],stage2_7[40]}
   );
   gpc615_5 gpc1628 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[92]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[17],stage2_9[25],stage2_8[28],stage2_7[41]}
   );
   gpc615_5 gpc1629 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[93]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[18],stage2_9[26],stage2_8[29],stage2_7[42]}
   );
   gpc615_5 gpc1630 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[94]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[19],stage2_9[27],stage2_8[30],stage2_7[43]}
   );
   gpc615_5 gpc1631 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[95]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[20],stage2_9[28],stage2_8[31],stage2_7[44]}
   );
   gpc606_5 gpc1632 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[6],stage2_10[21],stage2_9[29]}
   );
   gpc606_5 gpc1633 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[1],stage2_11[7],stage2_10[22],stage2_9[30]}
   );
   gpc606_5 gpc1634 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[2],stage2_11[8],stage2_10[23],stage2_9[31]}
   );
   gpc606_5 gpc1635 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[3],stage2_11[9],stage2_10[24],stage2_9[32]}
   );
   gpc606_5 gpc1636 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[4],stage2_11[10],stage2_10[25],stage2_9[33]}
   );
   gpc606_5 gpc1637 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[5],stage2_11[11],stage2_10[26],stage2_9[34]}
   );
   gpc606_5 gpc1638 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[6],stage2_11[12],stage2_10[27],stage2_9[35]}
   );
   gpc606_5 gpc1639 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[7],stage2_11[13],stage2_10[28],stage2_9[36]}
   );
   gpc606_5 gpc1640 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[8],stage2_11[14],stage2_10[29],stage2_9[37]}
   );
   gpc606_5 gpc1641 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[9],stage2_11[15],stage2_10[30],stage2_9[38]}
   );
   gpc606_5 gpc1642 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[10],stage2_11[16],stage2_10[31],stage2_9[39]}
   );
   gpc615_5 gpc1643 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106]},
      {stage1_10[0]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[11],stage2_11[17],stage2_10[32],stage2_9[40]}
   );
   gpc606_5 gpc1644 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[12],stage2_12[12],stage2_11[18],stage2_10[33]}
   );
   gpc606_5 gpc1645 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[13],stage2_12[13],stage2_11[19],stage2_10[34]}
   );
   gpc606_5 gpc1646 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[14],stage2_12[14],stage2_11[20],stage2_10[35]}
   );
   gpc606_5 gpc1647 (
      {stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[15],stage2_12[15],stage2_11[21],stage2_10[36]}
   );
   gpc606_5 gpc1648 (
      {stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[16],stage2_12[16],stage2_11[22],stage2_10[37]}
   );
   gpc606_5 gpc1649 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[17],stage2_12[17],stage2_11[23],stage2_10[38]}
   );
   gpc606_5 gpc1650 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[18],stage2_12[18],stage2_11[24],stage2_10[39]}
   );
   gpc606_5 gpc1651 (
      {stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[19],stage2_12[19],stage2_11[25],stage2_10[40]}
   );
   gpc606_5 gpc1652 (
      {stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[20],stage2_12[20],stage2_11[26],stage2_10[41]}
   );
   gpc606_5 gpc1653 (
      {stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[21],stage2_12[21],stage2_11[27],stage2_10[42]}
   );
   gpc606_5 gpc1654 (
      {stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[22],stage2_12[22],stage2_11[28],stage2_10[43]}
   );
   gpc606_5 gpc1655 (
      {stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[23],stage2_12[23],stage2_11[29],stage2_10[44]}
   );
   gpc606_5 gpc1656 (
      {stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[24],stage2_12[24],stage2_11[30],stage2_10[45]}
   );
   gpc606_5 gpc1657 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[25],stage2_12[25],stage2_11[31],stage2_10[46]}
   );
   gpc606_5 gpc1658 (
      {stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[26],stage2_12[26],stage2_11[32],stage2_10[47]}
   );
   gpc606_5 gpc1659 (
      {stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[27],stage2_12[27],stage2_11[33],stage2_10[48]}
   );
   gpc615_5 gpc1660 (
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76]},
      {stage1_12[96]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[16],stage2_13[28],stage2_12[28],stage2_11[34]}
   );
   gpc615_5 gpc1661 (
      {stage1_11[77], stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81]},
      {stage1_12[97]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[17],stage2_13[29],stage2_12[29],stage2_11[35]}
   );
   gpc615_5 gpc1662 (
      {stage1_11[82], stage1_11[83], stage1_11[84], stage1_11[85], stage1_11[86]},
      {stage1_12[98]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[18],stage2_13[30],stage2_12[30],stage2_11[36]}
   );
   gpc615_5 gpc1663 (
      {stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90], stage1_11[91]},
      {stage1_12[99]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[19],stage2_13[31],stage2_12[31],stage2_11[37]}
   );
   gpc615_5 gpc1664 (
      {stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_12[100]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[20],stage2_13[32],stage2_12[32],stage2_11[38]}
   );
   gpc615_5 gpc1665 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage1_12[101]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[21],stage2_13[33],stage2_12[33],stage2_11[39]}
   );
   gpc615_5 gpc1666 (
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106]},
      {stage1_12[102]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[22],stage2_13[34],stage2_12[34],stage2_11[40]}
   );
   gpc615_5 gpc1667 (
      {stage1_11[107], stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[103]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[23],stage2_13[35],stage2_12[35],stage2_11[41]}
   );
   gpc615_5 gpc1668 (
      {stage1_11[112], stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116]},
      {stage1_12[104]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[24],stage2_13[36],stage2_12[36],stage2_11[42]}
   );
   gpc615_5 gpc1669 (
      {stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121]},
      {stage1_12[105]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[25],stage2_13[37],stage2_12[37],stage2_11[43]}
   );
   gpc615_5 gpc1670 (
      {stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[106]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[26],stage2_13[38],stage2_12[38],stage2_11[44]}
   );
   gpc606_5 gpc1671 (
      {stage1_12[107], stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[11],stage2_14[27],stage2_13[39],stage2_12[39]}
   );
   gpc606_5 gpc1672 (
      {stage1_12[113], stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[12],stage2_14[28],stage2_13[40],stage2_12[40]}
   );
   gpc606_5 gpc1673 (
      {stage1_12[119], stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[13],stage2_14[29],stage2_13[41],stage2_12[41]}
   );
   gpc606_5 gpc1674 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[14],stage2_14[30],stage2_13[42],stage2_12[42]}
   );
   gpc606_5 gpc1675 (
      {stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[15],stage2_14[31],stage2_13[43],stage2_12[43]}
   );
   gpc606_5 gpc1676 (
      {stage1_12[137], stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[16],stage2_14[32],stage2_13[44],stage2_12[44]}
   );
   gpc606_5 gpc1677 (
      {stage1_12[143], stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[17],stage2_14[33],stage2_13[45],stage2_12[45]}
   );
   gpc606_5 gpc1678 (
      {stage1_12[149], stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[18],stage2_14[34],stage2_13[46],stage2_12[46]}
   );
   gpc606_5 gpc1679 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[19],stage2_14[35],stage2_13[47],stage2_12[47]}
   );
   gpc606_5 gpc1680 (
      {stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[20],stage2_14[36],stage2_13[48],stage2_12[48]}
   );
   gpc606_5 gpc1681 (
      {stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[21],stage2_14[37],stage2_13[49],stage2_12[49]}
   );
   gpc606_5 gpc1682 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[11],stage2_15[22],stage2_14[38],stage2_13[50]}
   );
   gpc606_5 gpc1683 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[12],stage2_15[23],stage2_14[39],stage2_13[51]}
   );
   gpc606_5 gpc1684 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[13],stage2_15[24],stage2_14[40],stage2_13[52]}
   );
   gpc606_5 gpc1685 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[14],stage2_15[25],stage2_14[41],stage2_13[53]}
   );
   gpc615_5 gpc1686 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[15],stage2_15[26]}
   );
   gpc615_5 gpc1687 (
      {stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[16],stage2_15[27]}
   );
   gpc615_5 gpc1688 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38]},
      {stage1_16[2]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[17],stage2_15[28]}
   );
   gpc615_5 gpc1689 (
      {stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_16[3]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[3],stage2_17[7],stage2_16[18],stage2_15[29]}
   );
   gpc615_5 gpc1690 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48]},
      {stage1_16[4]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[4],stage2_17[8],stage2_16[19],stage2_15[30]}
   );
   gpc615_5 gpc1691 (
      {stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[5]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[5],stage2_17[9],stage2_16[20],stage2_15[31]}
   );
   gpc615_5 gpc1692 (
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58]},
      {stage1_16[6]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[6],stage2_17[10],stage2_16[21],stage2_15[32]}
   );
   gpc615_5 gpc1693 (
      {stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63]},
      {stage1_16[7]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[7],stage2_17[11],stage2_16[22],stage2_15[33]}
   );
   gpc615_5 gpc1694 (
      {stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67], stage1_15[68]},
      {stage1_16[8]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[8],stage2_17[12],stage2_16[23],stage2_15[34]}
   );
   gpc615_5 gpc1695 (
      {stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_16[9]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[9],stage2_17[13],stage2_16[24],stage2_15[35]}
   );
   gpc615_5 gpc1696 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78]},
      {stage1_16[10]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[10],stage2_17[14],stage2_16[25],stage2_15[36]}
   );
   gpc615_5 gpc1697 (
      {stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[11]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[11],stage2_17[15],stage2_16[26],stage2_15[37]}
   );
   gpc606_5 gpc1698 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[12],stage2_17[16],stage2_16[27]}
   );
   gpc606_5 gpc1699 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[13],stage2_17[17],stage2_16[28]}
   );
   gpc606_5 gpc1700 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[14],stage2_17[18],stage2_16[29]}
   );
   gpc606_5 gpc1701 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[15],stage2_17[19],stage2_16[30]}
   );
   gpc606_5 gpc1702 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[16],stage2_17[20],stage2_16[31]}
   );
   gpc606_5 gpc1703 (
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[17],stage2_18[17],stage2_17[21],stage2_16[32]}
   );
   gpc606_5 gpc1704 (
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[18],stage2_18[18],stage2_17[22],stage2_16[33]}
   );
   gpc606_5 gpc1705 (
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[19],stage2_18[19],stage2_17[23],stage2_16[34]}
   );
   gpc606_5 gpc1706 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[20],stage2_18[20],stage2_17[24],stage2_16[35]}
   );
   gpc606_5 gpc1707 (
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[21],stage2_18[21],stage2_17[25],stage2_16[36]}
   );
   gpc606_5 gpc1708 (
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[22],stage2_18[22],stage2_17[26],stage2_16[37]}
   );
   gpc606_5 gpc1709 (
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[23],stage2_18[23],stage2_17[27],stage2_16[38]}
   );
   gpc606_5 gpc1710 (
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[24],stage2_18[24],stage2_17[28],stage2_16[39]}
   );
   gpc606_5 gpc1711 (
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[25],stage2_18[25],stage2_17[29],stage2_16[40]}
   );
   gpc606_5 gpc1712 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[14],stage2_19[26],stage2_18[26],stage2_17[30]}
   );
   gpc606_5 gpc1713 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[15],stage2_19[27],stage2_18[27],stage2_17[31]}
   );
   gpc606_5 gpc1714 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[16],stage2_19[28],stage2_18[28],stage2_17[32]}
   );
   gpc606_5 gpc1715 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[17],stage2_19[29],stage2_18[29],stage2_17[33]}
   );
   gpc606_5 gpc1716 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[18],stage2_19[30],stage2_18[30],stage2_17[34]}
   );
   gpc606_5 gpc1717 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[19],stage2_19[31],stage2_18[31],stage2_17[35]}
   );
   gpc615_5 gpc1718 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[36]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[20],stage2_19[32],stage2_18[32]}
   );
   gpc615_5 gpc1719 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[21],stage2_19[33],stage2_18[33]}
   );
   gpc615_5 gpc1720 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[12]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[2],stage2_21[8],stage2_20[22],stage2_19[34]}
   );
   gpc615_5 gpc1721 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[13]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[3],stage2_21[9],stage2_20[23],stage2_19[35]}
   );
   gpc615_5 gpc1722 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52]},
      {stage1_20[14]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[4],stage2_21[10],stage2_20[24],stage2_19[36]}
   );
   gpc615_5 gpc1723 (
      {stage1_19[53], stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57]},
      {stage1_20[15]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[5],stage2_21[11],stage2_20[25],stage2_19[37]}
   );
   gpc615_5 gpc1724 (
      {stage1_19[58], stage1_19[59], stage1_19[60], stage1_19[61], stage1_19[62]},
      {stage1_20[16]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[6],stage2_21[12],stage2_20[26],stage2_19[38]}
   );
   gpc615_5 gpc1725 (
      {stage1_19[63], stage1_19[64], stage1_19[65], stage1_19[66], stage1_19[67]},
      {stage1_20[17]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[7],stage2_21[13],stage2_20[27],stage2_19[39]}
   );
   gpc615_5 gpc1726 (
      {stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71], stage1_19[72]},
      {stage1_20[18]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[8],stage2_21[14],stage2_20[28],stage2_19[40]}
   );
   gpc615_5 gpc1727 (
      {stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage1_20[19]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[9],stage2_21[15],stage2_20[29],stage2_19[41]}
   );
   gpc615_5 gpc1728 (
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82]},
      {stage1_20[20]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[10],stage2_21[16],stage2_20[30],stage2_19[42]}
   );
   gpc615_5 gpc1729 (
      {stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_20[21]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[11],stage2_21[17],stage2_20[31],stage2_19[43]}
   );
   gpc615_5 gpc1730 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92]},
      {stage1_20[22]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[12],stage2_21[18],stage2_20[32],stage2_19[44]}
   );
   gpc606_5 gpc1731 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[11],stage2_22[13],stage2_21[19]}
   );
   gpc606_5 gpc1732 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[1],stage2_23[12],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc1733 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[2],stage2_23[13],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc1734 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[3],stage2_23[14],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc1735 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[4],stage2_23[15],stage2_22[17]}
   );
   gpc606_5 gpc1736 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[5],stage2_23[16],stage2_22[18]}
   );
   gpc606_5 gpc1737 (
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[6],stage2_23[17],stage2_22[19]}
   );
   gpc606_5 gpc1738 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[7],stage2_23[18],stage2_22[20]}
   );
   gpc606_5 gpc1739 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[8],stage2_23[19],stage2_22[21]}
   );
   gpc606_5 gpc1740 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[9],stage2_23[20],stage2_22[22]}
   );
   gpc606_5 gpc1741 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[10],stage2_23[21],stage2_22[23]}
   );
   gpc606_5 gpc1742 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[11],stage2_23[22],stage2_22[24]}
   );
   gpc606_5 gpc1743 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[12],stage2_23[23],stage2_22[25]}
   );
   gpc606_5 gpc1744 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[13],stage2_23[24],stage2_22[26]}
   );
   gpc606_5 gpc1745 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[14],stage2_23[25],stage2_22[27]}
   );
   gpc606_5 gpc1746 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[15],stage2_23[26],stage2_22[28]}
   );
   gpc615_5 gpc1747 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76]},
      {stage1_23[24]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[16],stage2_23[27],stage2_22[29]}
   );
   gpc606_5 gpc1748 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29], stage1_23[30]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[13],stage2_25[17],stage2_24[17],stage2_23[28]}
   );
   gpc606_5 gpc1749 (
      {stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[14],stage2_25[18],stage2_24[18],stage2_23[29]}
   );
   gpc606_5 gpc1750 (
      {stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[15],stage2_25[19],stage2_24[19],stage2_23[30]}
   );
   gpc606_5 gpc1751 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[16],stage2_25[20],stage2_24[20],stage2_23[31]}
   );
   gpc606_5 gpc1752 (
      {stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[17],stage2_25[21],stage2_24[21],stage2_23[32]}
   );
   gpc606_5 gpc1753 (
      {stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[18],stage2_25[22],stage2_24[22],stage2_23[33]}
   );
   gpc606_5 gpc1754 (
      {stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[19],stage2_25[23],stage2_24[23],stage2_23[34]}
   );
   gpc606_5 gpc1755 (
      {stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[20],stage2_25[24],stage2_24[24],stage2_23[35]}
   );
   gpc606_5 gpc1756 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[21],stage2_25[25],stage2_24[25]}
   );
   gpc615_5 gpc1757 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88]},
      {stage1_25[48]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[22],stage2_25[26],stage2_24[26]}
   );
   gpc615_5 gpc1758 (
      {stage1_24[89], stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93]},
      {stage1_25[49]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[23],stage2_25[27],stage2_24[27]}
   );
   gpc615_5 gpc1759 (
      {stage1_24[94], stage1_24[95], stage1_24[96], stage1_24[97], stage1_24[98]},
      {stage1_25[50]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[24],stage2_25[28],stage2_24[28]}
   );
   gpc615_5 gpc1760 (
      {stage1_24[99], stage1_24[100], stage1_24[101], stage1_24[102], stage1_24[103]},
      {stage1_25[51]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[12],stage2_26[25],stage2_25[29],stage2_24[29]}
   );
   gpc615_5 gpc1761 (
      {stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107], stage1_24[108]},
      {stage1_25[52]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[13],stage2_26[26],stage2_25[30],stage2_24[30]}
   );
   gpc615_5 gpc1762 (
      {stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_25[53]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[14],stage2_26[27],stage2_25[31],stage2_24[31]}
   );
   gpc615_5 gpc1763 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118]},
      {stage1_25[54]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[15],stage2_26[28],stage2_25[32],stage2_24[32]}
   );
   gpc615_5 gpc1764 (
      {stage1_24[119], stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123]},
      {stage1_25[55]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[16],stage2_26[29],stage2_25[33],stage2_24[33]}
   );
   gpc615_5 gpc1765 (
      {stage1_24[124], stage1_24[125], stage1_24[126], stage1_24[127], stage1_24[128]},
      {stage1_25[56]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[17],stage2_26[30],stage2_25[34],stage2_24[34]}
   );
   gpc615_5 gpc1766 (
      {stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132], stage1_24[133]},
      {stage1_25[57]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[18],stage2_26[31],stage2_25[35],stage2_24[35]}
   );
   gpc615_5 gpc1767 (
      {stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_25[58]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[19],stage2_26[32],stage2_25[36],stage2_24[36]}
   );
   gpc615_5 gpc1768 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_25[59]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[20],stage2_26[33],stage2_25[37],stage2_24[37]}
   );
   gpc615_5 gpc1769 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148]},
      {stage1_25[60]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[21],stage2_26[34],stage2_25[38],stage2_24[38]}
   );
   gpc615_5 gpc1770 (
      {stage1_24[149], stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153]},
      {stage1_25[61]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[22],stage2_26[35],stage2_25[39],stage2_24[39]}
   );
   gpc615_5 gpc1771 (
      {stage1_24[154], stage1_24[155], stage1_24[156], stage1_24[157], stage1_24[158]},
      {stage1_25[62]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[23],stage2_26[36],stage2_25[40],stage2_24[40]}
   );
   gpc615_5 gpc1772 (
      {stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162], stage1_24[163]},
      {stage1_25[63]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[24],stage2_26[37],stage2_25[41],stage2_24[41]}
   );
   gpc615_5 gpc1773 (
      {stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_25[64]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[25],stage2_26[38],stage2_25[42],stage2_24[42]}
   );
   gpc615_5 gpc1774 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[65]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[26],stage2_26[39],stage2_25[43],stage2_24[43]}
   );
   gpc615_5 gpc1775 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[66]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[27],stage2_26[40],stage2_25[44],stage2_24[44]}
   );
   gpc615_5 gpc1776 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[67]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[28],stage2_26[41],stage2_25[45],stage2_24[45]}
   );
   gpc615_5 gpc1777 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[68]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[29],stage2_26[42],stage2_25[46],stage2_24[46]}
   );
   gpc615_5 gpc1778 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[69]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[30],stage2_26[43],stage2_25[47],stage2_24[47]}
   );
   gpc615_5 gpc1779 (
      {stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_25[70]},
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143]},
      {stage2_28[23],stage2_27[31],stage2_26[44],stage2_25[48],stage2_24[48]}
   );
   gpc615_5 gpc1780 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_25[71]},
      {stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage2_28[24],stage2_27[32],stage2_26[45],stage2_25[49],stage2_24[49]}
   );
   gpc615_5 gpc1781 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208]},
      {stage1_25[72]},
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage2_28[25],stage2_27[33],stage2_26[46],stage2_25[50],stage2_24[50]}
   );
   gpc615_5 gpc1782 (
      {stage1_24[209], stage1_24[210], stage1_24[211], stage1_24[212], stage1_24[213]},
      {stage1_25[73]},
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161]},
      {stage2_28[26],stage2_27[34],stage2_26[47],stage2_25[51],stage2_24[51]}
   );
   gpc615_5 gpc1783 (
      {stage1_24[214], stage1_24[215], stage1_24[216], stage1_24[217], stage1_24[218]},
      {stage1_25[74]},
      {stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage2_28[27],stage2_27[35],stage2_26[48],stage2_25[52],stage2_24[52]}
   );
   gpc615_5 gpc1784 (
      {stage1_24[219], stage1_24[220], stage1_24[221], stage1_24[222], stage1_24[223]},
      {stage1_25[75]},
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173]},
      {stage2_28[28],stage2_27[36],stage2_26[49],stage2_25[53],stage2_24[53]}
   );
   gpc615_5 gpc1785 (
      {stage1_24[224], stage1_24[225], stage1_24[226], stage1_24[227], stage1_24[228]},
      {stage1_25[76]},
      {stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage2_28[29],stage2_27[37],stage2_26[50],stage2_25[54],stage2_24[54]}
   );
   gpc615_5 gpc1786 (
      {stage1_24[229], stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233]},
      {stage1_25[77]},
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage2_28[30],stage2_27[38],stage2_26[51],stage2_25[55],stage2_24[55]}
   );
   gpc615_5 gpc1787 (
      {stage1_24[234], stage1_24[235], stage1_24[236], stage1_24[237], stage1_24[238]},
      {stage1_25[78]},
      {stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191]},
      {stage2_28[31],stage2_27[39],stage2_26[52],stage2_25[56],stage2_24[56]}
   );
   gpc615_5 gpc1788 (
      {stage1_24[239], stage1_24[240], stage1_24[241], stage1_24[242], stage1_24[243]},
      {stage1_25[79]},
      {stage1_26[192], stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage2_28[32],stage2_27[40],stage2_26[53],stage2_25[57],stage2_24[57]}
   );
   gpc615_5 gpc1789 (
      {stage1_24[244], stage1_24[245], stage1_24[246], stage1_24[247], stage1_24[248]},
      {stage1_25[80]},
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203]},
      {stage2_28[33],stage2_27[41],stage2_26[54],stage2_25[58],stage2_24[58]}
   );
   gpc606_5 gpc1790 (
      {stage1_25[81], stage1_25[82], stage1_25[83], stage1_25[84], stage1_25[85], stage1_25[86]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[34],stage2_27[42],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc1791 (
      {stage1_25[87], stage1_25[88], stage1_25[89], stage1_25[90], stage1_25[91], stage1_25[92]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[35],stage2_27[43],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc1792 (
      {stage1_25[93], stage1_25[94], stage1_25[95], stage1_25[96], stage1_25[97], stage1_25[98]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[36],stage2_27[44],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc1793 (
      {stage1_25[99], stage1_25[100], stage1_25[101], stage1_25[102], stage1_25[103], stage1_25[104]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[37],stage2_27[45],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc1794 (
      {stage1_25[105], stage1_25[106], stage1_25[107], stage1_25[108], stage1_25[109], stage1_25[110]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[38],stage2_27[46],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc1795 (
      {stage1_25[111], stage1_25[112], stage1_25[113], stage1_25[114], stage1_25[115], stage1_25[116]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[39],stage2_27[47],stage2_26[60],stage2_25[64]}
   );
   gpc615_5 gpc1796 (
      {stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208]},
      {stage1_27[36]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[6],stage2_28[40],stage2_27[48],stage2_26[61]}
   );
   gpc615_5 gpc1797 (
      {stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213]},
      {stage1_27[37]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[7],stage2_28[41],stage2_27[49],stage2_26[62]}
   );
   gpc615_5 gpc1798 (
      {stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217], stage1_26[218]},
      {stage1_27[38]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[8],stage2_28[42],stage2_27[50],stage2_26[63]}
   );
   gpc615_5 gpc1799 (
      {stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222], stage1_26[223]},
      {stage1_27[39]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[9],stage2_28[43],stage2_27[51],stage2_26[64]}
   );
   gpc615_5 gpc1800 (
      {stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227], stage1_26[228]},
      {stage1_27[40]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[10],stage2_28[44],stage2_27[52],stage2_26[65]}
   );
   gpc615_5 gpc1801 (
      {stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232], stage1_26[233]},
      {stage1_27[41]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[11],stage2_28[45],stage2_27[53],stage2_26[66]}
   );
   gpc615_5 gpc1802 (
      {stage1_26[234], stage1_26[235], stage1_26[236], 1'b0, 1'b0},
      {stage1_27[42]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[12],stage2_28[46],stage2_27[54],stage2_26[67]}
   );
   gpc615_5 gpc1803 (
      {stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[13],stage2_28[47],stage2_27[55]}
   );
   gpc615_5 gpc1804 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[14],stage2_28[48],stage2_27[56]}
   );
   gpc615_5 gpc1805 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[44]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[9],stage2_29[15],stage2_28[49],stage2_27[57]}
   );
   gpc615_5 gpc1806 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[45]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[10],stage2_29[16],stage2_28[50],stage2_27[58]}
   );
   gpc615_5 gpc1807 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[46]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[11],stage2_29[17],stage2_28[51],stage2_27[59]}
   );
   gpc615_5 gpc1808 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[47]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[12],stage2_29[18],stage2_28[52],stage2_27[60]}
   );
   gpc606_5 gpc1809 (
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[6],stage2_30[13],stage2_29[19],stage2_28[53]}
   );
   gpc606_5 gpc1810 (
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[7],stage2_30[14],stage2_29[20],stage2_28[54]}
   );
   gpc606_5 gpc1811 (
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[8],stage2_30[15],stage2_29[21],stage2_28[55]}
   );
   gpc606_5 gpc1812 (
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[9],stage2_30[16],stage2_29[22],stage2_28[56]}
   );
   gpc606_5 gpc1813 (
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[10],stage2_30[17],stage2_29[23],stage2_28[57]}
   );
   gpc606_5 gpc1814 (
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[11],stage2_30[18],stage2_29[24],stage2_28[58]}
   );
   gpc606_5 gpc1815 (
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[12],stage2_30[19],stage2_29[25],stage2_28[59]}
   );
   gpc606_5 gpc1816 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[7],stage2_31[13],stage2_30[20],stage2_29[26]}
   );
   gpc606_5 gpc1817 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[8],stage2_31[14],stage2_30[21],stage2_29[27]}
   );
   gpc606_5 gpc1818 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[9],stage2_31[15],stage2_30[22],stage2_29[28]}
   );
   gpc606_5 gpc1819 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[10],stage2_31[16],stage2_30[23],stage2_29[29]}
   );
   gpc606_5 gpc1820 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[11],stage2_31[17],stage2_30[24],stage2_29[30]}
   );
   gpc606_5 gpc1821 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[12],stage2_31[18],stage2_30[25],stage2_29[31]}
   );
   gpc606_5 gpc1822 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[13],stage2_31[19],stage2_30[26],stage2_29[32]}
   );
   gpc606_5 gpc1823 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[14],stage2_31[20],stage2_30[27],stage2_29[33]}
   );
   gpc606_5 gpc1824 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[15],stage2_31[21],stage2_30[28],stage2_29[34]}
   );
   gpc606_5 gpc1825 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[16],stage2_31[22],stage2_30[29],stage2_29[35]}
   );
   gpc606_5 gpc1826 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[17],stage2_31[23],stage2_30[30],stage2_29[36]}
   );
   gpc606_5 gpc1827 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[18],stage2_31[24],stage2_30[31],stage2_29[37]}
   );
   gpc606_5 gpc1828 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[19],stage2_31[25],stage2_30[32],stage2_29[38]}
   );
   gpc606_5 gpc1829 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], 1'b0, 1'b0},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[20],stage2_31[26],stage2_30[33],stage2_29[39]}
   );
   gpc615_5 gpc1830 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46]},
      {stage1_31[84]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[14],stage2_32[21],stage2_31[27],stage2_30[34]}
   );
   gpc615_5 gpc1831 (
      {stage1_30[47], stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51]},
      {stage1_31[85]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[15],stage2_32[22],stage2_31[28],stage2_30[35]}
   );
   gpc615_5 gpc1832 (
      {stage1_30[52], stage1_30[53], stage1_30[54], stage1_30[55], stage1_30[56]},
      {stage1_31[86]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[16],stage2_32[23],stage2_31[29],stage2_30[36]}
   );
   gpc615_5 gpc1833 (
      {stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_31[87]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[17],stage2_32[24],stage2_31[30],stage2_30[37]}
   );
   gpc615_5 gpc1834 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66]},
      {stage1_31[88]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[18],stage2_32[25],stage2_31[31],stage2_30[38]}
   );
   gpc615_5 gpc1835 (
      {stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[19],stage2_32[26],stage2_31[32],stage2_30[39]}
   );
   gpc615_5 gpc1836 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76]},
      {stage1_31[90]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[20],stage2_32[27],stage2_31[33],stage2_30[40]}
   );
   gpc615_5 gpc1837 (
      {stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_31[91]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[21],stage2_32[28],stage2_31[34],stage2_30[41]}
   );
   gpc615_5 gpc1838 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86]},
      {stage1_31[92]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[22],stage2_32[29],stage2_31[35],stage2_30[42]}
   );
   gpc615_5 gpc1839 (
      {stage1_30[87], stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91]},
      {stage1_31[93]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[23],stage2_32[30],stage2_31[36],stage2_30[43]}
   );
   gpc615_5 gpc1840 (
      {stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95], stage1_30[96]},
      {stage1_31[94]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[24],stage2_32[31],stage2_31[37],stage2_30[44]}
   );
   gpc606_5 gpc1841 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[11],stage2_33[25],stage2_32[32],stage2_31[38]}
   );
   gpc606_5 gpc1842 (
      {stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[12],stage2_33[26],stage2_32[33],stage2_31[39]}
   );
   gpc606_5 gpc1843 (
      {stage1_31[107], stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[13],stage2_33[27],stage2_32[34],stage2_31[40]}
   );
   gpc606_5 gpc1844 (
      {stage1_31[113], stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[14],stage2_33[28],stage2_32[35],stage2_31[41]}
   );
   gpc615_5 gpc1845 (
      {stage1_31[119], stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123]},
      {stage1_32[66]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[15],stage2_33[29],stage2_32[36],stage2_31[42]}
   );
   gpc615_5 gpc1846 (
      {stage1_31[124], stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128]},
      {stage1_32[67]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], 1'b0, 1'b0},
      {stage2_35[5],stage2_34[16],stage2_33[30],stage2_32[37],stage2_31[43]}
   );
   gpc1_1 gpc1847 (
      {stage1_0[39]},
      {stage2_0[13]}
   );
   gpc1_1 gpc1848 (
      {stage1_0[40]},
      {stage2_0[14]}
   );
   gpc1_1 gpc1849 (
      {stage1_0[41]},
      {stage2_0[15]}
   );
   gpc1_1 gpc1850 (
      {stage1_0[42]},
      {stage2_0[16]}
   );
   gpc1_1 gpc1851 (
      {stage1_0[43]},
      {stage2_0[17]}
   );
   gpc1_1 gpc1852 (
      {stage1_0[44]},
      {stage2_0[18]}
   );
   gpc1_1 gpc1853 (
      {stage1_0[45]},
      {stage2_0[19]}
   );
   gpc1_1 gpc1854 (
      {stage1_0[46]},
      {stage2_0[20]}
   );
   gpc1_1 gpc1855 (
      {stage1_0[47]},
      {stage2_0[21]}
   );
   gpc1_1 gpc1856 (
      {stage1_0[48]},
      {stage2_0[22]}
   );
   gpc1_1 gpc1857 (
      {stage1_0[49]},
      {stage2_0[23]}
   );
   gpc1_1 gpc1858 (
      {stage1_1[78]},
      {stage2_1[13]}
   );
   gpc1_1 gpc1859 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc1860 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc1861 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc1862 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc1863 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc1864 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc1865 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc1866 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc1867 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc1868 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc1869 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc1870 (
      {stage1_1[90]},
      {stage2_1[25]}
   );
   gpc1_1 gpc1871 (
      {stage1_1[91]},
      {stage2_1[26]}
   );
   gpc1_1 gpc1872 (
      {stage1_1[92]},
      {stage2_1[27]}
   );
   gpc1_1 gpc1873 (
      {stage1_1[93]},
      {stage2_1[28]}
   );
   gpc1_1 gpc1874 (
      {stage1_1[94]},
      {stage2_1[29]}
   );
   gpc1_1 gpc1875 (
      {stage1_1[95]},
      {stage2_1[30]}
   );
   gpc1_1 gpc1876 (
      {stage1_1[96]},
      {stage2_1[31]}
   );
   gpc1_1 gpc1877 (
      {stage1_1[97]},
      {stage2_1[32]}
   );
   gpc1_1 gpc1878 (
      {stage1_2[84]},
      {stage2_2[27]}
   );
   gpc1_1 gpc1879 (
      {stage1_2[85]},
      {stage2_2[28]}
   );
   gpc1_1 gpc1880 (
      {stage1_2[86]},
      {stage2_2[29]}
   );
   gpc1_1 gpc1881 (
      {stage1_2[87]},
      {stage2_2[30]}
   );
   gpc1_1 gpc1882 (
      {stage1_2[88]},
      {stage2_2[31]}
   );
   gpc1_1 gpc1883 (
      {stage1_2[89]},
      {stage2_2[32]}
   );
   gpc1_1 gpc1884 (
      {stage1_2[90]},
      {stage2_2[33]}
   );
   gpc1_1 gpc1885 (
      {stage1_2[91]},
      {stage2_2[34]}
   );
   gpc1_1 gpc1886 (
      {stage1_3[87]},
      {stage2_3[39]}
   );
   gpc1_1 gpc1887 (
      {stage1_3[88]},
      {stage2_3[40]}
   );
   gpc1_1 gpc1888 (
      {stage1_3[89]},
      {stage2_3[41]}
   );
   gpc1_1 gpc1889 (
      {stage1_3[90]},
      {stage2_3[42]}
   );
   gpc1_1 gpc1890 (
      {stage1_4[118]},
      {stage2_4[43]}
   );
   gpc1_1 gpc1891 (
      {stage1_4[119]},
      {stage2_4[44]}
   );
   gpc1_1 gpc1892 (
      {stage1_4[120]},
      {stage2_4[45]}
   );
   gpc1_1 gpc1893 (
      {stage1_4[121]},
      {stage2_4[46]}
   );
   gpc1_1 gpc1894 (
      {stage1_4[122]},
      {stage2_4[47]}
   );
   gpc1_1 gpc1895 (
      {stage1_4[123]},
      {stage2_4[48]}
   );
   gpc1_1 gpc1896 (
      {stage1_4[124]},
      {stage2_4[49]}
   );
   gpc1_1 gpc1897 (
      {stage1_4[125]},
      {stage2_4[50]}
   );
   gpc1_1 gpc1898 (
      {stage1_4[126]},
      {stage2_4[51]}
   );
   gpc1_1 gpc1899 (
      {stage1_4[127]},
      {stage2_4[52]}
   );
   gpc1_1 gpc1900 (
      {stage1_4[128]},
      {stage2_4[53]}
   );
   gpc1_1 gpc1901 (
      {stage1_4[129]},
      {stage2_4[54]}
   );
   gpc1_1 gpc1902 (
      {stage1_4[130]},
      {stage2_4[55]}
   );
   gpc1_1 gpc1903 (
      {stage1_4[131]},
      {stage2_4[56]}
   );
   gpc1_1 gpc1904 (
      {stage1_4[132]},
      {stage2_4[57]}
   );
   gpc1_1 gpc1905 (
      {stage1_4[133]},
      {stage2_4[58]}
   );
   gpc1_1 gpc1906 (
      {stage1_4[134]},
      {stage2_4[59]}
   );
   gpc1_1 gpc1907 (
      {stage1_4[135]},
      {stage2_4[60]}
   );
   gpc1_1 gpc1908 (
      {stage1_4[136]},
      {stage2_4[61]}
   );
   gpc1_1 gpc1909 (
      {stage1_4[137]},
      {stage2_4[62]}
   );
   gpc1_1 gpc1910 (
      {stage1_4[138]},
      {stage2_4[63]}
   );
   gpc1_1 gpc1911 (
      {stage1_4[139]},
      {stage2_4[64]}
   );
   gpc1_1 gpc1912 (
      {stage1_4[140]},
      {stage2_4[65]}
   );
   gpc1_1 gpc1913 (
      {stage1_4[141]},
      {stage2_4[66]}
   );
   gpc1_1 gpc1914 (
      {stage1_4[142]},
      {stage2_4[67]}
   );
   gpc1_1 gpc1915 (
      {stage1_4[143]},
      {stage2_4[68]}
   );
   gpc1_1 gpc1916 (
      {stage1_4[144]},
      {stage2_4[69]}
   );
   gpc1_1 gpc1917 (
      {stage1_4[145]},
      {stage2_4[70]}
   );
   gpc1_1 gpc1918 (
      {stage1_4[146]},
      {stage2_4[71]}
   );
   gpc1_1 gpc1919 (
      {stage1_4[147]},
      {stage2_4[72]}
   );
   gpc1_1 gpc1920 (
      {stage1_4[148]},
      {stage2_4[73]}
   );
   gpc1_1 gpc1921 (
      {stage1_5[122]},
      {stage2_5[38]}
   );
   gpc1_1 gpc1922 (
      {stage1_5[123]},
      {stage2_5[39]}
   );
   gpc1_1 gpc1923 (
      {stage1_5[124]},
      {stage2_5[40]}
   );
   gpc1_1 gpc1924 (
      {stage1_5[125]},
      {stage2_5[41]}
   );
   gpc1_1 gpc1925 (
      {stage1_7[92]},
      {stage2_7[45]}
   );
   gpc1_1 gpc1926 (
      {stage1_7[93]},
      {stage2_7[46]}
   );
   gpc1_1 gpc1927 (
      {stage1_7[94]},
      {stage2_7[47]}
   );
   gpc1_1 gpc1928 (
      {stage1_7[95]},
      {stage2_7[48]}
   );
   gpc1_1 gpc1929 (
      {stage1_7[96]},
      {stage2_7[49]}
   );
   gpc1_1 gpc1930 (
      {stage1_7[97]},
      {stage2_7[50]}
   );
   gpc1_1 gpc1931 (
      {stage1_7[98]},
      {stage2_7[51]}
   );
   gpc1_1 gpc1932 (
      {stage1_7[99]},
      {stage2_7[52]}
   );
   gpc1_1 gpc1933 (
      {stage1_7[100]},
      {stage2_7[53]}
   );
   gpc1_1 gpc1934 (
      {stage1_8[96]},
      {stage2_8[32]}
   );
   gpc1_1 gpc1935 (
      {stage1_8[97]},
      {stage2_8[33]}
   );
   gpc1_1 gpc1936 (
      {stage1_8[98]},
      {stage2_8[34]}
   );
   gpc1_1 gpc1937 (
      {stage1_8[99]},
      {stage2_8[35]}
   );
   gpc1_1 gpc1938 (
      {stage1_8[100]},
      {stage2_8[36]}
   );
   gpc1_1 gpc1939 (
      {stage1_8[101]},
      {stage2_8[37]}
   );
   gpc1_1 gpc1940 (
      {stage1_8[102]},
      {stage2_8[38]}
   );
   gpc1_1 gpc1941 (
      {stage1_8[103]},
      {stage2_8[39]}
   );
   gpc1_1 gpc1942 (
      {stage1_8[104]},
      {stage2_8[40]}
   );
   gpc1_1 gpc1943 (
      {stage1_8[105]},
      {stage2_8[41]}
   );
   gpc1_1 gpc1944 (
      {stage1_8[106]},
      {stage2_8[42]}
   );
   gpc1_1 gpc1945 (
      {stage1_8[107]},
      {stage2_8[43]}
   );
   gpc1_1 gpc1946 (
      {stage1_8[108]},
      {stage2_8[44]}
   );
   gpc1_1 gpc1947 (
      {stage1_8[109]},
      {stage2_8[45]}
   );
   gpc1_1 gpc1948 (
      {stage1_8[110]},
      {stage2_8[46]}
   );
   gpc1_1 gpc1949 (
      {stage1_8[111]},
      {stage2_8[47]}
   );
   gpc1_1 gpc1950 (
      {stage1_8[112]},
      {stage2_8[48]}
   );
   gpc1_1 gpc1951 (
      {stage1_8[113]},
      {stage2_8[49]}
   );
   gpc1_1 gpc1952 (
      {stage1_8[114]},
      {stage2_8[50]}
   );
   gpc1_1 gpc1953 (
      {stage1_8[115]},
      {stage2_8[51]}
   );
   gpc1_1 gpc1954 (
      {stage1_8[116]},
      {stage2_8[52]}
   );
   gpc1_1 gpc1955 (
      {stage1_8[117]},
      {stage2_8[53]}
   );
   gpc1_1 gpc1956 (
      {stage1_8[118]},
      {stage2_8[54]}
   );
   gpc1_1 gpc1957 (
      {stage1_8[119]},
      {stage2_8[55]}
   );
   gpc1_1 gpc1958 (
      {stage1_9[107]},
      {stage2_9[41]}
   );
   gpc1_1 gpc1959 (
      {stage1_9[108]},
      {stage2_9[42]}
   );
   gpc1_1 gpc1960 (
      {stage1_9[109]},
      {stage2_9[43]}
   );
   gpc1_1 gpc1961 (
      {stage1_9[110]},
      {stage2_9[44]}
   );
   gpc1_1 gpc1962 (
      {stage1_9[111]},
      {stage2_9[45]}
   );
   gpc1_1 gpc1963 (
      {stage1_9[112]},
      {stage2_9[46]}
   );
   gpc1_1 gpc1964 (
      {stage1_9[113]},
      {stage2_9[47]}
   );
   gpc1_1 gpc1965 (
      {stage1_9[114]},
      {stage2_9[48]}
   );
   gpc1_1 gpc1966 (
      {stage1_9[115]},
      {stage2_9[49]}
   );
   gpc1_1 gpc1967 (
      {stage1_9[116]},
      {stage2_9[50]}
   );
   gpc1_1 gpc1968 (
      {stage1_9[117]},
      {stage2_9[51]}
   );
   gpc1_1 gpc1969 (
      {stage1_9[118]},
      {stage2_9[52]}
   );
   gpc1_1 gpc1970 (
      {stage1_9[119]},
      {stage2_9[53]}
   );
   gpc1_1 gpc1971 (
      {stage1_9[120]},
      {stage2_9[54]}
   );
   gpc1_1 gpc1972 (
      {stage1_9[121]},
      {stage2_9[55]}
   );
   gpc1_1 gpc1973 (
      {stage1_9[122]},
      {stage2_9[56]}
   );
   gpc1_1 gpc1974 (
      {stage1_9[123]},
      {stage2_9[57]}
   );
   gpc1_1 gpc1975 (
      {stage1_9[124]},
      {stage2_9[58]}
   );
   gpc1_1 gpc1976 (
      {stage1_9[125]},
      {stage2_9[59]}
   );
   gpc1_1 gpc1977 (
      {stage1_9[126]},
      {stage2_9[60]}
   );
   gpc1_1 gpc1978 (
      {stage1_9[127]},
      {stage2_9[61]}
   );
   gpc1_1 gpc1979 (
      {stage1_9[128]},
      {stage2_9[62]}
   );
   gpc1_1 gpc1980 (
      {stage1_9[129]},
      {stage2_9[63]}
   );
   gpc1_1 gpc1981 (
      {stage1_9[130]},
      {stage2_9[64]}
   );
   gpc1_1 gpc1982 (
      {stage1_9[131]},
      {stage2_9[65]}
   );
   gpc1_1 gpc1983 (
      {stage1_11[127]},
      {stage2_11[45]}
   );
   gpc1_1 gpc1984 (
      {stage1_11[128]},
      {stage2_11[46]}
   );
   gpc1_1 gpc1985 (
      {stage1_11[129]},
      {stage2_11[47]}
   );
   gpc1_1 gpc1986 (
      {stage1_11[130]},
      {stage2_11[48]}
   );
   gpc1_1 gpc1987 (
      {stage1_11[131]},
      {stage2_11[49]}
   );
   gpc1_1 gpc1988 (
      {stage1_11[132]},
      {stage2_11[50]}
   );
   gpc1_1 gpc1989 (
      {stage1_11[133]},
      {stage2_11[51]}
   );
   gpc1_1 gpc1990 (
      {stage1_11[134]},
      {stage2_11[52]}
   );
   gpc1_1 gpc1991 (
      {stage1_11[135]},
      {stage2_11[53]}
   );
   gpc1_1 gpc1992 (
      {stage1_11[136]},
      {stage2_11[54]}
   );
   gpc1_1 gpc1993 (
      {stage1_11[137]},
      {stage2_11[55]}
   );
   gpc1_1 gpc1994 (
      {stage1_11[138]},
      {stage2_11[56]}
   );
   gpc1_1 gpc1995 (
      {stage1_11[139]},
      {stage2_11[57]}
   );
   gpc1_1 gpc1996 (
      {stage1_12[173]},
      {stage2_12[50]}
   );
   gpc1_1 gpc1997 (
      {stage1_12[174]},
      {stage2_12[51]}
   );
   gpc1_1 gpc1998 (
      {stage1_12[175]},
      {stage2_12[52]}
   );
   gpc1_1 gpc1999 (
      {stage1_12[176]},
      {stage2_12[53]}
   );
   gpc1_1 gpc2000 (
      {stage1_12[177]},
      {stage2_12[54]}
   );
   gpc1_1 gpc2001 (
      {stage1_12[178]},
      {stage2_12[55]}
   );
   gpc1_1 gpc2002 (
      {stage1_12[179]},
      {stage2_12[56]}
   );
   gpc1_1 gpc2003 (
      {stage1_12[180]},
      {stage2_12[57]}
   );
   gpc1_1 gpc2004 (
      {stage1_12[181]},
      {stage2_12[58]}
   );
   gpc1_1 gpc2005 (
      {stage1_12[182]},
      {stage2_12[59]}
   );
   gpc1_1 gpc2006 (
      {stage1_12[183]},
      {stage2_12[60]}
   );
   gpc1_1 gpc2007 (
      {stage1_12[184]},
      {stage2_12[61]}
   );
   gpc1_1 gpc2008 (
      {stage1_12[185]},
      {stage2_12[62]}
   );
   gpc1_1 gpc2009 (
      {stage1_12[186]},
      {stage2_12[63]}
   );
   gpc1_1 gpc2010 (
      {stage1_12[187]},
      {stage2_12[64]}
   );
   gpc1_1 gpc2011 (
      {stage1_12[188]},
      {stage2_12[65]}
   );
   gpc1_1 gpc2012 (
      {stage1_12[189]},
      {stage2_12[66]}
   );
   gpc1_1 gpc2013 (
      {stage1_12[190]},
      {stage2_12[67]}
   );
   gpc1_1 gpc2014 (
      {stage1_12[191]},
      {stage2_12[68]}
   );
   gpc1_1 gpc2015 (
      {stage1_12[192]},
      {stage2_12[69]}
   );
   gpc1_1 gpc2016 (
      {stage1_12[193]},
      {stage2_12[70]}
   );
   gpc1_1 gpc2017 (
      {stage1_12[194]},
      {stage2_12[71]}
   );
   gpc1_1 gpc2018 (
      {stage1_12[195]},
      {stage2_12[72]}
   );
   gpc1_1 gpc2019 (
      {stage1_12[196]},
      {stage2_12[73]}
   );
   gpc1_1 gpc2020 (
      {stage1_12[197]},
      {stage2_12[74]}
   );
   gpc1_1 gpc2021 (
      {stage1_13[90]},
      {stage2_13[54]}
   );
   gpc1_1 gpc2022 (
      {stage1_13[91]},
      {stage2_13[55]}
   );
   gpc1_1 gpc2023 (
      {stage1_13[92]},
      {stage2_13[56]}
   );
   gpc1_1 gpc2024 (
      {stage1_14[66]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2025 (
      {stage1_14[67]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2026 (
      {stage1_14[68]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2027 (
      {stage1_14[69]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2028 (
      {stage1_14[70]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2029 (
      {stage1_14[71]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2030 (
      {stage1_14[72]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2031 (
      {stage1_14[73]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2032 (
      {stage1_14[74]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2033 (
      {stage1_14[75]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2034 (
      {stage1_14[76]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2035 (
      {stage1_14[77]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2036 (
      {stage1_14[78]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2037 (
      {stage1_14[79]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2038 (
      {stage1_14[80]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2039 (
      {stage1_14[81]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2040 (
      {stage1_14[82]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2041 (
      {stage1_14[83]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2042 (
      {stage1_14[84]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2043 (
      {stage1_14[85]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2044 (
      {stage1_14[86]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2045 (
      {stage1_14[87]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2046 (
      {stage1_14[88]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2047 (
      {stage1_14[89]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2048 (
      {stage1_14[90]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2049 (
      {stage1_14[91]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2050 (
      {stage1_14[92]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2051 (
      {stage1_14[93]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2052 (
      {stage1_14[94]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2053 (
      {stage1_14[95]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2054 (
      {stage1_14[96]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2055 (
      {stage1_14[97]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2056 (
      {stage1_14[98]},
      {stage2_14[74]}
   );
   gpc1_1 gpc2057 (
      {stage1_14[99]},
      {stage2_14[75]}
   );
   gpc1_1 gpc2058 (
      {stage1_14[100]},
      {stage2_14[76]}
   );
   gpc1_1 gpc2059 (
      {stage1_14[101]},
      {stage2_14[77]}
   );
   gpc1_1 gpc2060 (
      {stage1_14[102]},
      {stage2_14[78]}
   );
   gpc1_1 gpc2061 (
      {stage1_14[103]},
      {stage2_14[79]}
   );
   gpc1_1 gpc2062 (
      {stage1_14[104]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2063 (
      {stage1_14[105]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2064 (
      {stage1_14[106]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2065 (
      {stage1_14[107]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2066 (
      {stage1_14[108]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2067 (
      {stage1_14[109]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2068 (
      {stage1_14[110]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2069 (
      {stage1_14[111]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2070 (
      {stage1_14[112]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2071 (
      {stage1_14[113]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2072 (
      {stage1_15[84]},
      {stage2_15[38]}
   );
   gpc1_1 gpc2073 (
      {stage1_15[85]},
      {stage2_15[39]}
   );
   gpc1_1 gpc2074 (
      {stage1_15[86]},
      {stage2_15[40]}
   );
   gpc1_1 gpc2075 (
      {stage1_15[87]},
      {stage2_15[41]}
   );
   gpc1_1 gpc2076 (
      {stage1_15[88]},
      {stage2_15[42]}
   );
   gpc1_1 gpc2077 (
      {stage1_15[89]},
      {stage2_15[43]}
   );
   gpc1_1 gpc2078 (
      {stage1_15[90]},
      {stage2_15[44]}
   );
   gpc1_1 gpc2079 (
      {stage1_15[91]},
      {stage2_15[45]}
   );
   gpc1_1 gpc2080 (
      {stage1_15[92]},
      {stage2_15[46]}
   );
   gpc1_1 gpc2081 (
      {stage1_17[108]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2082 (
      {stage1_17[109]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2083 (
      {stage1_17[110]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2084 (
      {stage1_17[111]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2085 (
      {stage1_17[112]},
      {stage2_17[40]}
   );
   gpc1_1 gpc2086 (
      {stage1_17[113]},
      {stage2_17[41]}
   );
   gpc1_1 gpc2087 (
      {stage1_17[114]},
      {stage2_17[42]}
   );
   gpc1_1 gpc2088 (
      {stage1_17[115]},
      {stage2_17[43]}
   );
   gpc1_1 gpc2089 (
      {stage1_17[116]},
      {stage2_17[44]}
   );
   gpc1_1 gpc2090 (
      {stage1_17[117]},
      {stage2_17[45]}
   );
   gpc1_1 gpc2091 (
      {stage1_17[118]},
      {stage2_17[46]}
   );
   gpc1_1 gpc2092 (
      {stage1_17[119]},
      {stage2_17[47]}
   );
   gpc1_1 gpc2093 (
      {stage1_17[120]},
      {stage2_17[48]}
   );
   gpc1_1 gpc2094 (
      {stage1_17[121]},
      {stage2_17[49]}
   );
   gpc1_1 gpc2095 (
      {stage1_17[122]},
      {stage2_17[50]}
   );
   gpc1_1 gpc2096 (
      {stage1_17[123]},
      {stage2_17[51]}
   );
   gpc1_1 gpc2097 (
      {stage1_17[124]},
      {stage2_17[52]}
   );
   gpc1_1 gpc2098 (
      {stage1_17[125]},
      {stage2_17[53]}
   );
   gpc1_1 gpc2099 (
      {stage1_17[126]},
      {stage2_17[54]}
   );
   gpc1_1 gpc2100 (
      {stage1_18[94]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2101 (
      {stage1_18[95]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2102 (
      {stage1_18[96]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2103 (
      {stage1_18[97]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2104 (
      {stage1_18[98]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2105 (
      {stage1_18[99]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2106 (
      {stage1_18[100]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2107 (
      {stage1_18[101]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2108 (
      {stage1_18[102]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2109 (
      {stage1_18[103]},
      {stage2_18[43]}
   );
   gpc1_1 gpc2110 (
      {stage1_18[104]},
      {stage2_18[44]}
   );
   gpc1_1 gpc2111 (
      {stage1_18[105]},
      {stage2_18[45]}
   );
   gpc1_1 gpc2112 (
      {stage1_18[106]},
      {stage2_18[46]}
   );
   gpc1_1 gpc2113 (
      {stage1_18[107]},
      {stage2_18[47]}
   );
   gpc1_1 gpc2114 (
      {stage1_18[108]},
      {stage2_18[48]}
   );
   gpc1_1 gpc2115 (
      {stage1_18[109]},
      {stage2_18[49]}
   );
   gpc1_1 gpc2116 (
      {stage1_18[110]},
      {stage2_18[50]}
   );
   gpc1_1 gpc2117 (
      {stage1_18[111]},
      {stage2_18[51]}
   );
   gpc1_1 gpc2118 (
      {stage1_18[112]},
      {stage2_18[52]}
   );
   gpc1_1 gpc2119 (
      {stage1_18[113]},
      {stage2_18[53]}
   );
   gpc1_1 gpc2120 (
      {stage1_18[114]},
      {stage2_18[54]}
   );
   gpc1_1 gpc2121 (
      {stage1_18[115]},
      {stage2_18[55]}
   );
   gpc1_1 gpc2122 (
      {stage1_18[116]},
      {stage2_18[56]}
   );
   gpc1_1 gpc2123 (
      {stage1_18[117]},
      {stage2_18[57]}
   );
   gpc1_1 gpc2124 (
      {stage1_18[118]},
      {stage2_18[58]}
   );
   gpc1_1 gpc2125 (
      {stage1_18[119]},
      {stage2_18[59]}
   );
   gpc1_1 gpc2126 (
      {stage1_18[120]},
      {stage2_18[60]}
   );
   gpc1_1 gpc2127 (
      {stage1_18[121]},
      {stage2_18[61]}
   );
   gpc1_1 gpc2128 (
      {stage1_18[122]},
      {stage2_18[62]}
   );
   gpc1_1 gpc2129 (
      {stage1_18[123]},
      {stage2_18[63]}
   );
   gpc1_1 gpc2130 (
      {stage1_18[124]},
      {stage2_18[64]}
   );
   gpc1_1 gpc2131 (
      {stage1_18[125]},
      {stage2_18[65]}
   );
   gpc1_1 gpc2132 (
      {stage1_18[126]},
      {stage2_18[66]}
   );
   gpc1_1 gpc2133 (
      {stage1_18[127]},
      {stage2_18[67]}
   );
   gpc1_1 gpc2134 (
      {stage1_18[128]},
      {stage2_18[68]}
   );
   gpc1_1 gpc2135 (
      {stage1_18[129]},
      {stage2_18[69]}
   );
   gpc1_1 gpc2136 (
      {stage1_18[130]},
      {stage2_18[70]}
   );
   gpc1_1 gpc2137 (
      {stage1_18[131]},
      {stage2_18[71]}
   );
   gpc1_1 gpc2138 (
      {stage1_18[132]},
      {stage2_18[72]}
   );
   gpc1_1 gpc2139 (
      {stage1_18[133]},
      {stage2_18[73]}
   );
   gpc1_1 gpc2140 (
      {stage1_18[134]},
      {stage2_18[74]}
   );
   gpc1_1 gpc2141 (
      {stage1_18[135]},
      {stage2_18[75]}
   );
   gpc1_1 gpc2142 (
      {stage1_18[136]},
      {stage2_18[76]}
   );
   gpc1_1 gpc2143 (
      {stage1_18[137]},
      {stage2_18[77]}
   );
   gpc1_1 gpc2144 (
      {stage1_18[138]},
      {stage2_18[78]}
   );
   gpc1_1 gpc2145 (
      {stage1_18[139]},
      {stage2_18[79]}
   );
   gpc1_1 gpc2146 (
      {stage1_18[140]},
      {stage2_18[80]}
   );
   gpc1_1 gpc2147 (
      {stage1_18[141]},
      {stage2_18[81]}
   );
   gpc1_1 gpc2148 (
      {stage1_18[142]},
      {stage2_18[82]}
   );
   gpc1_1 gpc2149 (
      {stage1_18[143]},
      {stage2_18[83]}
   );
   gpc1_1 gpc2150 (
      {stage1_18[144]},
      {stage2_18[84]}
   );
   gpc1_1 gpc2151 (
      {stage1_18[145]},
      {stage2_18[85]}
   );
   gpc1_1 gpc2152 (
      {stage1_18[146]},
      {stage2_18[86]}
   );
   gpc1_1 gpc2153 (
      {stage1_18[147]},
      {stage2_18[87]}
   );
   gpc1_1 gpc2154 (
      {stage1_18[148]},
      {stage2_18[88]}
   );
   gpc1_1 gpc2155 (
      {stage1_18[149]},
      {stage2_18[89]}
   );
   gpc1_1 gpc2156 (
      {stage1_18[150]},
      {stage2_18[90]}
   );
   gpc1_1 gpc2157 (
      {stage1_19[93]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2158 (
      {stage1_20[23]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2159 (
      {stage1_20[24]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2160 (
      {stage1_20[25]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2161 (
      {stage1_20[26]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2162 (
      {stage1_20[27]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2163 (
      {stage1_20[28]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2164 (
      {stage1_20[29]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2165 (
      {stage1_20[30]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2166 (
      {stage1_20[31]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2167 (
      {stage1_20[32]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2168 (
      {stage1_20[33]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2169 (
      {stage1_20[34]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2170 (
      {stage1_20[35]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2171 (
      {stage1_20[36]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2172 (
      {stage1_20[37]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2173 (
      {stage1_20[38]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2174 (
      {stage1_20[39]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2175 (
      {stage1_20[40]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2176 (
      {stage1_20[41]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2177 (
      {stage1_20[42]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2178 (
      {stage1_20[43]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2179 (
      {stage1_20[44]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2180 (
      {stage1_20[45]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2181 (
      {stage1_20[46]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2182 (
      {stage1_20[47]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2183 (
      {stage1_20[48]},
      {stage2_20[58]}
   );
   gpc1_1 gpc2184 (
      {stage1_20[49]},
      {stage2_20[59]}
   );
   gpc1_1 gpc2185 (
      {stage1_20[50]},
      {stage2_20[60]}
   );
   gpc1_1 gpc2186 (
      {stage1_20[51]},
      {stage2_20[61]}
   );
   gpc1_1 gpc2187 (
      {stage1_20[52]},
      {stage2_20[62]}
   );
   gpc1_1 gpc2188 (
      {stage1_20[53]},
      {stage2_20[63]}
   );
   gpc1_1 gpc2189 (
      {stage1_20[54]},
      {stage2_20[64]}
   );
   gpc1_1 gpc2190 (
      {stage1_20[55]},
      {stage2_20[65]}
   );
   gpc1_1 gpc2191 (
      {stage1_20[56]},
      {stage2_20[66]}
   );
   gpc1_1 gpc2192 (
      {stage1_20[57]},
      {stage2_20[67]}
   );
   gpc1_1 gpc2193 (
      {stage1_20[58]},
      {stage2_20[68]}
   );
   gpc1_1 gpc2194 (
      {stage1_20[59]},
      {stage2_20[69]}
   );
   gpc1_1 gpc2195 (
      {stage1_20[60]},
      {stage2_20[70]}
   );
   gpc1_1 gpc2196 (
      {stage1_20[61]},
      {stage2_20[71]}
   );
   gpc1_1 gpc2197 (
      {stage1_20[62]},
      {stage2_20[72]}
   );
   gpc1_1 gpc2198 (
      {stage1_20[63]},
      {stage2_20[73]}
   );
   gpc1_1 gpc2199 (
      {stage1_20[64]},
      {stage2_20[74]}
   );
   gpc1_1 gpc2200 (
      {stage1_20[65]},
      {stage2_20[75]}
   );
   gpc1_1 gpc2201 (
      {stage1_20[66]},
      {stage2_20[76]}
   );
   gpc1_1 gpc2202 (
      {stage1_20[67]},
      {stage2_20[77]}
   );
   gpc1_1 gpc2203 (
      {stage1_20[68]},
      {stage2_20[78]}
   );
   gpc1_1 gpc2204 (
      {stage1_20[69]},
      {stage2_20[79]}
   );
   gpc1_1 gpc2205 (
      {stage1_20[70]},
      {stage2_20[80]}
   );
   gpc1_1 gpc2206 (
      {stage1_20[71]},
      {stage2_20[81]}
   );
   gpc1_1 gpc2207 (
      {stage1_20[72]},
      {stage2_20[82]}
   );
   gpc1_1 gpc2208 (
      {stage1_20[73]},
      {stage2_20[83]}
   );
   gpc1_1 gpc2209 (
      {stage1_20[74]},
      {stage2_20[84]}
   );
   gpc1_1 gpc2210 (
      {stage1_20[75]},
      {stage2_20[85]}
   );
   gpc1_1 gpc2211 (
      {stage1_20[76]},
      {stage2_20[86]}
   );
   gpc1_1 gpc2212 (
      {stage1_20[77]},
      {stage2_20[87]}
   );
   gpc1_1 gpc2213 (
      {stage1_20[78]},
      {stage2_20[88]}
   );
   gpc1_1 gpc2214 (
      {stage1_20[79]},
      {stage2_20[89]}
   );
   gpc1_1 gpc2215 (
      {stage1_20[80]},
      {stage2_20[90]}
   );
   gpc1_1 gpc2216 (
      {stage1_20[81]},
      {stage2_20[91]}
   );
   gpc1_1 gpc2217 (
      {stage1_20[82]},
      {stage2_20[92]}
   );
   gpc1_1 gpc2218 (
      {stage1_20[83]},
      {stage2_20[93]}
   );
   gpc1_1 gpc2219 (
      {stage1_20[84]},
      {stage2_20[94]}
   );
   gpc1_1 gpc2220 (
      {stage1_20[85]},
      {stage2_20[95]}
   );
   gpc1_1 gpc2221 (
      {stage1_20[86]},
      {stage2_20[96]}
   );
   gpc1_1 gpc2222 (
      {stage1_20[87]},
      {stage2_20[97]}
   );
   gpc1_1 gpc2223 (
      {stage1_20[88]},
      {stage2_20[98]}
   );
   gpc1_1 gpc2224 (
      {stage1_20[89]},
      {stage2_20[99]}
   );
   gpc1_1 gpc2225 (
      {stage1_20[90]},
      {stage2_20[100]}
   );
   gpc1_1 gpc2226 (
      {stage1_20[91]},
      {stage2_20[101]}
   );
   gpc1_1 gpc2227 (
      {stage1_20[92]},
      {stage2_20[102]}
   );
   gpc1_1 gpc2228 (
      {stage1_20[93]},
      {stage2_20[103]}
   );
   gpc1_1 gpc2229 (
      {stage1_20[94]},
      {stage2_20[104]}
   );
   gpc1_1 gpc2230 (
      {stage1_20[95]},
      {stage2_20[105]}
   );
   gpc1_1 gpc2231 (
      {stage1_20[96]},
      {stage2_20[106]}
   );
   gpc1_1 gpc2232 (
      {stage1_20[97]},
      {stage2_20[107]}
   );
   gpc1_1 gpc2233 (
      {stage1_20[98]},
      {stage2_20[108]}
   );
   gpc1_1 gpc2234 (
      {stage1_20[99]},
      {stage2_20[109]}
   );
   gpc1_1 gpc2235 (
      {stage1_20[100]},
      {stage2_20[110]}
   );
   gpc1_1 gpc2236 (
      {stage1_20[101]},
      {stage2_20[111]}
   );
   gpc1_1 gpc2237 (
      {stage1_20[102]},
      {stage2_20[112]}
   );
   gpc1_1 gpc2238 (
      {stage1_20[103]},
      {stage2_20[113]}
   );
   gpc1_1 gpc2239 (
      {stage1_20[104]},
      {stage2_20[114]}
   );
   gpc1_1 gpc2240 (
      {stage1_20[105]},
      {stage2_20[115]}
   );
   gpc1_1 gpc2241 (
      {stage1_20[106]},
      {stage2_20[116]}
   );
   gpc1_1 gpc2242 (
      {stage1_20[107]},
      {stage2_20[117]}
   );
   gpc1_1 gpc2243 (
      {stage1_20[108]},
      {stage2_20[118]}
   );
   gpc1_1 gpc2244 (
      {stage1_20[109]},
      {stage2_20[119]}
   );
   gpc1_1 gpc2245 (
      {stage1_20[110]},
      {stage2_20[120]}
   );
   gpc1_1 gpc2246 (
      {stage1_20[111]},
      {stage2_20[121]}
   );
   gpc1_1 gpc2247 (
      {stage1_20[112]},
      {stage2_20[122]}
   );
   gpc1_1 gpc2248 (
      {stage1_20[113]},
      {stage2_20[123]}
   );
   gpc1_1 gpc2249 (
      {stage1_20[114]},
      {stage2_20[124]}
   );
   gpc1_1 gpc2250 (
      {stage1_20[115]},
      {stage2_20[125]}
   );
   gpc1_1 gpc2251 (
      {stage1_21[90]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2252 (
      {stage1_21[91]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2253 (
      {stage1_21[92]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2254 (
      {stage1_21[93]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2255 (
      {stage1_21[94]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2256 (
      {stage1_21[95]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2257 (
      {stage1_21[96]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2258 (
      {stage1_21[97]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2259 (
      {stage1_21[98]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2260 (
      {stage1_21[99]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2261 (
      {stage1_21[100]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2262 (
      {stage1_21[101]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2263 (
      {stage1_21[102]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2264 (
      {stage1_21[103]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2265 (
      {stage1_21[104]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2266 (
      {stage1_21[105]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2267 (
      {stage1_21[106]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2268 (
      {stage1_21[107]},
      {stage2_21[40]}
   );
   gpc1_1 gpc2269 (
      {stage1_21[108]},
      {stage2_21[41]}
   );
   gpc1_1 gpc2270 (
      {stage1_21[109]},
      {stage2_21[42]}
   );
   gpc1_1 gpc2271 (
      {stage1_21[110]},
      {stage2_21[43]}
   );
   gpc1_1 gpc2272 (
      {stage1_21[111]},
      {stage2_21[44]}
   );
   gpc1_1 gpc2273 (
      {stage1_21[112]},
      {stage2_21[45]}
   );
   gpc1_1 gpc2274 (
      {stage1_21[113]},
      {stage2_21[46]}
   );
   gpc1_1 gpc2275 (
      {stage1_21[114]},
      {stage2_21[47]}
   );
   gpc1_1 gpc2276 (
      {stage1_21[115]},
      {stage2_21[48]}
   );
   gpc1_1 gpc2277 (
      {stage1_21[116]},
      {stage2_21[49]}
   );
   gpc1_1 gpc2278 (
      {stage1_21[117]},
      {stage2_21[50]}
   );
   gpc1_1 gpc2279 (
      {stage1_21[118]},
      {stage2_21[51]}
   );
   gpc1_1 gpc2280 (
      {stage1_21[119]},
      {stage2_21[52]}
   );
   gpc1_1 gpc2281 (
      {stage1_21[120]},
      {stage2_21[53]}
   );
   gpc1_1 gpc2282 (
      {stage1_21[121]},
      {stage2_21[54]}
   );
   gpc1_1 gpc2283 (
      {stage1_21[122]},
      {stage2_21[55]}
   );
   gpc1_1 gpc2284 (
      {stage1_21[123]},
      {stage2_21[56]}
   );
   gpc1_1 gpc2285 (
      {stage1_21[124]},
      {stage2_21[57]}
   );
   gpc1_1 gpc2286 (
      {stage1_21[125]},
      {stage2_21[58]}
   );
   gpc1_1 gpc2287 (
      {stage1_21[126]},
      {stage2_21[59]}
   );
   gpc1_1 gpc2288 (
      {stage1_21[127]},
      {stage2_21[60]}
   );
   gpc1_1 gpc2289 (
      {stage1_21[128]},
      {stage2_21[61]}
   );
   gpc1_1 gpc2290 (
      {stage1_21[129]},
      {stage2_21[62]}
   );
   gpc1_1 gpc2291 (
      {stage1_21[130]},
      {stage2_21[63]}
   );
   gpc1_1 gpc2292 (
      {stage1_21[131]},
      {stage2_21[64]}
   );
   gpc1_1 gpc2293 (
      {stage1_21[132]},
      {stage2_21[65]}
   );
   gpc1_1 gpc2294 (
      {stage1_21[133]},
      {stage2_21[66]}
   );
   gpc1_1 gpc2295 (
      {stage1_21[134]},
      {stage2_21[67]}
   );
   gpc1_1 gpc2296 (
      {stage1_21[135]},
      {stage2_21[68]}
   );
   gpc1_1 gpc2297 (
      {stage1_21[136]},
      {stage2_21[69]}
   );
   gpc1_1 gpc2298 (
      {stage1_21[137]},
      {stage2_21[70]}
   );
   gpc1_1 gpc2299 (
      {stage1_21[138]},
      {stage2_21[71]}
   );
   gpc1_1 gpc2300 (
      {stage1_22[77]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2301 (
      {stage1_22[78]},
      {stage2_22[31]}
   );
   gpc1_1 gpc2302 (
      {stage1_22[79]},
      {stage2_22[32]}
   );
   gpc1_1 gpc2303 (
      {stage1_22[80]},
      {stage2_22[33]}
   );
   gpc1_1 gpc2304 (
      {stage1_22[81]},
      {stage2_22[34]}
   );
   gpc1_1 gpc2305 (
      {stage1_22[82]},
      {stage2_22[35]}
   );
   gpc1_1 gpc2306 (
      {stage1_22[83]},
      {stage2_22[36]}
   );
   gpc1_1 gpc2307 (
      {stage1_22[84]},
      {stage2_22[37]}
   );
   gpc1_1 gpc2308 (
      {stage1_22[85]},
      {stage2_22[38]}
   );
   gpc1_1 gpc2309 (
      {stage1_22[86]},
      {stage2_22[39]}
   );
   gpc1_1 gpc2310 (
      {stage1_22[87]},
      {stage2_22[40]}
   );
   gpc1_1 gpc2311 (
      {stage1_22[88]},
      {stage2_22[41]}
   );
   gpc1_1 gpc2312 (
      {stage1_22[89]},
      {stage2_22[42]}
   );
   gpc1_1 gpc2313 (
      {stage1_22[90]},
      {stage2_22[43]}
   );
   gpc1_1 gpc2314 (
      {stage1_22[91]},
      {stage2_22[44]}
   );
   gpc1_1 gpc2315 (
      {stage1_22[92]},
      {stage2_22[45]}
   );
   gpc1_1 gpc2316 (
      {stage1_22[93]},
      {stage2_22[46]}
   );
   gpc1_1 gpc2317 (
      {stage1_23[73]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2318 (
      {stage1_23[74]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2319 (
      {stage1_23[75]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2320 (
      {stage1_23[76]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2321 (
      {stage1_23[77]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2322 (
      {stage1_23[78]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2323 (
      {stage1_23[79]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2324 (
      {stage1_23[80]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2325 (
      {stage1_23[81]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2326 (
      {stage1_23[82]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2327 (
      {stage1_23[83]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2328 (
      {stage1_23[84]},
      {stage2_23[47]}
   );
   gpc1_1 gpc2329 (
      {stage1_23[85]},
      {stage2_23[48]}
   );
   gpc1_1 gpc2330 (
      {stage1_23[86]},
      {stage2_23[49]}
   );
   gpc1_1 gpc2331 (
      {stage1_23[87]},
      {stage2_23[50]}
   );
   gpc1_1 gpc2332 (
      {stage1_23[88]},
      {stage2_23[51]}
   );
   gpc1_1 gpc2333 (
      {stage1_23[89]},
      {stage2_23[52]}
   );
   gpc1_1 gpc2334 (
      {stage1_23[90]},
      {stage2_23[53]}
   );
   gpc1_1 gpc2335 (
      {stage1_23[91]},
      {stage2_23[54]}
   );
   gpc1_1 gpc2336 (
      {stage1_23[92]},
      {stage2_23[55]}
   );
   gpc1_1 gpc2337 (
      {stage1_23[93]},
      {stage2_23[56]}
   );
   gpc1_1 gpc2338 (
      {stage1_24[249]},
      {stage2_24[59]}
   );
   gpc1_1 gpc2339 (
      {stage1_24[250]},
      {stage2_24[60]}
   );
   gpc1_1 gpc2340 (
      {stage1_24[251]},
      {stage2_24[61]}
   );
   gpc1_1 gpc2341 (
      {stage1_24[252]},
      {stage2_24[62]}
   );
   gpc1_1 gpc2342 (
      {stage1_24[253]},
      {stage2_24[63]}
   );
   gpc1_1 gpc2343 (
      {stage1_25[117]},
      {stage2_25[65]}
   );
   gpc1_1 gpc2344 (
      {stage1_27[73]},
      {stage2_27[61]}
   );
   gpc1_1 gpc2345 (
      {stage1_27[74]},
      {stage2_27[62]}
   );
   gpc1_1 gpc2346 (
      {stage1_27[75]},
      {stage2_27[63]}
   );
   gpc1_1 gpc2347 (
      {stage1_27[76]},
      {stage2_27[64]}
   );
   gpc1_1 gpc2348 (
      {stage1_27[77]},
      {stage2_27[65]}
   );
   gpc1_1 gpc2349 (
      {stage1_27[78]},
      {stage2_27[66]}
   );
   gpc1_1 gpc2350 (
      {stage1_27[79]},
      {stage2_27[67]}
   );
   gpc1_1 gpc2351 (
      {stage1_27[80]},
      {stage2_27[68]}
   );
   gpc1_1 gpc2352 (
      {stage1_27[81]},
      {stage2_27[69]}
   );
   gpc1_1 gpc2353 (
      {stage1_27[82]},
      {stage2_27[70]}
   );
   gpc1_1 gpc2354 (
      {stage1_27[83]},
      {stage2_27[71]}
   );
   gpc1_1 gpc2355 (
      {stage1_27[84]},
      {stage2_27[72]}
   );
   gpc1_1 gpc2356 (
      {stage1_27[85]},
      {stage2_27[73]}
   );
   gpc1_1 gpc2357 (
      {stage1_27[86]},
      {stage2_27[74]}
   );
   gpc1_1 gpc2358 (
      {stage1_27[87]},
      {stage2_27[75]}
   );
   gpc1_1 gpc2359 (
      {stage1_27[88]},
      {stage2_27[76]}
   );
   gpc1_1 gpc2360 (
      {stage1_27[89]},
      {stage2_27[77]}
   );
   gpc1_1 gpc2361 (
      {stage1_27[90]},
      {stage2_27[78]}
   );
   gpc1_1 gpc2362 (
      {stage1_27[91]},
      {stage2_27[79]}
   );
   gpc1_1 gpc2363 (
      {stage1_27[92]},
      {stage2_27[80]}
   );
   gpc1_1 gpc2364 (
      {stage1_27[93]},
      {stage2_27[81]}
   );
   gpc1_1 gpc2365 (
      {stage1_27[94]},
      {stage2_27[82]}
   );
   gpc1_1 gpc2366 (
      {stage1_27[95]},
      {stage2_27[83]}
   );
   gpc1_1 gpc2367 (
      {stage1_27[96]},
      {stage2_27[84]}
   );
   gpc1_1 gpc2368 (
      {stage1_27[97]},
      {stage2_27[85]}
   );
   gpc1_1 gpc2369 (
      {stage1_27[98]},
      {stage2_27[86]}
   );
   gpc1_1 gpc2370 (
      {stage1_27[99]},
      {stage2_27[87]}
   );
   gpc1_1 gpc2371 (
      {stage1_27[100]},
      {stage2_27[88]}
   );
   gpc1_1 gpc2372 (
      {stage1_27[101]},
      {stage2_27[89]}
   );
   gpc1_1 gpc2373 (
      {stage1_27[102]},
      {stage2_27[90]}
   );
   gpc1_1 gpc2374 (
      {stage1_27[103]},
      {stage2_27[91]}
   );
   gpc1_1 gpc2375 (
      {stage1_27[104]},
      {stage2_27[92]}
   );
   gpc1_1 gpc2376 (
      {stage1_27[105]},
      {stage2_27[93]}
   );
   gpc1_1 gpc2377 (
      {stage1_27[106]},
      {stage2_27[94]}
   );
   gpc1_1 gpc2378 (
      {stage1_27[107]},
      {stage2_27[95]}
   );
   gpc1_1 gpc2379 (
      {stage1_28[90]},
      {stage2_28[60]}
   );
   gpc1_1 gpc2380 (
      {stage1_28[91]},
      {stage2_28[61]}
   );
   gpc1_1 gpc2381 (
      {stage1_28[92]},
      {stage2_28[62]}
   );
   gpc1_1 gpc2382 (
      {stage1_28[93]},
      {stage2_28[63]}
   );
   gpc1_1 gpc2383 (
      {stage1_28[94]},
      {stage2_28[64]}
   );
   gpc1_1 gpc2384 (
      {stage1_28[95]},
      {stage2_28[65]}
   );
   gpc1_1 gpc2385 (
      {stage1_28[96]},
      {stage2_28[66]}
   );
   gpc1_1 gpc2386 (
      {stage1_28[97]},
      {stage2_28[67]}
   );
   gpc1_1 gpc2387 (
      {stage1_28[98]},
      {stage2_28[68]}
   );
   gpc1_1 gpc2388 (
      {stage1_28[99]},
      {stage2_28[69]}
   );
   gpc1_1 gpc2389 (
      {stage1_28[100]},
      {stage2_28[70]}
   );
   gpc1_1 gpc2390 (
      {stage1_28[101]},
      {stage2_28[71]}
   );
   gpc1_1 gpc2391 (
      {stage1_31[129]},
      {stage2_31[44]}
   );
   gpc1_1 gpc2392 (
      {stage1_31[130]},
      {stage2_31[45]}
   );
   gpc1_1 gpc2393 (
      {stage1_31[131]},
      {stage2_31[46]}
   );
   gpc1_1 gpc2394 (
      {stage1_31[132]},
      {stage2_31[47]}
   );
   gpc1_1 gpc2395 (
      {stage1_32[68]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2396 (
      {stage1_32[69]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2397 (
      {stage1_32[70]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2398 (
      {stage1_32[71]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2399 (
      {stage1_32[72]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2400 (
      {stage1_32[73]},
      {stage2_32[43]}
   );
   gpc117_4 gpc2401 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_1[0]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc117_4 gpc2402 (
      {stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[1]},
      {stage2_2[1]},
      {stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc2403 (
      {stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc2404 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21]},
      {stage2_1[8]},
      {stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage3_4[1],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc2405 (
      {stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc2406 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3],stage3_3[5]}
   );
   gpc615_5 gpc2407 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[2],stage3_4[4],stage3_3[6]}
   );
   gpc615_5 gpc2408 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[3],stage3_4[5],stage3_3[7]}
   );
   gpc606_5 gpc2409 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[4],stage3_4[6]}
   );
   gpc606_5 gpc2410 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc2411 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[6],stage3_4[8]}
   );
   gpc615_5 gpc2412 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[7],stage3_5[7],stage3_4[9]}
   );
   gpc615_5 gpc2413 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[8],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc2414 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[9],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc2415 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[10],stage3_5[10],stage3_4[12]}
   );
   gpc615_5 gpc2416 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[11],stage3_5[11],stage3_4[13]}
   );
   gpc606_5 gpc2417 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[12],stage3_5[12]}
   );
   gpc606_5 gpc2418 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[13],stage3_5[13]}
   );
   gpc606_5 gpc2419 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[14],stage3_5[14]}
   );
   gpc615_5 gpc2420 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[11],stage3_7[14]}
   );
   gpc615_5 gpc2421 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[12],stage3_7[15]}
   );
   gpc615_5 gpc2422 (
      {stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[2]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc2423 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37]},
      {stage2_8[3]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[3],stage3_9[6],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc2424 (
      {stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42]},
      {stage2_8[4]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[4],stage3_9[7],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc2425 (
      {stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage2_8[5]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[5],stage3_9[8],stage3_8[16],stage3_7[19]}
   );
   gpc623_5 gpc2426 (
      {stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[6], stage2_8[7]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[6],stage3_9[9],stage3_8[17],stage3_7[20]}
   );
   gpc606_5 gpc2427 (
      {stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[7],stage3_10[7],stage3_9[10],stage3_8[18]}
   );
   gpc606_5 gpc2428 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[8],stage3_10[8],stage3_9[11],stage3_8[19]}
   );
   gpc606_5 gpc2429 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[9],stage3_10[9],stage3_9[12],stage3_8[20]}
   );
   gpc606_5 gpc2430 (
      {stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[10],stage3_10[10],stage3_9[13],stage3_8[21]}
   );
   gpc606_5 gpc2431 (
      {stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[11],stage3_10[11],stage3_9[14],stage3_8[22]}
   );
   gpc606_5 gpc2432 (
      {stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[12],stage3_10[12],stage3_9[15],stage3_8[23]}
   );
   gpc606_5 gpc2433 (
      {stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[13],stage3_10[13],stage3_9[16],stage3_8[24]}
   );
   gpc615_5 gpc2434 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[42]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[14],stage3_10[14],stage3_9[17],stage3_8[25]}
   );
   gpc606_5 gpc2435 (
      {stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[8],stage3_11[15],stage3_10[15],stage3_9[18]}
   );
   gpc606_5 gpc2436 (
      {stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[9],stage3_11[16],stage3_10[16],stage3_9[19]}
   );
   gpc606_5 gpc2437 (
      {stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[10],stage3_11[17],stage3_10[17],stage3_9[20]}
   );
   gpc615_5 gpc2438 (
      {stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[48]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[11],stage3_11[18],stage3_10[18],stage3_9[21]}
   );
   gpc615_5 gpc2439 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[12],stage3_11[19]}
   );
   gpc615_5 gpc2440 (
      {stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_12[1]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[13],stage3_11[20]}
   );
   gpc615_5 gpc2441 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_12[2]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[14],stage3_11[21]}
   );
   gpc615_5 gpc2442 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_12[3]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[15],stage3_11[22]}
   );
   gpc615_5 gpc2443 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48]},
      {stage2_12[4]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[16],stage3_11[23]}
   );
   gpc615_5 gpc2444 (
      {stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage2_12[5]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[17],stage3_11[24]}
   );
   gpc615_5 gpc2445 (
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], 1'b0},
      {stage2_12[6]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[6],stage3_13[10],stage3_12[18],stage3_11[25]}
   );
   gpc606_5 gpc2446 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[7],stage3_13[11],stage3_12[19]}
   );
   gpc606_5 gpc2447 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[8],stage3_13[12],stage3_12[20]}
   );
   gpc606_5 gpc2448 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[9],stage3_13[13],stage3_12[21]}
   );
   gpc606_5 gpc2449 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[10],stage3_13[14],stage3_12[22]}
   );
   gpc606_5 gpc2450 (
      {stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[11],stage3_14[11],stage3_13[15],stage3_12[23]}
   );
   gpc606_5 gpc2451 (
      {stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[12],stage3_14[12],stage3_13[16],stage3_12[24]}
   );
   gpc606_5 gpc2452 (
      {stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[13],stage3_14[13],stage3_13[17],stage3_12[25]}
   );
   gpc606_5 gpc2453 (
      {stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[14],stage3_14[14],stage3_13[18],stage3_12[26]}
   );
   gpc606_5 gpc2454 (
      {stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[15],stage3_14[15],stage3_13[19],stage3_12[27]}
   );
   gpc606_5 gpc2455 (
      {stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[16],stage3_14[16],stage3_13[20],stage3_12[28]}
   );
   gpc606_5 gpc2456 (
      {stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[17],stage3_14[17],stage3_13[21],stage3_12[29]}
   );
   gpc615_5 gpc2457 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[11],stage3_15[18],stage3_14[18]}
   );
   gpc615_5 gpc2458 (
      {stage2_14[71], stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[12],stage3_15[19],stage3_14[19]}
   );
   gpc615_5 gpc2459 (
      {stage2_14[76], stage2_14[77], stage2_14[78], stage2_14[79], stage2_14[80]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[13],stage3_15[20],stage3_14[20]}
   );
   gpc615_5 gpc2460 (
      {stage2_14[81], stage2_14[82], stage2_14[83], stage2_14[84], stage2_14[85]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[14],stage3_15[21],stage3_14[21]}
   );
   gpc615_5 gpc2461 (
      {stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8]},
      {stage2_16[24]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[4],stage3_17[4],stage3_16[15],stage3_15[22]}
   );
   gpc615_5 gpc2462 (
      {stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13]},
      {stage2_16[25]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[5],stage3_17[5],stage3_16[16],stage3_15[23]}
   );
   gpc615_5 gpc2463 (
      {stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18]},
      {stage2_16[26]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[6],stage3_17[6],stage3_16[17],stage3_15[24]}
   );
   gpc615_5 gpc2464 (
      {stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage2_16[27]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[7],stage3_17[7],stage3_16[18],stage3_15[25]}
   );
   gpc615_5 gpc2465 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[28]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[8],stage3_17[8],stage3_16[19],stage3_15[26]}
   );
   gpc615_5 gpc2466 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[29]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[9],stage3_17[9],stage3_16[20],stage3_15[27]}
   );
   gpc615_5 gpc2467 (
      {stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38]},
      {stage2_16[30]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[10],stage3_17[10],stage3_16[21],stage3_15[28]}
   );
   gpc615_5 gpc2468 (
      {stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43]},
      {stage2_16[31]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[11],stage3_17[11],stage3_16[22],stage3_15[29]}
   );
   gpc606_5 gpc2469 (
      {stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35], stage2_16[36], stage2_16[37]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[12],stage3_17[12],stage3_16[23]}
   );
   gpc615_5 gpc2470 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[0]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[9],stage3_18[13]}
   );
   gpc615_5 gpc2471 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[1]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[10],stage3_18[14]}
   );
   gpc615_5 gpc2472 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[2]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[11],stage3_18[15]}
   );
   gpc615_5 gpc2473 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[3]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[12],stage3_18[16]}
   );
   gpc615_5 gpc2474 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[4]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[13],stage3_18[17]}
   );
   gpc615_5 gpc2475 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage2_19[5]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[14],stage3_18[18]}
   );
   gpc615_5 gpc2476 (
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40]},
      {stage2_19[6]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[15],stage3_18[19]}
   );
   gpc615_5 gpc2477 (
      {stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45]},
      {stage2_19[7]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[16],stage3_18[20]}
   );
   gpc615_5 gpc2478 (
      {stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50]},
      {stage2_19[8]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[17],stage3_18[21]}
   );
   gpc615_5 gpc2479 (
      {stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55]},
      {stage2_19[9]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[18],stage3_18[22]}
   );
   gpc615_5 gpc2480 (
      {stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_19[10]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[19],stage3_18[23]}
   );
   gpc615_5 gpc2481 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65]},
      {stage2_19[11]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[20],stage3_18[24]}
   );
   gpc615_5 gpc2482 (
      {stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70]},
      {stage2_19[12]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[21],stage3_18[25]}
   );
   gpc615_5 gpc2483 (
      {stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75]},
      {stage2_19[13]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[22],stage3_18[26]}
   );
   gpc615_5 gpc2484 (
      {stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80]},
      {stage2_19[14]},
      {stage2_20[84], stage2_20[85], stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89]},
      {stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[23],stage3_18[27]}
   );
   gpc615_5 gpc2485 (
      {stage2_19[15], stage2_19[16], stage2_19[17], stage2_19[18], stage2_19[19]},
      {stage2_20[90]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[24]}
   );
   gpc615_5 gpc2486 (
      {stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23], stage2_19[24]},
      {stage2_20[91]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[25]}
   );
   gpc615_5 gpc2487 (
      {stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[92]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[26]}
   );
   gpc615_5 gpc2488 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34]},
      {stage2_20[93]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[27]}
   );
   gpc615_5 gpc2489 (
      {stage2_19[35], stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39]},
      {stage2_20[94]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[28]}
   );
   gpc606_5 gpc2490 (
      {stage2_20[95], stage2_20[96], stage2_20[97], stage2_20[98], stage2_20[99], stage2_20[100]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[20],stage3_21[20],stage3_20[21]}
   );
   gpc606_5 gpc2491 (
      {stage2_20[101], stage2_20[102], stage2_20[103], stage2_20[104], stage2_20[105], stage2_20[106]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[21],stage3_21[21],stage3_20[22]}
   );
   gpc606_5 gpc2492 (
      {stage2_20[107], stage2_20[108], stage2_20[109], stage2_20[110], stage2_20[111], stage2_20[112]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc1343_5 gpc2493 (
      {stage2_21[30], stage2_21[31], stage2_21[32]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[0], stage2_23[1], stage2_23[2]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[3],stage3_23[8],stage3_22[23],stage3_21[23]}
   );
   gpc1343_5 gpc2494 (
      {stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage2_22[22], stage2_22[23], stage2_22[24], stage2_22[25]},
      {stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[4],stage3_23[9],stage3_22[24],stage3_21[24]}
   );
   gpc1343_5 gpc2495 (
      {stage2_21[36], stage2_21[37], stage2_21[38]},
      {stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_23[6], stage2_23[7], stage2_23[8]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[5],stage3_23[10],stage3_22[25],stage3_21[25]}
   );
   gpc615_5 gpc2496 (
      {stage2_21[39], stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43]},
      {stage2_22[30]},
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage3_25[3],stage3_24[6],stage3_23[11],stage3_22[26],stage3_21[26]}
   );
   gpc615_5 gpc2497 (
      {stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47], stage2_21[48]},
      {stage2_22[31]},
      {stage2_23[15], stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage3_25[4],stage3_24[7],stage3_23[12],stage3_22[27],stage3_21[27]}
   );
   gpc615_5 gpc2498 (
      {stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage2_22[32]},
      {stage2_23[21], stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage3_25[5],stage3_24[8],stage3_23[13],stage3_22[28],stage3_21[28]}
   );
   gpc615_5 gpc2499 (
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58]},
      {stage2_22[33]},
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32]},
      {stage3_25[6],stage3_24[9],stage3_23[14],stage3_22[29],stage3_21[29]}
   );
   gpc615_5 gpc2500 (
      {stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_22[34]},
      {stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage3_25[7],stage3_24[10],stage3_23[15],stage3_22[30],stage3_21[30]}
   );
   gpc615_5 gpc2501 (
      {stage2_21[64], stage2_21[65], stage2_21[66], stage2_21[67], stage2_21[68]},
      {stage2_22[35]},
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage3_25[8],stage3_24[11],stage3_23[16],stage3_22[31],stage3_21[31]}
   );
   gpc615_5 gpc2502 (
      {stage2_21[69], stage2_21[70], stage2_21[71], 1'b0, 1'b0},
      {stage2_22[36]},
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage3_25[9],stage3_24[12],stage3_23[17],stage3_22[32],stage3_21[32]}
   );
   gpc615_5 gpc2503 (
      {stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[51]},
      {stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7], stage2_24[8]},
      {stage3_26[0],stage3_25[10],stage3_24[13],stage3_23[18],stage3_22[33]}
   );
   gpc615_5 gpc2504 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[52]},
      {stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13], stage2_24[14]},
      {stage3_26[1],stage3_25[11],stage3_24[14],stage3_23[19],stage3_22[34]}
   );
   gpc615_5 gpc2505 (
      {stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56], 1'b0},
      {stage2_24[15]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[2],stage3_25[12],stage3_24[15],stage3_23[20]}
   );
   gpc606_5 gpc2506 (
      {stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[3],stage3_25[13],stage3_24[16]}
   );
   gpc606_5 gpc2507 (
      {stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[2],stage3_26[4],stage3_25[14],stage3_24[17]}
   );
   gpc606_5 gpc2508 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[3],stage3_26[5],stage3_25[15],stage3_24[18]}
   );
   gpc606_5 gpc2509 (
      {stage2_24[34], stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[4],stage3_26[6],stage3_25[16],stage3_24[19]}
   );
   gpc606_5 gpc2510 (
      {stage2_24[40], stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[5],stage3_26[7],stage3_25[17],stage3_24[20]}
   );
   gpc606_5 gpc2511 (
      {stage2_24[46], stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[6],stage3_26[8],stage3_25[18],stage3_24[21]}
   );
   gpc606_5 gpc2512 (
      {stage2_24[52], stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[7],stage3_26[9],stage3_25[19],stage3_24[22]}
   );
   gpc606_5 gpc2513 (
      {stage2_24[58], stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[8],stage3_26[10],stage3_25[20],stage3_24[23]}
   );
   gpc606_5 gpc2514 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[8],stage3_27[9],stage3_26[11],stage3_25[21]}
   );
   gpc606_5 gpc2515 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[9],stage3_27[10],stage3_26[12],stage3_25[22]}
   );
   gpc606_5 gpc2516 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[10],stage3_27[11],stage3_26[13],stage3_25[23]}
   );
   gpc606_5 gpc2517 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[11],stage3_27[12],stage3_26[14],stage3_25[24]}
   );
   gpc606_5 gpc2518 (
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[12],stage3_27[13],stage3_26[15],stage3_25[25]}
   );
   gpc606_5 gpc2519 (
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage3_29[5],stage3_28[13],stage3_27[14],stage3_26[16],stage3_25[26]}
   );
   gpc606_5 gpc2520 (
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage3_29[6],stage3_28[14],stage3_27[15],stage3_26[17],stage3_25[27]}
   );
   gpc606_5 gpc2521 (
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage3_29[7],stage3_28[15],stage3_27[16],stage3_26[18],stage3_25[28]}
   );
   gpc606_5 gpc2522 (
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage3_29[8],stage3_28[16],stage3_27[17],stage3_26[19],stage3_25[29]}
   );
   gpc615_5 gpc2523 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[9],stage3_28[17],stage3_27[18],stage3_26[20]}
   );
   gpc615_5 gpc2524 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[55]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[10],stage3_28[18],stage3_27[19],stage3_26[21]}
   );
   gpc615_5 gpc2525 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[56]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[11],stage3_28[19],stage3_27[20],stage3_26[22]}
   );
   gpc615_5 gpc2526 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[57]},
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage3_30[3],stage3_29[12],stage3_28[20],stage3_27[21],stage3_26[23]}
   );
   gpc606_5 gpc2527 (
      {stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[4],stage3_29[13],stage3_28[21],stage3_27[22]}
   );
   gpc615_5 gpc2528 (
      {stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[24]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[5],stage3_29[14],stage3_28[22],stage3_27[23]}
   );
   gpc615_5 gpc2529 (
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73]},
      {stage2_28[25]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[6],stage3_29[15],stage3_28[23],stage3_27[24]}
   );
   gpc615_5 gpc2530 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78]},
      {stage2_28[26]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[7],stage3_29[16],stage3_28[24],stage3_27[25]}
   );
   gpc615_5 gpc2531 (
      {stage2_27[79], stage2_27[80], stage2_27[81], stage2_27[82], stage2_27[83]},
      {stage2_28[27]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[8],stage3_29[17],stage3_28[25],stage3_27[26]}
   );
   gpc606_5 gpc2532 (
      {stage2_28[28], stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[5],stage3_30[9],stage3_29[18],stage3_28[26]}
   );
   gpc606_5 gpc2533 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[6],stage3_30[10],stage3_29[19],stage3_28[27]}
   );
   gpc606_5 gpc2534 (
      {stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[7],stage3_30[11],stage3_29[20],stage3_28[28]}
   );
   gpc606_5 gpc2535 (
      {stage2_28[46], stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[8],stage3_30[12],stage3_29[21],stage3_28[29]}
   );
   gpc606_5 gpc2536 (
      {stage2_28[52], stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[9],stage3_30[13],stage3_29[22],stage3_28[30]}
   );
   gpc606_5 gpc2537 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[5],stage3_31[10],stage3_30[14],stage3_29[23]}
   );
   gpc615_5 gpc2538 (
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[6],stage3_31[11],stage3_30[15]}
   );
   gpc615_5 gpc2539 (
      {stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39]},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[7],stage3_31[12],stage3_30[16]}
   );
   gpc615_5 gpc2540 (
      {stage2_30[40], stage2_30[41], stage2_30[42], stage2_30[43], stage2_30[44]},
      {stage2_31[8]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[3],stage3_32[8],stage3_31[13],stage3_30[17]}
   );
   gpc615_5 gpc2541 (
      {stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12], stage2_31[13]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[4],stage3_32[9],stage3_31[14]}
   );
   gpc615_5 gpc2542 (
      {stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17], stage2_31[18]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[5],stage3_32[10],stage3_31[15]}
   );
   gpc615_5 gpc2543 (
      {stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[6],stage3_32[11],stage3_31[16]}
   );
   gpc615_5 gpc2544 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[7],stage3_32[12],stage3_31[17]}
   );
   gpc606_5 gpc2545 (
      {stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[7],stage3_33[8],stage3_32[13]}
   );
   gpc606_5 gpc2546 (
      {stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[8],stage3_33[9],stage3_32[14]}
   );
   gpc606_5 gpc2547 (
      {stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], 1'b0},
      {stage3_36[2],stage3_35[6],stage3_34[9],stage3_33[10],stage3_32[15]}
   );
   gpc1_1 gpc2548 (
      {stage2_0[22]},
      {stage3_0[4]}
   );
   gpc1_1 gpc2549 (
      {stage2_0[23]},
      {stage3_0[5]}
   );
   gpc1_1 gpc2550 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc2551 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc2552 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc2553 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc2554 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc2555 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc2556 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc2557 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc2558 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc2559 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc2560 (
      {stage2_1[19]},
      {stage3_1[14]}
   );
   gpc1_1 gpc2561 (
      {stage2_1[20]},
      {stage3_1[15]}
   );
   gpc1_1 gpc2562 (
      {stage2_1[21]},
      {stage3_1[16]}
   );
   gpc1_1 gpc2563 (
      {stage2_1[22]},
      {stage3_1[17]}
   );
   gpc1_1 gpc2564 (
      {stage2_1[23]},
      {stage3_1[18]}
   );
   gpc1_1 gpc2565 (
      {stage2_1[24]},
      {stage3_1[19]}
   );
   gpc1_1 gpc2566 (
      {stage2_1[25]},
      {stage3_1[20]}
   );
   gpc1_1 gpc2567 (
      {stage2_1[26]},
      {stage3_1[21]}
   );
   gpc1_1 gpc2568 (
      {stage2_1[27]},
      {stage3_1[22]}
   );
   gpc1_1 gpc2569 (
      {stage2_1[28]},
      {stage3_1[23]}
   );
   gpc1_1 gpc2570 (
      {stage2_1[29]},
      {stage3_1[24]}
   );
   gpc1_1 gpc2571 (
      {stage2_1[30]},
      {stage3_1[25]}
   );
   gpc1_1 gpc2572 (
      {stage2_1[31]},
      {stage3_1[26]}
   );
   gpc1_1 gpc2573 (
      {stage2_1[32]},
      {stage3_1[27]}
   );
   gpc1_1 gpc2574 (
      {stage2_2[15]},
      {stage3_2[5]}
   );
   gpc1_1 gpc2575 (
      {stage2_2[16]},
      {stage3_2[6]}
   );
   gpc1_1 gpc2576 (
      {stage2_2[17]},
      {stage3_2[7]}
   );
   gpc1_1 gpc2577 (
      {stage2_2[18]},
      {stage3_2[8]}
   );
   gpc1_1 gpc2578 (
      {stage2_2[19]},
      {stage3_2[9]}
   );
   gpc1_1 gpc2579 (
      {stage2_2[20]},
      {stage3_2[10]}
   );
   gpc1_1 gpc2580 (
      {stage2_2[21]},
      {stage3_2[11]}
   );
   gpc1_1 gpc2581 (
      {stage2_2[22]},
      {stage3_2[12]}
   );
   gpc1_1 gpc2582 (
      {stage2_2[23]},
      {stage3_2[13]}
   );
   gpc1_1 gpc2583 (
      {stage2_2[24]},
      {stage3_2[14]}
   );
   gpc1_1 gpc2584 (
      {stage2_2[25]},
      {stage3_2[15]}
   );
   gpc1_1 gpc2585 (
      {stage2_2[26]},
      {stage3_2[16]}
   );
   gpc1_1 gpc2586 (
      {stage2_2[27]},
      {stage3_2[17]}
   );
   gpc1_1 gpc2587 (
      {stage2_2[28]},
      {stage3_2[18]}
   );
   gpc1_1 gpc2588 (
      {stage2_2[29]},
      {stage3_2[19]}
   );
   gpc1_1 gpc2589 (
      {stage2_2[30]},
      {stage3_2[20]}
   );
   gpc1_1 gpc2590 (
      {stage2_2[31]},
      {stage3_2[21]}
   );
   gpc1_1 gpc2591 (
      {stage2_2[32]},
      {stage3_2[22]}
   );
   gpc1_1 gpc2592 (
      {stage2_2[33]},
      {stage3_2[23]}
   );
   gpc1_1 gpc2593 (
      {stage2_2[34]},
      {stage3_2[24]}
   );
   gpc1_1 gpc2594 (
      {stage2_3[16]},
      {stage3_3[8]}
   );
   gpc1_1 gpc2595 (
      {stage2_3[17]},
      {stage3_3[9]}
   );
   gpc1_1 gpc2596 (
      {stage2_3[18]},
      {stage3_3[10]}
   );
   gpc1_1 gpc2597 (
      {stage2_3[19]},
      {stage3_3[11]}
   );
   gpc1_1 gpc2598 (
      {stage2_3[20]},
      {stage3_3[12]}
   );
   gpc1_1 gpc2599 (
      {stage2_3[21]},
      {stage3_3[13]}
   );
   gpc1_1 gpc2600 (
      {stage2_3[22]},
      {stage3_3[14]}
   );
   gpc1_1 gpc2601 (
      {stage2_3[23]},
      {stage3_3[15]}
   );
   gpc1_1 gpc2602 (
      {stage2_3[24]},
      {stage3_3[16]}
   );
   gpc1_1 gpc2603 (
      {stage2_3[25]},
      {stage3_3[17]}
   );
   gpc1_1 gpc2604 (
      {stage2_3[26]},
      {stage3_3[18]}
   );
   gpc1_1 gpc2605 (
      {stage2_3[27]},
      {stage3_3[19]}
   );
   gpc1_1 gpc2606 (
      {stage2_3[28]},
      {stage3_3[20]}
   );
   gpc1_1 gpc2607 (
      {stage2_3[29]},
      {stage3_3[21]}
   );
   gpc1_1 gpc2608 (
      {stage2_3[30]},
      {stage3_3[22]}
   );
   gpc1_1 gpc2609 (
      {stage2_3[31]},
      {stage3_3[23]}
   );
   gpc1_1 gpc2610 (
      {stage2_3[32]},
      {stage3_3[24]}
   );
   gpc1_1 gpc2611 (
      {stage2_3[33]},
      {stage3_3[25]}
   );
   gpc1_1 gpc2612 (
      {stage2_3[34]},
      {stage3_3[26]}
   );
   gpc1_1 gpc2613 (
      {stage2_3[35]},
      {stage3_3[27]}
   );
   gpc1_1 gpc2614 (
      {stage2_3[36]},
      {stage3_3[28]}
   );
   gpc1_1 gpc2615 (
      {stage2_3[37]},
      {stage3_3[29]}
   );
   gpc1_1 gpc2616 (
      {stage2_3[38]},
      {stage3_3[30]}
   );
   gpc1_1 gpc2617 (
      {stage2_3[39]},
      {stage3_3[31]}
   );
   gpc1_1 gpc2618 (
      {stage2_3[40]},
      {stage3_3[32]}
   );
   gpc1_1 gpc2619 (
      {stage2_3[41]},
      {stage3_3[33]}
   );
   gpc1_1 gpc2620 (
      {stage2_3[42]},
      {stage3_3[34]}
   );
   gpc1_1 gpc2621 (
      {stage2_4[52]},
      {stage3_4[14]}
   );
   gpc1_1 gpc2622 (
      {stage2_4[53]},
      {stage3_4[15]}
   );
   gpc1_1 gpc2623 (
      {stage2_4[54]},
      {stage3_4[16]}
   );
   gpc1_1 gpc2624 (
      {stage2_4[55]},
      {stage3_4[17]}
   );
   gpc1_1 gpc2625 (
      {stage2_4[56]},
      {stage3_4[18]}
   );
   gpc1_1 gpc2626 (
      {stage2_4[57]},
      {stage3_4[19]}
   );
   gpc1_1 gpc2627 (
      {stage2_4[58]},
      {stage3_4[20]}
   );
   gpc1_1 gpc2628 (
      {stage2_4[59]},
      {stage3_4[21]}
   );
   gpc1_1 gpc2629 (
      {stage2_4[60]},
      {stage3_4[22]}
   );
   gpc1_1 gpc2630 (
      {stage2_4[61]},
      {stage3_4[23]}
   );
   gpc1_1 gpc2631 (
      {stage2_4[62]},
      {stage3_4[24]}
   );
   gpc1_1 gpc2632 (
      {stage2_4[63]},
      {stage3_4[25]}
   );
   gpc1_1 gpc2633 (
      {stage2_4[64]},
      {stage3_4[26]}
   );
   gpc1_1 gpc2634 (
      {stage2_4[65]},
      {stage3_4[27]}
   );
   gpc1_1 gpc2635 (
      {stage2_4[66]},
      {stage3_4[28]}
   );
   gpc1_1 gpc2636 (
      {stage2_4[67]},
      {stage3_4[29]}
   );
   gpc1_1 gpc2637 (
      {stage2_4[68]},
      {stage3_4[30]}
   );
   gpc1_1 gpc2638 (
      {stage2_4[69]},
      {stage3_4[31]}
   );
   gpc1_1 gpc2639 (
      {stage2_4[70]},
      {stage3_4[32]}
   );
   gpc1_1 gpc2640 (
      {stage2_4[71]},
      {stage3_4[33]}
   );
   gpc1_1 gpc2641 (
      {stage2_4[72]},
      {stage3_4[34]}
   );
   gpc1_1 gpc2642 (
      {stage2_4[73]},
      {stage3_4[35]}
   );
   gpc1_1 gpc2643 (
      {stage2_5[41]},
      {stage3_5[15]}
   );
   gpc1_1 gpc2644 (
      {stage2_6[48]},
      {stage3_6[15]}
   );
   gpc1_1 gpc2645 (
      {stage2_6[49]},
      {stage3_6[16]}
   );
   gpc1_1 gpc2646 (
      {stage2_6[50]},
      {stage3_6[17]}
   );
   gpc1_1 gpc2647 (
      {stage2_6[51]},
      {stage3_6[18]}
   );
   gpc1_1 gpc2648 (
      {stage2_6[52]},
      {stage3_6[19]}
   );
   gpc1_1 gpc2649 (
      {stage2_7[51]},
      {stage3_7[21]}
   );
   gpc1_1 gpc2650 (
      {stage2_7[52]},
      {stage3_7[22]}
   );
   gpc1_1 gpc2651 (
      {stage2_7[53]},
      {stage3_7[23]}
   );
   gpc1_1 gpc2652 (
      {stage2_8[55]},
      {stage3_8[26]}
   );
   gpc1_1 gpc2653 (
      {stage2_12[73]},
      {stage3_12[30]}
   );
   gpc1_1 gpc2654 (
      {stage2_12[74]},
      {stage3_12[31]}
   );
   gpc1_1 gpc2655 (
      {stage2_13[42]},
      {stage3_13[22]}
   );
   gpc1_1 gpc2656 (
      {stage2_13[43]},
      {stage3_13[23]}
   );
   gpc1_1 gpc2657 (
      {stage2_13[44]},
      {stage3_13[24]}
   );
   gpc1_1 gpc2658 (
      {stage2_13[45]},
      {stage3_13[25]}
   );
   gpc1_1 gpc2659 (
      {stage2_13[46]},
      {stage3_13[26]}
   );
   gpc1_1 gpc2660 (
      {stage2_13[47]},
      {stage3_13[27]}
   );
   gpc1_1 gpc2661 (
      {stage2_13[48]},
      {stage3_13[28]}
   );
   gpc1_1 gpc2662 (
      {stage2_13[49]},
      {stage3_13[29]}
   );
   gpc1_1 gpc2663 (
      {stage2_13[50]},
      {stage3_13[30]}
   );
   gpc1_1 gpc2664 (
      {stage2_13[51]},
      {stage3_13[31]}
   );
   gpc1_1 gpc2665 (
      {stage2_13[52]},
      {stage3_13[32]}
   );
   gpc1_1 gpc2666 (
      {stage2_13[53]},
      {stage3_13[33]}
   );
   gpc1_1 gpc2667 (
      {stage2_13[54]},
      {stage3_13[34]}
   );
   gpc1_1 gpc2668 (
      {stage2_13[55]},
      {stage3_13[35]}
   );
   gpc1_1 gpc2669 (
      {stage2_13[56]},
      {stage3_13[36]}
   );
   gpc1_1 gpc2670 (
      {stage2_14[86]},
      {stage3_14[22]}
   );
   gpc1_1 gpc2671 (
      {stage2_14[87]},
      {stage3_14[23]}
   );
   gpc1_1 gpc2672 (
      {stage2_14[88]},
      {stage3_14[24]}
   );
   gpc1_1 gpc2673 (
      {stage2_14[89]},
      {stage3_14[25]}
   );
   gpc1_1 gpc2674 (
      {stage2_15[44]},
      {stage3_15[30]}
   );
   gpc1_1 gpc2675 (
      {stage2_15[45]},
      {stage3_15[31]}
   );
   gpc1_1 gpc2676 (
      {stage2_15[46]},
      {stage3_15[32]}
   );
   gpc1_1 gpc2677 (
      {stage2_16[38]},
      {stage3_16[24]}
   );
   gpc1_1 gpc2678 (
      {stage2_16[39]},
      {stage3_16[25]}
   );
   gpc1_1 gpc2679 (
      {stage2_16[40]},
      {stage3_16[26]}
   );
   gpc1_1 gpc2680 (
      {stage2_17[48]},
      {stage3_17[13]}
   );
   gpc1_1 gpc2681 (
      {stage2_17[49]},
      {stage3_17[14]}
   );
   gpc1_1 gpc2682 (
      {stage2_17[50]},
      {stage3_17[15]}
   );
   gpc1_1 gpc2683 (
      {stage2_17[51]},
      {stage3_17[16]}
   );
   gpc1_1 gpc2684 (
      {stage2_17[52]},
      {stage3_17[17]}
   );
   gpc1_1 gpc2685 (
      {stage2_17[53]},
      {stage3_17[18]}
   );
   gpc1_1 gpc2686 (
      {stage2_17[54]},
      {stage3_17[19]}
   );
   gpc1_1 gpc2687 (
      {stage2_18[81]},
      {stage3_18[28]}
   );
   gpc1_1 gpc2688 (
      {stage2_18[82]},
      {stage3_18[29]}
   );
   gpc1_1 gpc2689 (
      {stage2_18[83]},
      {stage3_18[30]}
   );
   gpc1_1 gpc2690 (
      {stage2_18[84]},
      {stage3_18[31]}
   );
   gpc1_1 gpc2691 (
      {stage2_18[85]},
      {stage3_18[32]}
   );
   gpc1_1 gpc2692 (
      {stage2_18[86]},
      {stage3_18[33]}
   );
   gpc1_1 gpc2693 (
      {stage2_18[87]},
      {stage3_18[34]}
   );
   gpc1_1 gpc2694 (
      {stage2_18[88]},
      {stage3_18[35]}
   );
   gpc1_1 gpc2695 (
      {stage2_18[89]},
      {stage3_18[36]}
   );
   gpc1_1 gpc2696 (
      {stage2_18[90]},
      {stage3_18[37]}
   );
   gpc1_1 gpc2697 (
      {stage2_19[40]},
      {stage3_19[29]}
   );
   gpc1_1 gpc2698 (
      {stage2_19[41]},
      {stage3_19[30]}
   );
   gpc1_1 gpc2699 (
      {stage2_19[42]},
      {stage3_19[31]}
   );
   gpc1_1 gpc2700 (
      {stage2_19[43]},
      {stage3_19[32]}
   );
   gpc1_1 gpc2701 (
      {stage2_19[44]},
      {stage3_19[33]}
   );
   gpc1_1 gpc2702 (
      {stage2_19[45]},
      {stage3_19[34]}
   );
   gpc1_1 gpc2703 (
      {stage2_20[113]},
      {stage3_20[24]}
   );
   gpc1_1 gpc2704 (
      {stage2_20[114]},
      {stage3_20[25]}
   );
   gpc1_1 gpc2705 (
      {stage2_20[115]},
      {stage3_20[26]}
   );
   gpc1_1 gpc2706 (
      {stage2_20[116]},
      {stage3_20[27]}
   );
   gpc1_1 gpc2707 (
      {stage2_20[117]},
      {stage3_20[28]}
   );
   gpc1_1 gpc2708 (
      {stage2_20[118]},
      {stage3_20[29]}
   );
   gpc1_1 gpc2709 (
      {stage2_20[119]},
      {stage3_20[30]}
   );
   gpc1_1 gpc2710 (
      {stage2_20[120]},
      {stage3_20[31]}
   );
   gpc1_1 gpc2711 (
      {stage2_20[121]},
      {stage3_20[32]}
   );
   gpc1_1 gpc2712 (
      {stage2_20[122]},
      {stage3_20[33]}
   );
   gpc1_1 gpc2713 (
      {stage2_20[123]},
      {stage3_20[34]}
   );
   gpc1_1 gpc2714 (
      {stage2_20[124]},
      {stage3_20[35]}
   );
   gpc1_1 gpc2715 (
      {stage2_20[125]},
      {stage3_20[36]}
   );
   gpc1_1 gpc2716 (
      {stage2_25[60]},
      {stage3_25[30]}
   );
   gpc1_1 gpc2717 (
      {stage2_25[61]},
      {stage3_25[31]}
   );
   gpc1_1 gpc2718 (
      {stage2_25[62]},
      {stage3_25[32]}
   );
   gpc1_1 gpc2719 (
      {stage2_25[63]},
      {stage3_25[33]}
   );
   gpc1_1 gpc2720 (
      {stage2_25[64]},
      {stage3_25[34]}
   );
   gpc1_1 gpc2721 (
      {stage2_25[65]},
      {stage3_25[35]}
   );
   gpc1_1 gpc2722 (
      {stage2_27[84]},
      {stage3_27[27]}
   );
   gpc1_1 gpc2723 (
      {stage2_27[85]},
      {stage3_27[28]}
   );
   gpc1_1 gpc2724 (
      {stage2_27[86]},
      {stage3_27[29]}
   );
   gpc1_1 gpc2725 (
      {stage2_27[87]},
      {stage3_27[30]}
   );
   gpc1_1 gpc2726 (
      {stage2_27[88]},
      {stage3_27[31]}
   );
   gpc1_1 gpc2727 (
      {stage2_27[89]},
      {stage3_27[32]}
   );
   gpc1_1 gpc2728 (
      {stage2_27[90]},
      {stage3_27[33]}
   );
   gpc1_1 gpc2729 (
      {stage2_27[91]},
      {stage3_27[34]}
   );
   gpc1_1 gpc2730 (
      {stage2_27[92]},
      {stage3_27[35]}
   );
   gpc1_1 gpc2731 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc2732 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc2733 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc2734 (
      {stage2_28[58]},
      {stage3_28[31]}
   );
   gpc1_1 gpc2735 (
      {stage2_28[59]},
      {stage3_28[32]}
   );
   gpc1_1 gpc2736 (
      {stage2_28[60]},
      {stage3_28[33]}
   );
   gpc1_1 gpc2737 (
      {stage2_28[61]},
      {stage3_28[34]}
   );
   gpc1_1 gpc2738 (
      {stage2_28[62]},
      {stage3_28[35]}
   );
   gpc1_1 gpc2739 (
      {stage2_28[63]},
      {stage3_28[36]}
   );
   gpc1_1 gpc2740 (
      {stage2_28[64]},
      {stage3_28[37]}
   );
   gpc1_1 gpc2741 (
      {stage2_28[65]},
      {stage3_28[38]}
   );
   gpc1_1 gpc2742 (
      {stage2_28[66]},
      {stage3_28[39]}
   );
   gpc1_1 gpc2743 (
      {stage2_28[67]},
      {stage3_28[40]}
   );
   gpc1_1 gpc2744 (
      {stage2_28[68]},
      {stage3_28[41]}
   );
   gpc1_1 gpc2745 (
      {stage2_28[69]},
      {stage3_28[42]}
   );
   gpc1_1 gpc2746 (
      {stage2_28[70]},
      {stage3_28[43]}
   );
   gpc1_1 gpc2747 (
      {stage2_28[71]},
      {stage3_28[44]}
   );
   gpc1_1 gpc2748 (
      {stage2_29[36]},
      {stage3_29[24]}
   );
   gpc1_1 gpc2749 (
      {stage2_29[37]},
      {stage3_29[25]}
   );
   gpc1_1 gpc2750 (
      {stage2_29[38]},
      {stage3_29[26]}
   );
   gpc1_1 gpc2751 (
      {stage2_29[39]},
      {stage3_29[27]}
   );
   gpc1_1 gpc2752 (
      {stage2_31[29]},
      {stage3_31[18]}
   );
   gpc1_1 gpc2753 (
      {stage2_31[30]},
      {stage3_31[19]}
   );
   gpc1_1 gpc2754 (
      {stage2_31[31]},
      {stage3_31[20]}
   );
   gpc1_1 gpc2755 (
      {stage2_31[32]},
      {stage3_31[21]}
   );
   gpc1_1 gpc2756 (
      {stage2_31[33]},
      {stage3_31[22]}
   );
   gpc1_1 gpc2757 (
      {stage2_31[34]},
      {stage3_31[23]}
   );
   gpc1_1 gpc2758 (
      {stage2_31[35]},
      {stage3_31[24]}
   );
   gpc1_1 gpc2759 (
      {stage2_31[36]},
      {stage3_31[25]}
   );
   gpc1_1 gpc2760 (
      {stage2_31[37]},
      {stage3_31[26]}
   );
   gpc1_1 gpc2761 (
      {stage2_31[38]},
      {stage3_31[27]}
   );
   gpc1_1 gpc2762 (
      {stage2_31[39]},
      {stage3_31[28]}
   );
   gpc1_1 gpc2763 (
      {stage2_31[40]},
      {stage3_31[29]}
   );
   gpc1_1 gpc2764 (
      {stage2_31[41]},
      {stage3_31[30]}
   );
   gpc1_1 gpc2765 (
      {stage2_31[42]},
      {stage3_31[31]}
   );
   gpc1_1 gpc2766 (
      {stage2_31[43]},
      {stage3_31[32]}
   );
   gpc1_1 gpc2767 (
      {stage2_31[44]},
      {stage3_31[33]}
   );
   gpc1_1 gpc2768 (
      {stage2_31[45]},
      {stage3_31[34]}
   );
   gpc1_1 gpc2769 (
      {stage2_31[46]},
      {stage3_31[35]}
   );
   gpc1_1 gpc2770 (
      {stage2_31[47]},
      {stage3_31[36]}
   );
   gpc1_1 gpc2771 (
      {stage2_32[40]},
      {stage3_32[16]}
   );
   gpc1_1 gpc2772 (
      {stage2_32[41]},
      {stage3_32[17]}
   );
   gpc1_1 gpc2773 (
      {stage2_32[42]},
      {stage3_32[18]}
   );
   gpc1_1 gpc2774 (
      {stage2_32[43]},
      {stage3_32[19]}
   );
   gpc1_1 gpc2775 (
      {stage2_33[24]},
      {stage3_33[11]}
   );
   gpc1_1 gpc2776 (
      {stage2_33[25]},
      {stage3_33[12]}
   );
   gpc1_1 gpc2777 (
      {stage2_33[26]},
      {stage3_33[13]}
   );
   gpc1_1 gpc2778 (
      {stage2_33[27]},
      {stage3_33[14]}
   );
   gpc1_1 gpc2779 (
      {stage2_33[28]},
      {stage3_33[15]}
   );
   gpc1_1 gpc2780 (
      {stage2_33[29]},
      {stage3_33[16]}
   );
   gpc1_1 gpc2781 (
      {stage2_33[30]},
      {stage3_33[17]}
   );
   gpc1_1 gpc2782 (
      {stage2_35[0]},
      {stage3_35[7]}
   );
   gpc1_1 gpc2783 (
      {stage2_35[1]},
      {stage3_35[8]}
   );
   gpc1_1 gpc2784 (
      {stage2_35[2]},
      {stage3_35[9]}
   );
   gpc1_1 gpc2785 (
      {stage2_35[3]},
      {stage3_35[10]}
   );
   gpc1_1 gpc2786 (
      {stage2_35[4]},
      {stage3_35[11]}
   );
   gpc1_1 gpc2787 (
      {stage2_35[5]},
      {stage3_35[12]}
   );
   gpc606_5 gpc2788 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc2789 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc2790 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc2791 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc2792 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc2793 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc2794 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc207_4 gpc2795 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_5[0], stage3_5[1]},
      {stage4_6[4],stage4_5[7],stage4_4[7],stage4_3[7]}
   );
   gpc207_4 gpc2796 (
      {stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30], stage3_3[31]},
      {stage3_5[2], stage3_5[3]},
      {stage4_6[5],stage4_5[8],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc2797 (
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[6],stage4_5[9],stage4_4[9]}
   );
   gpc606_5 gpc2798 (
      {stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc2799 (
      {stage3_5[10], stage3_5[11], stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[8],stage4_5[11]}
   );
   gpc615_5 gpc2800 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[12]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[2],stage4_8[3],stage4_7[3],stage4_6[9]}
   );
   gpc615_5 gpc2801 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[13]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[3],stage4_8[4],stage4_7[4],stage4_6[10]}
   );
   gpc135_4 gpc2802 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc2803 (
      {stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[3],stage4_9[5],stage4_8[6]}
   );
   gpc135_4 gpc2804 (
      {stage3_8[22], stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26]},
      {stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[2]},
      {stage4_11[2],stage4_10[4],stage4_9[6],stage4_8[7]}
   );
   gpc606_5 gpc2805 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[7]}
   );
   gpc606_5 gpc2806 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[4],stage4_10[6],stage4_9[8]}
   );
   gpc615_5 gpc2807 (
      {stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[5],stage4_10[7]}
   );
   gpc615_5 gpc2808 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[6],stage4_10[8]}
   );
   gpc615_5 gpc2809 (
      {stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17], stage3_11[18]},
      {stage3_12[12]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[2],stage4_13[4],stage4_12[4],stage4_11[7]}
   );
   gpc615_5 gpc2810 (
      {stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage3_12[13]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[3],stage4_13[5],stage4_12[5],stage4_11[8]}
   );
   gpc615_5 gpc2811 (
      {stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18]},
      {stage3_13[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[4],stage4_13[6],stage4_12[6]}
   );
   gpc615_5 gpc2812 (
      {stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[13]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[5],stage4_13[7],stage4_12[7]}
   );
   gpc615_5 gpc2813 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_13[14]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[4],stage4_14[6],stage4_13[8],stage4_12[8]}
   );
   gpc606_5 gpc2814 (
      {stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[3],stage4_15[5],stage4_14[7],stage4_13[9]}
   );
   gpc606_5 gpc2815 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[4],stage4_15[6],stage4_14[8],stage4_13[10]}
   );
   gpc606_5 gpc2816 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[5],stage4_15[7],stage4_14[9]}
   );
   gpc615_5 gpc2817 (
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16]},
      {stage3_16[6]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[3],stage4_16[6],stage4_15[8]}
   );
   gpc615_5 gpc2818 (
      {stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage3_16[7]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[2],stage4_17[4],stage4_16[7],stage4_15[9]}
   );
   gpc615_5 gpc2819 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[8]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[3],stage4_17[5],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc2820 (
      {stage3_16[9], stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13]},
      {stage3_17[18]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[4],stage4_17[6],stage4_16[9]}
   );
   gpc615_5 gpc2821 (
      {stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[19]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[5],stage4_17[7],stage4_16[10]}
   );
   gpc1163_5 gpc2822 (
      {stage3_18[12], stage3_18[13], stage3_18[14]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[0]},
      {stage3_21[0]},
      {stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[6]}
   );
   gpc1163_5 gpc2823 (
      {stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage3_20[1]},
      {stage3_21[1]},
      {stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[7]}
   );
   gpc1163_5 gpc2824 (
      {stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage3_20[2]},
      {stage3_21[2]},
      {stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[7],stage4_18[8]}
   );
   gpc615_5 gpc2825 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage3_19[18]},
      {stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8]},
      {stage4_22[3],stage4_21[3],stage4_20[5],stage4_19[8],stage4_18[9]}
   );
   gpc615_5 gpc2826 (
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30]},
      {stage3_19[19]},
      {stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14]},
      {stage4_22[4],stage4_21[4],stage4_20[6],stage4_19[9],stage4_18[10]}
   );
   gpc615_5 gpc2827 (
      {stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35]},
      {stage3_19[20]},
      {stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20]},
      {stage4_22[5],stage4_21[5],stage4_20[7],stage4_19[10],stage4_18[11]}
   );
   gpc615_5 gpc2828 (
      {stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_20[21]},
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage4_23[0],stage4_22[6],stage4_21[6],stage4_20[8],stage4_19[11]}
   );
   gpc615_5 gpc2829 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[22]},
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage4_23[1],stage4_22[7],stage4_21[7],stage4_20[9],stage4_19[12]}
   );
   gpc615_5 gpc2830 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], 1'b0},
      {stage3_20[23]},
      {stage3_21[15], stage3_21[16], stage3_21[17], stage3_21[18], stage3_21[19], stage3_21[20]},
      {stage4_23[2],stage4_22[8],stage4_21[8],stage4_20[10],stage4_19[13]}
   );
   gpc606_5 gpc2831 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[3],stage4_22[9],stage4_21[9],stage4_20[11]}
   );
   gpc606_5 gpc2832 (
      {stage3_21[21], stage3_21[22], stage3_21[23], stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[1],stage4_23[4],stage4_22[10],stage4_21[10]}
   );
   gpc606_5 gpc2833 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[2],stage4_23[5],stage4_22[11],stage4_21[11]}
   );
   gpc615_5 gpc2834 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[12]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[2],stage4_24[3],stage4_23[6],stage4_22[12]}
   );
   gpc615_5 gpc2835 (
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15]},
      {stage3_23[13]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[3],stage4_24[4],stage4_23[7],stage4_22[13]}
   );
   gpc615_5 gpc2836 (
      {stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20]},
      {stage3_23[14]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[4],stage4_24[5],stage4_23[8],stage4_22[14]}
   );
   gpc615_5 gpc2837 (
      {stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25]},
      {stage3_23[15]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[5],stage4_24[6],stage4_23[9],stage4_22[15]}
   );
   gpc615_5 gpc2838 (
      {stage3_23[16], stage3_23[17], stage3_23[18], stage3_23[19], stage3_23[20]},
      {1'b0},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[6],stage4_24[7],stage4_23[10]}
   );
   gpc606_5 gpc2839 (
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[5],stage4_25[7]}
   );
   gpc606_5 gpc2840 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[2],stage4_26[6],stage4_25[8]}
   );
   gpc606_5 gpc2841 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[3],stage4_26[7],stage4_25[9]}
   );
   gpc606_5 gpc2842 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[3],stage4_27[4],stage4_26[8],stage4_25[10]}
   );
   gpc606_5 gpc2843 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage4_29[4],stage4_28[4],stage4_27[5],stage4_26[9],stage4_25[11]}
   );
   gpc606_5 gpc2844 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[5],stage4_28[5],stage4_27[6],stage4_26[10]}
   );
   gpc606_5 gpc2845 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[6],stage4_28[6],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc2846 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16]},
      {stage3_27[30]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[7],stage4_28[7],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc2847 (
      {stage3_26[17], stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21]},
      {stage3_27[31]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[8],stage4_28[8],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc2848 (
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[0],stage4_30[4],stage4_29[9],stage4_28[9]}
   );
   gpc606_5 gpc2849 (
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[1],stage4_30[5],stage4_29[10],stage4_28[10]}
   );
   gpc606_5 gpc2850 (
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[6],stage4_29[11]}
   );
   gpc606_5 gpc2851 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[3],stage4_30[7],stage4_29[12]}
   );
   gpc606_5 gpc2852 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[4],stage4_30[8],stage4_29[13]}
   );
   gpc606_5 gpc2853 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[5],stage4_30[9]}
   );
   gpc615_5 gpc2854 (
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage3_32[6]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6],stage4_31[6]}
   );
   gpc615_5 gpc2855 (
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage3_32[7]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7],stage4_31[7]}
   );
   gpc606_5 gpc2856 (
      {stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc2857 (
      {stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], 1'b0, 1'b0},
      {stage4_36[1],stage4_35[3],stage4_34[4],stage4_33[7],stage4_32[9]}
   );
   gpc606_5 gpc2858 (
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1_1 gpc2859 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc2860 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc2861 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc2862 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc2863 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc2864 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc2865 (
      {stage3_1[18]},
      {stage4_1[3]}
   );
   gpc1_1 gpc2866 (
      {stage3_1[19]},
      {stage4_1[4]}
   );
   gpc1_1 gpc2867 (
      {stage3_1[20]},
      {stage4_1[5]}
   );
   gpc1_1 gpc2868 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc2869 (
      {stage3_1[22]},
      {stage4_1[7]}
   );
   gpc1_1 gpc2870 (
      {stage3_1[23]},
      {stage4_1[8]}
   );
   gpc1_1 gpc2871 (
      {stage3_1[24]},
      {stage4_1[9]}
   );
   gpc1_1 gpc2872 (
      {stage3_1[25]},
      {stage4_1[10]}
   );
   gpc1_1 gpc2873 (
      {stage3_1[26]},
      {stage4_1[11]}
   );
   gpc1_1 gpc2874 (
      {stage3_1[27]},
      {stage4_1[12]}
   );
   gpc1_1 gpc2875 (
      {stage3_2[24]},
      {stage4_2[7]}
   );
   gpc1_1 gpc2876 (
      {stage3_3[32]},
      {stage4_3[9]}
   );
   gpc1_1 gpc2877 (
      {stage3_3[33]},
      {stage4_3[10]}
   );
   gpc1_1 gpc2878 (
      {stage3_3[34]},
      {stage4_3[11]}
   );
   gpc1_1 gpc2879 (
      {stage3_4[30]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2880 (
      {stage3_4[31]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2881 (
      {stage3_4[32]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2882 (
      {stage3_4[33]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2883 (
      {stage3_4[34]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2884 (
      {stage3_4[35]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2885 (
      {stage3_6[16]},
      {stage4_6[11]}
   );
   gpc1_1 gpc2886 (
      {stage3_6[17]},
      {stage4_6[12]}
   );
   gpc1_1 gpc2887 (
      {stage3_6[18]},
      {stage4_6[13]}
   );
   gpc1_1 gpc2888 (
      {stage3_6[19]},
      {stage4_6[14]}
   );
   gpc1_1 gpc2889 (
      {stage3_7[14]},
      {stage4_7[5]}
   );
   gpc1_1 gpc2890 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc2891 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc2892 (
      {stage3_7[17]},
      {stage4_7[8]}
   );
   gpc1_1 gpc2893 (
      {stage3_7[18]},
      {stage4_7[9]}
   );
   gpc1_1 gpc2894 (
      {stage3_7[19]},
      {stage4_7[10]}
   );
   gpc1_1 gpc2895 (
      {stage3_7[20]},
      {stage4_7[11]}
   );
   gpc1_1 gpc2896 (
      {stage3_7[21]},
      {stage4_7[12]}
   );
   gpc1_1 gpc2897 (
      {stage3_7[22]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2898 (
      {stage3_7[23]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2899 (
      {stage3_9[21]},
      {stage4_9[9]}
   );
   gpc1_1 gpc2900 (
      {stage3_10[13]},
      {stage4_10[9]}
   );
   gpc1_1 gpc2901 (
      {stage3_10[14]},
      {stage4_10[10]}
   );
   gpc1_1 gpc2902 (
      {stage3_10[15]},
      {stage4_10[11]}
   );
   gpc1_1 gpc2903 (
      {stage3_10[16]},
      {stage4_10[12]}
   );
   gpc1_1 gpc2904 (
      {stage3_10[17]},
      {stage4_10[13]}
   );
   gpc1_1 gpc2905 (
      {stage3_10[18]},
      {stage4_10[14]}
   );
   gpc1_1 gpc2906 (
      {stage3_11[24]},
      {stage4_11[9]}
   );
   gpc1_1 gpc2907 (
      {stage3_11[25]},
      {stage4_11[10]}
   );
   gpc1_1 gpc2908 (
      {stage3_12[29]},
      {stage4_12[9]}
   );
   gpc1_1 gpc2909 (
      {stage3_12[30]},
      {stage4_12[10]}
   );
   gpc1_1 gpc2910 (
      {stage3_12[31]},
      {stage4_12[11]}
   );
   gpc1_1 gpc2911 (
      {stage3_13[27]},
      {stage4_13[11]}
   );
   gpc1_1 gpc2912 (
      {stage3_13[28]},
      {stage4_13[12]}
   );
   gpc1_1 gpc2913 (
      {stage3_13[29]},
      {stage4_13[13]}
   );
   gpc1_1 gpc2914 (
      {stage3_13[30]},
      {stage4_13[14]}
   );
   gpc1_1 gpc2915 (
      {stage3_13[31]},
      {stage4_13[15]}
   );
   gpc1_1 gpc2916 (
      {stage3_13[32]},
      {stage4_13[16]}
   );
   gpc1_1 gpc2917 (
      {stage3_13[33]},
      {stage4_13[17]}
   );
   gpc1_1 gpc2918 (
      {stage3_13[34]},
      {stage4_13[18]}
   );
   gpc1_1 gpc2919 (
      {stage3_13[35]},
      {stage4_13[19]}
   );
   gpc1_1 gpc2920 (
      {stage3_13[36]},
      {stage4_13[20]}
   );
   gpc1_1 gpc2921 (
      {stage3_14[24]},
      {stage4_14[10]}
   );
   gpc1_1 gpc2922 (
      {stage3_14[25]},
      {stage4_14[11]}
   );
   gpc1_1 gpc2923 (
      {stage3_15[27]},
      {stage4_15[11]}
   );
   gpc1_1 gpc2924 (
      {stage3_15[28]},
      {stage4_15[12]}
   );
   gpc1_1 gpc2925 (
      {stage3_15[29]},
      {stage4_15[13]}
   );
   gpc1_1 gpc2926 (
      {stage3_15[30]},
      {stage4_15[14]}
   );
   gpc1_1 gpc2927 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc2928 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc2929 (
      {stage3_16[19]},
      {stage4_16[11]}
   );
   gpc1_1 gpc2930 (
      {stage3_16[20]},
      {stage4_16[12]}
   );
   gpc1_1 gpc2931 (
      {stage3_16[21]},
      {stage4_16[13]}
   );
   gpc1_1 gpc2932 (
      {stage3_16[22]},
      {stage4_16[14]}
   );
   gpc1_1 gpc2933 (
      {stage3_16[23]},
      {stage4_16[15]}
   );
   gpc1_1 gpc2934 (
      {stage3_16[24]},
      {stage4_16[16]}
   );
   gpc1_1 gpc2935 (
      {stage3_16[25]},
      {stage4_16[17]}
   );
   gpc1_1 gpc2936 (
      {stage3_16[26]},
      {stage4_16[18]}
   );
   gpc1_1 gpc2937 (
      {stage3_18[36]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2938 (
      {stage3_18[37]},
      {stage4_18[13]}
   );
   gpc1_1 gpc2939 (
      {stage3_20[30]},
      {stage4_20[12]}
   );
   gpc1_1 gpc2940 (
      {stage3_20[31]},
      {stage4_20[13]}
   );
   gpc1_1 gpc2941 (
      {stage3_20[32]},
      {stage4_20[14]}
   );
   gpc1_1 gpc2942 (
      {stage3_20[33]},
      {stage4_20[15]}
   );
   gpc1_1 gpc2943 (
      {stage3_20[34]},
      {stage4_20[16]}
   );
   gpc1_1 gpc2944 (
      {stage3_20[35]},
      {stage4_20[17]}
   );
   gpc1_1 gpc2945 (
      {stage3_20[36]},
      {stage4_20[18]}
   );
   gpc1_1 gpc2946 (
      {stage3_22[26]},
      {stage4_22[16]}
   );
   gpc1_1 gpc2947 (
      {stage3_22[27]},
      {stage4_22[17]}
   );
   gpc1_1 gpc2948 (
      {stage3_22[28]},
      {stage4_22[18]}
   );
   gpc1_1 gpc2949 (
      {stage3_22[29]},
      {stage4_22[19]}
   );
   gpc1_1 gpc2950 (
      {stage3_22[30]},
      {stage4_22[20]}
   );
   gpc1_1 gpc2951 (
      {stage3_22[31]},
      {stage4_22[21]}
   );
   gpc1_1 gpc2952 (
      {stage3_22[32]},
      {stage4_22[22]}
   );
   gpc1_1 gpc2953 (
      {stage3_22[33]},
      {stage4_22[23]}
   );
   gpc1_1 gpc2954 (
      {stage3_22[34]},
      {stage4_22[24]}
   );
   gpc1_1 gpc2955 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc2956 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc2957 (
      {stage3_27[32]},
      {stage4_27[10]}
   );
   gpc1_1 gpc2958 (
      {stage3_27[33]},
      {stage4_27[11]}
   );
   gpc1_1 gpc2959 (
      {stage3_27[34]},
      {stage4_27[12]}
   );
   gpc1_1 gpc2960 (
      {stage3_27[35]},
      {stage4_27[13]}
   );
   gpc1_1 gpc2961 (
      {stage3_27[36]},
      {stage4_27[14]}
   );
   gpc1_1 gpc2962 (
      {stage3_27[37]},
      {stage4_27[15]}
   );
   gpc1_1 gpc2963 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc2964 (
      {stage3_28[36]},
      {stage4_28[11]}
   );
   gpc1_1 gpc2965 (
      {stage3_28[37]},
      {stage4_28[12]}
   );
   gpc1_1 gpc2966 (
      {stage3_28[38]},
      {stage4_28[13]}
   );
   gpc1_1 gpc2967 (
      {stage3_28[39]},
      {stage4_28[14]}
   );
   gpc1_1 gpc2968 (
      {stage3_28[40]},
      {stage4_28[15]}
   );
   gpc1_1 gpc2969 (
      {stage3_28[41]},
      {stage4_28[16]}
   );
   gpc1_1 gpc2970 (
      {stage3_28[42]},
      {stage4_28[17]}
   );
   gpc1_1 gpc2971 (
      {stage3_28[43]},
      {stage4_28[18]}
   );
   gpc1_1 gpc2972 (
      {stage3_28[44]},
      {stage4_28[19]}
   );
   gpc1_1 gpc2973 (
      {stage3_29[18]},
      {stage4_29[14]}
   );
   gpc1_1 gpc2974 (
      {stage3_29[19]},
      {stage4_29[15]}
   );
   gpc1_1 gpc2975 (
      {stage3_29[20]},
      {stage4_29[16]}
   );
   gpc1_1 gpc2976 (
      {stage3_29[21]},
      {stage4_29[17]}
   );
   gpc1_1 gpc2977 (
      {stage3_29[22]},
      {stage4_29[18]}
   );
   gpc1_1 gpc2978 (
      {stage3_29[23]},
      {stage4_29[19]}
   );
   gpc1_1 gpc2979 (
      {stage3_29[24]},
      {stage4_29[20]}
   );
   gpc1_1 gpc2980 (
      {stage3_29[25]},
      {stage4_29[21]}
   );
   gpc1_1 gpc2981 (
      {stage3_29[26]},
      {stage4_29[22]}
   );
   gpc1_1 gpc2982 (
      {stage3_29[27]},
      {stage4_29[23]}
   );
   gpc1_1 gpc2983 (
      {stage3_31[28]},
      {stage4_31[8]}
   );
   gpc1_1 gpc2984 (
      {stage3_31[29]},
      {stage4_31[9]}
   );
   gpc1_1 gpc2985 (
      {stage3_31[30]},
      {stage4_31[10]}
   );
   gpc1_1 gpc2986 (
      {stage3_31[31]},
      {stage4_31[11]}
   );
   gpc1_1 gpc2987 (
      {stage3_31[32]},
      {stage4_31[12]}
   );
   gpc1_1 gpc2988 (
      {stage3_31[33]},
      {stage4_31[13]}
   );
   gpc1_1 gpc2989 (
      {stage3_31[34]},
      {stage4_31[14]}
   );
   gpc1_1 gpc2990 (
      {stage3_31[35]},
      {stage4_31[15]}
   );
   gpc1_1 gpc2991 (
      {stage3_31[36]},
      {stage4_31[16]}
   );
   gpc1_1 gpc2992 (
      {stage3_35[6]},
      {stage4_35[5]}
   );
   gpc1_1 gpc2993 (
      {stage3_35[7]},
      {stage4_35[6]}
   );
   gpc1_1 gpc2994 (
      {stage3_35[8]},
      {stage4_35[7]}
   );
   gpc1_1 gpc2995 (
      {stage3_35[9]},
      {stage4_35[8]}
   );
   gpc1_1 gpc2996 (
      {stage3_35[10]},
      {stage4_35[9]}
   );
   gpc1_1 gpc2997 (
      {stage3_35[11]},
      {stage4_35[10]}
   );
   gpc1_1 gpc2998 (
      {stage3_35[12]},
      {stage4_35[11]}
   );
   gpc1_1 gpc2999 (
      {stage3_36[0]},
      {stage4_36[3]}
   );
   gpc1_1 gpc3000 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc3001 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc606_5 gpc3002 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc3003 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc3004 (
      {stage4_1[6], stage4_1[7], stage4_1[8], stage4_1[9], stage4_1[10], stage4_1[11]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2],stage5_1[2]}
   );
   gpc606_5 gpc3005 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc3006 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc3007 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[2],stage5_7[2],stage5_6[2],stage5_5[4]}
   );
   gpc606_5 gpc3008 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[3],stage5_7[3],stage5_6[3],stage5_5[5]}
   );
   gpc606_5 gpc3009 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[2],stage5_8[4]}
   );
   gpc615_5 gpc3010 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1]}
   );
   gpc606_5 gpc3011 (
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc606_5 gpc3012 (
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2],stage5_12[3]}
   );
   gpc606_5 gpc3013 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[2],stage5_14[3],stage5_13[3]}
   );
   gpc606_5 gpc3014 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[2],stage5_15[3],stage5_14[4],stage5_13[4]}
   );
   gpc615_5 gpc3015 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[12]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[2],stage5_16[3],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc3016 (
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[0],stage5_18[1],stage5_17[3],stage5_16[4]}
   );
   gpc606_5 gpc3017 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6], stage4_18[7]},
      {stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[4],stage5_16[5]}
   );
   gpc606_5 gpc3018 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[5]}
   );
   gpc615_5 gpc3019 (
      {stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc615_5 gpc3020 (
      {stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage4_20[6]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[4]}
   );
   gpc623_5 gpc3021 (
      {stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[6], stage4_21[7]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[1],stage5_22[2],stage5_21[3],stage5_20[4]}
   );
   gpc623_5 gpc3022 (
      {stage4_20[10], stage4_20[11], stage4_20[12]},
      {stage4_21[8], stage4_21[9]},
      {stage4_22[6], stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage5_24[1],stage5_23[2],stage5_22[3],stage5_21[4],stage5_20[5]}
   );
   gpc623_5 gpc3023 (
      {stage4_20[13], stage4_20[14], stage4_20[15]},
      {stage4_21[10], stage4_21[11]},
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage5_24[2],stage5_23[3],stage5_22[4],stage5_21[5],stage5_20[6]}
   );
   gpc615_5 gpc3024 (
      {stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[3],stage5_23[4],stage5_22[5]}
   );
   gpc615_5 gpc3025 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[6]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[1],stage5_25[1],stage5_24[4],stage5_23[5]}
   );
   gpc615_5 gpc3026 (
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10]},
      {stage4_24[7]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[2],stage5_25[2],stage5_24[5],stage5_23[6]}
   );
   gpc606_5 gpc3027 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[3]}
   );
   gpc615_5 gpc3028 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[4]}
   );
   gpc615_5 gpc3029 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[5]}
   );
   gpc615_5 gpc3030 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[18]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[3],stage5_29[3],stage5_28[3],stage5_27[5]}
   );
   gpc615_5 gpc3031 (
      {stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage4_28[19]},
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11]},
      {stage5_31[1],stage5_30[4],stage5_29[4],stage5_28[4],stage5_27[6]}
   );
   gpc615_5 gpc3032 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {1'b0},
      {stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage5_31[2],stage5_30[5],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc606_5 gpc3033 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22], stage4_29[23]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[3],stage5_30[6],stage5_29[6]}
   );
   gpc1163_5 gpc3034 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage4_32[0]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[4],stage5_30[7]}
   );
   gpc1163_5 gpc3035 (
      {stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], 1'b0},
      {stage4_32[1]},
      {stage4_33[1]},
      {stage5_34[1],stage5_33[2],stage5_32[2],stage5_31[5],stage5_30[8]}
   );
   gpc606_5 gpc3036 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[3],stage5_32[3]}
   );
   gpc606_5 gpc3037 (
      {stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5], stage4_33[6], stage4_33[7]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[4]}
   );
   gpc1_1 gpc3038 (
      {stage4_1[12]},
      {stage5_1[3]}
   );
   gpc1_1 gpc3039 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc3040 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc3041 (
      {stage4_4[12]},
      {stage5_4[5]}
   );
   gpc1_1 gpc3042 (
      {stage4_4[13]},
      {stage5_4[6]}
   );
   gpc1_1 gpc3043 (
      {stage4_4[14]},
      {stage5_4[7]}
   );
   gpc1_1 gpc3044 (
      {stage4_4[15]},
      {stage5_4[8]}
   );
   gpc1_1 gpc3045 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc3046 (
      {stage4_6[13]},
      {stage5_6[5]}
   );
   gpc1_1 gpc3047 (
      {stage4_6[14]},
      {stage5_6[6]}
   );
   gpc1_1 gpc3048 (
      {stage4_7[12]},
      {stage5_7[4]}
   );
   gpc1_1 gpc3049 (
      {stage4_7[13]},
      {stage5_7[5]}
   );
   gpc1_1 gpc3050 (
      {stage4_7[14]},
      {stage5_7[6]}
   );
   gpc1_1 gpc3051 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc3052 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc3053 (
      {stage4_9[0]},
      {stage5_9[3]}
   );
   gpc1_1 gpc3054 (
      {stage4_9[1]},
      {stage5_9[4]}
   );
   gpc1_1 gpc3055 (
      {stage4_9[2]},
      {stage5_9[5]}
   );
   gpc1_1 gpc3056 (
      {stage4_9[3]},
      {stage5_9[6]}
   );
   gpc1_1 gpc3057 (
      {stage4_9[4]},
      {stage5_9[7]}
   );
   gpc1_1 gpc3058 (
      {stage4_9[5]},
      {stage5_9[8]}
   );
   gpc1_1 gpc3059 (
      {stage4_9[6]},
      {stage5_9[9]}
   );
   gpc1_1 gpc3060 (
      {stage4_9[7]},
      {stage5_9[10]}
   );
   gpc1_1 gpc3061 (
      {stage4_9[8]},
      {stage5_9[11]}
   );
   gpc1_1 gpc3062 (
      {stage4_9[9]},
      {stage5_9[12]}
   );
   gpc1_1 gpc3063 (
      {stage4_10[11]},
      {stage5_10[2]}
   );
   gpc1_1 gpc3064 (
      {stage4_10[12]},
      {stage5_10[3]}
   );
   gpc1_1 gpc3065 (
      {stage4_10[13]},
      {stage5_10[4]}
   );
   gpc1_1 gpc3066 (
      {stage4_10[14]},
      {stage5_10[5]}
   );
   gpc1_1 gpc3067 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc3068 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc3069 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc3070 (
      {stage4_11[10]},
      {stage5_11[6]}
   );
   gpc1_1 gpc3071 (
      {stage4_13[18]},
      {stage5_13[5]}
   );
   gpc1_1 gpc3072 (
      {stage4_13[19]},
      {stage5_13[6]}
   );
   gpc1_1 gpc3073 (
      {stage4_13[20]},
      {stage5_13[7]}
   );
   gpc1_1 gpc3074 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc3075 (
      {stage4_15[13]},
      {stage5_15[5]}
   );
   gpc1_1 gpc3076 (
      {stage4_15[14]},
      {stage5_15[6]}
   );
   gpc1_1 gpc3077 (
      {stage4_15[15]},
      {stage5_15[7]}
   );
   gpc1_1 gpc3078 (
      {stage4_15[16]},
      {stage5_15[8]}
   );
   gpc1_1 gpc3079 (
      {stage4_17[6]},
      {stage5_17[6]}
   );
   gpc1_1 gpc3080 (
      {stage4_17[7]},
      {stage5_17[7]}
   );
   gpc1_1 gpc3081 (
      {stage4_18[13]},
      {stage5_18[5]}
   );
   gpc1_1 gpc3082 (
      {stage4_19[12]},
      {stage5_19[5]}
   );
   gpc1_1 gpc3083 (
      {stage4_19[13]},
      {stage5_19[6]}
   );
   gpc1_1 gpc3084 (
      {stage4_20[16]},
      {stage5_20[7]}
   );
   gpc1_1 gpc3085 (
      {stage4_20[17]},
      {stage5_20[8]}
   );
   gpc1_1 gpc3086 (
      {stage4_20[18]},
      {stage5_20[9]}
   );
   gpc1_1 gpc3087 (
      {stage4_22[23]},
      {stage5_22[6]}
   );
   gpc1_1 gpc3088 (
      {stage4_22[24]},
      {stage5_22[7]}
   );
   gpc1_1 gpc3089 (
      {stage4_30[6]},
      {stage5_30[9]}
   );
   gpc1_1 gpc3090 (
      {stage4_30[7]},
      {stage5_30[10]}
   );
   gpc1_1 gpc3091 (
      {stage4_30[8]},
      {stage5_30[11]}
   );
   gpc1_1 gpc3092 (
      {stage4_30[9]},
      {stage5_30[12]}
   );
   gpc1_1 gpc3093 (
      {stage4_32[8]},
      {stage5_32[4]}
   );
   gpc1_1 gpc3094 (
      {stage4_32[9]},
      {stage5_32[5]}
   );
   gpc1_1 gpc3095 (
      {stage4_33[8]},
      {stage5_33[5]}
   );
   gpc1_1 gpc3096 (
      {stage4_35[6]},
      {stage5_35[2]}
   );
   gpc1_1 gpc3097 (
      {stage4_35[7]},
      {stage5_35[3]}
   );
   gpc1_1 gpc3098 (
      {stage4_35[8]},
      {stage5_35[4]}
   );
   gpc1_1 gpc3099 (
      {stage4_35[9]},
      {stage5_35[5]}
   );
   gpc1_1 gpc3100 (
      {stage4_35[10]},
      {stage5_35[6]}
   );
   gpc1_1 gpc3101 (
      {stage4_35[11]},
      {stage5_35[7]}
   );
   gpc1_1 gpc3102 (
      {stage4_36[0]},
      {stage5_36[2]}
   );
   gpc1_1 gpc3103 (
      {stage4_36[1]},
      {stage5_36[3]}
   );
   gpc1_1 gpc3104 (
      {stage4_36[2]},
      {stage5_36[4]}
   );
   gpc1_1 gpc3105 (
      {stage4_36[3]},
      {stage5_36[5]}
   );
   gpc1_1 gpc3106 (
      {stage4_36[4]},
      {stage5_36[6]}
   );
   gpc1_1 gpc3107 (
      {stage4_36[5]},
      {stage5_36[7]}
   );
   gpc1_1 gpc3108 (
      {stage4_37[0]},
      {stage5_37[1]}
   );
   gpc1343_5 gpc3109 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc606_5 gpc3110 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc3111 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1],stage6_5[2]}
   );
   gpc1163_5 gpc3112 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2]}
   );
   gpc1163_5 gpc3113 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[1]},
      {stage5_11[1]},
      {stage6_12[1],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc615_5 gpc3114 (
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[2]}
   );
   gpc1343_5 gpc3115 (
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1]}
   );
   gpc1343_5 gpc3116 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[2]}
   );
   gpc606_5 gpc3117 (
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[2]}
   );
   gpc615_5 gpc3118 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[3]}
   );
   gpc606_5 gpc3119 (
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage6_25[0],stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[2]}
   );
   gpc615_5 gpc3120 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[6]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[1],stage6_24[1],stage6_23[1],stage6_22[2]}
   );
   gpc1163_5 gpc3121 (
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage5_27[0]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1],stage6_25[2]}
   );
   gpc117_4 gpc3122 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc3123 (
      {stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], 1'b0, 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[2],stage6_28[2]}
   );
   gpc606_5 gpc3124 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[2],stage6_29[3]}
   );
   gpc615_5 gpc3125 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {1'b0},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[2],stage6_31[2],stage6_30[3]}
   );
   gpc606_5 gpc3126 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc3127 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {stage5_35[6]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[2]}
   );
   gpc1_1 gpc3128 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc3129 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc3130 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc3131 (
      {stage5_4[7]},
      {stage6_4[2]}
   );
   gpc1_1 gpc3132 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc3133 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc3134 (
      {stage5_7[6]},
      {stage6_7[2]}
   );
   gpc1_1 gpc3135 (
      {stage5_8[6]},
      {stage6_8[4]}
   );
   gpc1_1 gpc3136 (
      {stage5_9[12]},
      {stage6_9[3]}
   );
   gpc1_1 gpc3137 (
      {stage5_10[2]},
      {stage6_10[2]}
   );
   gpc1_1 gpc3138 (
      {stage5_10[3]},
      {stage6_10[3]}
   );
   gpc1_1 gpc3139 (
      {stage5_10[4]},
      {stage6_10[4]}
   );
   gpc1_1 gpc3140 (
      {stage5_10[5]},
      {stage6_10[5]}
   );
   gpc1_1 gpc3141 (
      {stage5_12[1]},
      {stage6_12[3]}
   );
   gpc1_1 gpc3142 (
      {stage5_12[2]},
      {stage6_12[4]}
   );
   gpc1_1 gpc3143 (
      {stage5_12[3]},
      {stage6_12[5]}
   );
   gpc1_1 gpc3144 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc3145 (
      {stage5_13[7]},
      {stage6_13[2]}
   );
   gpc1_1 gpc3146 (
      {stage5_14[6]},
      {stage6_14[3]}
   );
   gpc1_1 gpc3147 (
      {stage5_15[8]},
      {stage6_15[3]}
   );
   gpc1_1 gpc3148 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc3149 (
      {stage5_20[6]},
      {stage6_20[2]}
   );
   gpc1_1 gpc3150 (
      {stage5_20[7]},
      {stage6_20[3]}
   );
   gpc1_1 gpc3151 (
      {stage5_20[8]},
      {stage6_20[4]}
   );
   gpc1_1 gpc3152 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc3153 (
      {stage5_22[5]},
      {stage6_22[3]}
   );
   gpc1_1 gpc3154 (
      {stage5_22[6]},
      {stage6_22[4]}
   );
   gpc1_1 gpc3155 (
      {stage5_22[7]},
      {stage6_22[5]}
   );
   gpc1_1 gpc3156 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc3157 (
      {stage5_30[12]},
      {stage6_30[5]}
   );
   gpc1_1 gpc3158 (
      {stage5_35[7]},
      {stage6_35[2]}
   );
   gpc1_1 gpc3159 (
      {stage5_36[6]},
      {stage6_36[2]}
   );
   gpc1_1 gpc3160 (
      {stage5_36[7]},
      {stage6_36[3]}
   );
   gpc1_1 gpc3161 (
      {stage5_37[0]},
      {stage6_37[2]}
   );
   gpc1_1 gpc3162 (
      {stage5_37[1]},
      {stage6_37[3]}
   );
   gpc223_4 gpc3163 (
      {stage6_4[0], stage6_4[1], stage6_4[2]},
      {stage6_5[0], stage6_5[1]},
      {stage6_6[0], stage6_6[1]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc23_3 gpc3164 (
      {stage6_7[0], stage6_7[1], stage6_7[2]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc3165 (
      {stage6_8[2], stage6_8[3], stage6_8[4]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[1]}
   );
   gpc623_5 gpc3166 (
      {stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[1]}
   );
   gpc1343_5 gpc3167 (
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc3_2 gpc3168 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage7_18[0],stage7_17[1]}
   );
   gpc1415_5 gpc3169 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4]},
      {stage6_19[0]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc623_5 gpc3170 (
      {stage6_20[4], stage6_20[5], 1'b0},
      {stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1]}
   );
   gpc1343_5 gpc3171 (
      {stage6_23[0], stage6_23[1], 1'b0},
      {stage6_24[0], stage6_24[1], 1'b0, 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2]},
      {stage6_26[0]},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[1],stage7_23[1]}
   );
   gpc223_4 gpc3172 (
      {stage6_27[0], stage6_27[1], 1'b0},
      {stage6_28[0], stage6_28[1]},
      {stage6_29[0], stage6_29[1]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[1]}
   );
   gpc623_5 gpc3173 (
      {stage6_28[2], 1'b0, 1'b0},
      {stage6_29[2], stage6_29[3]},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[1],stage7_29[1],stage7_28[1]}
   );
   gpc1163_5 gpc3174 (
      {stage6_31[0], stage6_31[1], stage6_31[2]},
      {stage6_32[0], stage6_32[1], stage6_32[2], 1'b0, 1'b0, 1'b0},
      {stage6_33[0]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc1343_5 gpc3175 (
      {stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[1], stage6_34[2], 1'b0, 1'b0},
      {stage6_35[0], stage6_35[1], stage6_35[2]},
      {stage6_36[0]},
      {stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1],stage7_33[1]}
   );
   gpc1163_5 gpc3176 (
      {stage6_36[1], stage6_36[2], stage6_36[3]},
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], 1'b0, 1'b0},
      {stage6_38[0]},
      {1'b0},
      {stage7_39[0],stage7_38[0],stage7_37[1],stage7_36[1]}
   );
   gpc1_1 gpc3177 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc3178 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc3179 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc3180 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc3181 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc3182 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc3183 (
      {stage6_4[3]},
      {stage7_4[1]}
   );
   gpc1_1 gpc3184 (
      {stage6_5[2]},
      {stage7_5[1]}
   );
   gpc1_1 gpc3185 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc3186 (
      {stage6_15[3]},
      {stage7_15[1]}
   );
   gpc1_1 gpc3187 (
      {stage6_16[1]},
      {stage7_16[1]}
   );
   gpc1_1 gpc3188 (
      {stage6_19[1]},
      {stage7_19[1]}
   );
   gpc1_1 gpc3189 (
      {stage6_26[1]},
      {stage7_26[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor_CLA256_32 compressor_CLA256_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8a39080463ab377ddd1e36a9beeee63bf6819ed7cf061b6838f7ddd7a66ddda2a2599056de7d528a8490f3b91b60b951d3b9e5bf2204b582b0ca7073a30b4098943a04b137110dc1fb4f067aacff65e83034bd1662d0ce688927215744e970f9e47a5d3d6f31841a40225935c807d4753c056c41edf5cd8ac323e3078c913b903b6472c85c23575136dbe1052c3a3092a6d6bca3f219702d231f4501ba1333b78f966c3a5afd0528de752fe3202437e6830e2f843c9a3b7e4b4604f04bd24ece3ce40a200c9ae6091e5193004df85083e173d736b0bbabd18189f51c8b7b757fbea6126ab21bea481fefb6b0a261b5cf22c4dde5ec700ab8e302a758955780f0a1ce18776546812ff415b6a6775d1e80b2dfc53bce91bddf8f2009980a8c1d457f0719f1506f4ed2f0a92ae974ba4aaa060b1a2cabfc3a6ba176f4f1b0a93c46d583d309f7ad294632468560e19a6e9dccfaffccd54e0ec4e2c2cbee778569e565068c80ee009cbf2f116fadd94c0386f4da5ccb932f9d502f21cf01e7a737a85d0e80fbb91935b3a7ce39f5215bd78f396dc8a739f924ea73f2ecc42f9cb2086027ac94b502a8701e6887f4346e96cae7210ac9e75e21891d8e82841b0004b1854c6d34aaf4aa3bbe25f316b7a889d253ab15b0dae47a59666a9c1584c59a5db5b193cf72eed41384199f9329d4b4fc47b8625032fee2b5cfcb91eb406e3f251dd34f924eed90625eb431e1c1d8815dfa7ff3b1bde812c148c1705d2556f687e5b55403195a06f5188367e215a49c65325e5b0a1ca453bef59469239f9d4417753c141ccaea8413e6d42cce9f7d51efdce97a7cf794e264efdb639a3c42de50d477b24664a75be13bc16cc729a1df4b9ea3a02b0910811ee73cb3dad0282f68c56e4b0a459534481c16c17c5f99c92f3bc5522a2afdc18a28428b23b3868833cbe3a03797c8c3fc883caa9f92ec534f0a38fecb0846fe2da14587d362ecbc026096db0547308f9dd8d5057d523ecb93a8cd430d65a46550ea89f7f984e54765f8eb0e18de71b1bcbca6e64e8e30b7ab43415ce9078dab6677d546e9bb8d1353173fc8ce2581af41990460b83f0c310a99b34f2158bff46801255c18c8c6e45f8b0adb45c3717c2a6c57474e3089662968835aff6b70d512b7761e40da756916c5e5509aa8daae8b8e7196b8a3b93c4e5af9197660f78755dc10c8a01bd73c29720e403c6670ac5d2114c72eb589e846592512949329f40b5862c1b2de168dfcca92a804bb31b18b391450e4b63efb38440bc33bf92e243fe322c47a7098256f5c549d84e07b143d6cdf33e3965e2c9777257956188d745a12a0e57c17ea4448fe182dfefec64198c3a0bca8fa177e9ee9e0f77851f0ad04b3df063639debcc92e9b19aeab80ee63cb2636630a245413ad87fb4b257b7942354123ac59da1eca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h85ec8cf3a54da0f44bd4e2477a302da447174131c9bd80b655885957ec974609be5f86ff7b557baa82104737ab5cdc421b82d9f3ff0a11400e5ea01b73169efccedcd44d46a1a1d723dd5e20bbf8291e9958b5b0544ba631f37b6500a70049fa1a1ab34ee241024a1c0307e58d63163baa3972e6448d8b5970653d7cf7371be63baeb7788ebc1c424068415fb6759b04bc12f940e9488ef3facb7b43a6ff2b87a7352729fe4f3a94358593f25429bfccc41a554608d7e85e84e74b5bd581f075e30c244bc5d96d0005d7e2c33c1a54cfbb6708aa284c631415b41e81c031a8ac29165792034fa9b78cbbadfdc5d7f3d9afb10e4b5c4635efc93d49c44e8e820ef88033fc76aeff51017b5dc1d809fa62966cbe7d3450b67cdd4a87222f364aa23eed79ec2e7707158a15a568f21317fb16d0184440740fe0b99f5fd2b51220c116f167f87863ecb9951a9124d86726284c489bb47ec281e68042908a12517e333a63400d502cf55eb3647990075d9f0bf11d3d479b5739cf6cdf737a29b1d4068bb762948aa6bdbf8879973b963f07627ed99961bea6ba6fb507816f9cd42d1221c96e3a46f39ba771da6cbb8afcd91bf4fb2a1deee277a56838af9340cae1119985d1b07e3c2eb2ecf2795137479e152cce97aa8492567ed82b2b020db8f154a87ececf613597deaa097134db03ccb56693f6b0c12fa4727d5804517a0de485774c0e040b908778a5e27f6dfec19bb933fe0d84bf1da2f4766283d7580078ac2aec0206b0f9cc73741b171ef92327a0000d00175c26d6a9cfcef134457d804ba84424c05cb4f1c4b997427e530c70d84208825d2d82b70e778e4e2be4116e13f5e82160fa244373c1ab7921a982cba7e6420ac5c88d9ba75a333a5953e80fe317f71066069860c9164a6332aa5c4949ee73021599a9b5ad007a8e6ef0152c215a86670d508e2d5508b8c374eb209384921a1a6f9de4ecbab9576e5e6c35955a255217afd7488ed366f56f421ee45c9e653740fcf36ad6e5b49699cd8bd302f735cd7a13176eda80be939b5936a96276ae4b41129b747e661d5e91a7b7a34d8034e3514e003149179df8b52edee55873378ac165a2c352361071a5bf96b18f0e8e69e39a7e7c7f08c1f7f785b49f826fecf36270d84eeb84aa730b6e58a75f69803e5d4fe84ec0f0c7bcff90010b8abffc6416406d28b3a668218ef0e83876b428b39321fa2f83542eccabdbc7e7032c01a3dc3a4997a9a547b9702d774e3aea32ff5ba2bc85480ae09a8c8975d717baed57f4189553083a1834677b5439b56dd366d249fd187d17cfd89e7cb68b0ee7e5f818a919584038e3f570d45b0f034b23998be9b9c17c1d54b87f84fa80074beb47b8913b94b12af4ca0eff67012ea0194c09cd1bb374b9ab7be4d53fce6c42b7b89bda6fd4488bfdc5a1d97c8dc7ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf6b7e09813c6c152e90b12f74c027259a895be5801b02a2a12f99817bae7454d436ad568a671eaaac33e818c800616715346865783af34af4105fa38d165998520cf320e6944d9a0829d23531edc1be0bc812727ea4208941fea72b1673d81d3fc913d10fb3816cf5513013d99215c0b18943ed7497a895e2c9684688babdca71431e7e58c5c5b6afbb56b845076776eb0573c1f3146af59d129c59b820596925172b39147d555711fd8c9e83b1abb3c67d5075ff992a24c1d56332c78bf7a1fc565600c245cc4cdad0711523598996bb0b31cb00244d0e150a7efbab29f5bb435be8ba8e970bf93d4d513115215b1cb1107d1ce00a57cd814c53ebf1df5c47a927f281b3631864eb5363a5503b1b546b4af76a29cd3f354123b76fb13c2bfee2d2ffe4b089f1ee818d5bf550bb1739ed400974a2230149159dca16e21bfce5de957d2309f940509e748f09a33675526c27cdbaa66d10831ca28a764c972f1293deb455c4eb365b8885e99c5e8e1d5a17a7f8e328935cf709e6a33ebdbe247748fb3d6d94130e91e728858b174b73d8642b91fab587ce3c507f0907f5b3c77806ebf5bc7fbd86dea3230942b113558ba65911fb7e365a5ac09d06b52477fd418db2e5fc750b5a9488744ab4d3b880c1fa7e25dc9744c5a2ef2f59d1dc991e8d05836bbbca2955a1800e0ae2c89b70fa6a47cef155445ee84883bc4537d96b3383b660d3534f25bc29d254739dd5606fd4b5c836982cf82d563ad37b742ada0b051a6656aa4a1acec2d5013c8b0cf570ee7483edf25f7056de9162a3f62de5a6a8d75f1dadbe1faf46d0d60f036dfaca27a63dc3759a240342ced1d6bd6f245cf027ab1504f4865cca5b632d3227d25d8b514499b9cd724facb1d08e4d81f779615bf64bec347067f2d7d22f2f74ecde5a7e27132eb14fdde7f77688aa84629b73e928dea3d68082d97fff2b82380b7380380cfc2ea4fcf3f223b500aac6d648efccf093df0ea070020006834d09c1592e77271fca919ff595a273f6c89ca3713992d3416e94b7181637ff27f396901af9b557485eac5c4a82011be476ff2bf287dca9a5571add417ec0024f9d026a942fd92b8931944c8a7b07dc6bc88585d495789db07e543020b5f43205c7e3ae071045aa82774f8db2e2ad200d83c14d3e70539782c6a11abd19ea53431f710d336caf8e2974e066386d96f5940d57027ce048d8eb2455dbd4a61d2f192730098883082d74029d213485336fe4f78d336f0839d49fbe4ead652d852ff6b47451ef2a3bef1afe809309a8c8a40a26d9b81c5df2961a8ea8b5e027d873e0b56eed6de4e9d52d5df91c77841e5713b4b2a66835c8dacbae181818aa909334864e77c0971b647a20a8efab95004e9b2db9eeca759c3d3a065490a0e9bb57d3c151100ed468b7b21555a56801895e8541d97ef10;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc7eb3d1339e2103f72ad3502a29e0b397fad3019fddc7fed3899fad0ae04f5f0db44ccd89c251523571f5b2646865a008db9caacbd81681a46c5a06f3a75c614b2f42cbc87f512c9c998849d4a5fec83d4fcbf91cae87bd2951bb814494827138505a62f8d47725325f8349305909830754e7d141740ffef3694246496cd651ade0fc2af4ea3d71b8391ec5adbbc0f81beb3d831b9ead743883f2439d838a997ef83185d69fea0a2ef9cb2636f15050c5f71bfd80b727b6514d71e2baef084a71cc0b1069af56c899dfc93fdbfca06b2d370dda9b4b8ae6299d2602fe6abcd2fa58ea539c2b211d7e19781853607121ede892c9df28bf6c2bf1d1dc1ad6c815bc91d520fc815d1b38c3ac1ef6d09abf7fd2026109d9de282c0dc06e02d6f7a0e521d570fcb5e30107eecb1d0bafb846f4798ebbb7473be123a169d3e9644a84273c3067e32abefdfb8f2b69497e2463362f9236018d0f946d531a1a74ff124f9a0c8479c8af2caaac10d181d7f3e56778c11f84845824d9b150d5b2a2ed37dd06bc626e2767c444c9ef95dde16c96a3bb4ce3af7eb73db3dcdbacb19ff2c96a1fe52eb825e2245cf267aa10950d2a5efe993d31b5c664c56b1969d633c2c0207311968eeb6cb946c434f843a5923c90394b5bedf26f6995f4aebcc3b2b243f72343c79ea11a686cbee8496b47f02a5b5427dc4cf6ccb89b2c8f8f2a06d36727dcde298953cd87680651129cc905ea4c3961124713d0a73d85902c754294c5d26662e5a42b066ed017219d9e57023367b6a132a812eb7dce601eac1a7834ccbac646432f33eef3f5ba8207e4620eb31d0a830218e2b758ad1b14fa142513916067dfcfe5ef25ed82744b0536fc607f9f4f66121740cf9b3c63180569e4e1a514e59cc6c238136c2ea7de8ddd6832e2fe7e3b6a4274671e568c6fa9cf51a5475ecc9a74931d11d258098786ba0aa443cb0cdde1da174e7f5bf873d04b2139442d713b257d06b0d2f0d084f62bc0deaa82a8890c4b8348982e94319cb683167f658f11ba53ce9a67d67ead57193bfe993e43179f2ad105d43d9dde09a90441317fb33c106ddf612bf538ded52b8796f047e8b0b49a93e7d4f77ab4829bf20d2578cd244260a8d098ab8edea808260a70862b85d4acf055f909b03588854e4aca247944f40e2149e996d1647c9a46e4b66fd8e7343890d1c1af0e3f514153d56cb135e14942df5d403c752684325341b8f50658fc59f9727e1994f7b350d137ae4a5022a826f62abf9147459ecab4c8ac9cc76f31c75f82807f20b488ee49631aae9802c78e788ab6e3efbe5aa84a8d1bf102a2d236c4cbf2853073d0c06b5fa92fccde2b459bceb5e9e8c148c4f6c482806b69da79912729bada0035f76d8be4e065c945007f34353c62a6b43a6bcfd0208561aef2a43db334d57c185baee1b9aa7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1edab326f50d3656d8152b8ef6bacd4b7acfb4e34a20a4ed00c856ececdd357a492779c89bbcb4b724c782a44df7e3b939cf090016965b1a5980b36e6fd19d02ad14a8842f1a7d3c1b017eaa931b6c4aaffe8b840058f873281516ad4b83e19d9f9807d64856554ccdd7ce0ebc6ddc99339f4a6950fcfad4489c1b59fd5f43d672d0b71558d1211768e0d4add2a849fa915237a44a6be8bb3d9e40a488522de0e25b485975631c98a00cc538596d784654ab4f321b51ae02eb0e08e82185e9f3558da6f6e58372a5594778772583a4a0bc490097b6d5c56289c005cc3ac3961e9c81c8c95fee40c4029408b1c1e89ae2127d5325f4d3e7feffd1e13486861f4a8c377c650f0ab7ee9cba3239e1d38e834c84440a502db6883ce8711d59dd80ba32eadf380a3a04bc2504d3b573660c47dd8cdd543d52a8566f537758e4d41b601b2fbc4cd7252221a614a79a7eacb7b484ac4b07901a5676e2678aa600be3f6f4fe525ab3263ee9602758484aec3caabc3f53edfa9747a9b6c488c2ccb113ce388e57299e2eb94396f68547316ccf12e2f7645a96c9e52f72cdb03476d0a59d178b97ccf4115bc90695ccdc33cacfae4ff108a782ff15e15476b59702dc708fdda9cef91f6b30ba6e5b47298da9eed1283fe9ba0f1a8c7594baf475d1d0806bde53fb05d294cc7629389ef76704ef359527705edb6d893e7ad100fa5aa6e8f7106ab73cda9f4709cfe44f77804a4ac0dc9206e4a7175ac7b5f2ae80df795c6ccc25c35c428195c8d6671588a0e0bce2586a099492757283888b98c1224ebd02c5107d4c381473462ced1613c7f782a3b1d903a6899c99edace9a139a85bef259fc3dd22909d0752d7fbec0e51d84b73ee27d74b5b0d98a79e096ecd108f4d0c8dd3e0c8e7029ab1f7ba72fdafaaafa254820cc61b3f64b3e162a2da185a29b8094ecd02be4fea21d53d628d6e463d2ce03e83e8acc85a4fa30ccbeeb4c86c1b09db9125db15c11492313eab424a9e7ba2cc94b635fdb8641b5c995b15bf7f808c0080863c6347ea1cf2f04d6f39dd44af821da8446e4b0322ddf6fe77c7119580975e2d1ba30391c271f38bce0039e77e64eba9c31e7ccbbb289cba1dd3d8e651017e642aabebc847e3f45af45e51dafc1debb68e698f226b2be79731f67fa41a5f692c1233c8f603be3c028a54fa70e456eb91bf26b5e2f035172a1a20f44f47127b655d1eb8dd035e762fb0790ca1405d322776c0d6ef18cc2b3ab2fcc615b5724c3bb327a4405fe71a16d2fc8d9d15ebe61a97eec645a9e2177a236ae0009f00a3f6042295a6a75a8057f5504301e09d628fd87086a0da7fd16ea66b8aac30dc90fc7d22682eb4500217a3f293481443d74d2a27d339b6411297e6a62ac1c1bd652a8ae0e47ff0e70d5beb18911a82210583adc62e3e795e95bf0a34108f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcdab951f4d3cf574fdd3e9aea2b2b1524bd709c79e09b74cf840b168d508e91af02f9b80597700124f55065ae0b75c83c8ceba88a7bfc0aa20cc7dca0252b5cdd2c6e682718b694b79ec22bde6ca4c9828ccaf1e208fec6e9c5097e32dd12885dd2ecc5abb392bebb601a815fc4f081fca18ed2ae92e7c2ba31535acb40a4a1c8b39716935451d53e6994ec0a5f727245807e0afe39c0d0d413f4af2fadec9ae9bc3b92a9f79a09b1a5390c30148463dbb2bd59caf56698b16b85f15668e0d6618619a0e01b4581e7dc47b276aa8cbe767577deea0769336051bbaa9e657002938e2343997752573d8b9355c7f2ecdc59973f6013993ecf336ea854b4056d094f0c7f22ec9bc75888dcc1f1ab02fb2b446f660506e1b78ac1500742780b9a2e9be9d80f01ea2ede278254c1875a5f0cb6b044aed72bc112ed41e5d1d6861b2642f00b78153fe428243a5a1d307b190246c046816f3da993048328cfe6ea181e2c582a100e95de839ca25f3a6e70a3bcc8b03547dea7af0c0882310ccc3080282b28c8052ddba30116f668d0d9321bdba81d2d5bfa8cea2ed999be7dac78ea29b2d7245fabb31456ff44171cd1adf5d282158824a8602b08349c77c5d2865ce8f763365bb676ae325cef5156c4d8e3921c660cbb17d1040d3636b7a7fda25d16a0e57e7703c00a58027deb92726414c20471df0ba6cdee26e123302f77d01abb9d22f6ed590e7d349e2c69ccd7cdf7d374c07caa234fd9dc00a07e9a3e3ab89e96d4c3a56de78246a08cda3dbb2e31240511daee69e65cd8b042af62e573d7793552256e99081f27922d4de73ef6c8b550653d7f819a4f8ce3082c96102565c017761f47b4f4a2d725d09c026a59b8a843a61242067bcc557b85ba159aa737745103ea4250cf2353ab884bb5fc44ff792ec45a1c100b413f506b82d4e03b7b8c4bd6acb8f5f3417216c95e9a1ad7116f672f43e9bd665d8cfce859016de9dae7590ed564aaa6712fca6602272ccb745e3839ae9eebc0028014778fb45c02f0a2b0bc2803603187454e8f5dabf02388c41d33937d5ba3f7f3856ad4ce562e75c98b3a86f45385e59c55017ec10d035edd6dd9dc2a6945558d94eb95f7701942548eca56f0dd0ea7e9d39fa5c4ed091a9fff5dadd0dabe03e07164d7ffb783fa0368d496a255c528ef5374f648cb0403de400d2cafcb9bd75fbfa174968442339388e552c454bdbdd22db268376b3e2957c02f0deac1f4a4b78753d797349b4e1c4487f62c175049078709ca0e432c423ea3a16f1bd3a594a838981f48308f265288bb1b55fea3b2a93e1045560ae84fcdbed90c22b24ab4ab8bd9068f8ad521f773ac2d43fdcfa22bdd6cfab8b203b337dc4b201ca4976834aa6b0503071503d6bf3a0b5a8ddeaf2e75ef4e9f68d4dc28fe70d116c8baaf185e5e87fd2ca001ce9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc1531486c1fbaabaa7af8e9691e3512d8a22ae2bdd4c91add69673805f810c9478e5fb958e88387c7391121d3d4231fcbdc95c28c447cde95354abce50c6a7d7edd3a4b34c68c5874b3f50522c449bf07960b0d8ca13b216d32cb9eb3d315d8a239713f425a0d51c686dc787e1d885b249f6784a9d632688c7af5d3d560ce0ec857837da884bfb728ff2ebae8360150819211a0ba06ebafb865134cbe8e3c64ad09a95698e6a23fa7f3c3d4e1c3ab0330d9bf12cb4b31378b6d4810aa3fe6442b9119761d7221958b94584ecb302c01b4117f559f193d550b06c7ca1d2bd4aaa6b81ed3044d06de09b1dee7fe79deaa3d1e04cbdface5151450a842a7ed0c89b5e262c4a8392c88bfa3034a1785a5189b79f8779c5b55ea5f9ba9dfb444c9d108feb44e13366da678c2321828ab5f046ebf5cbbc82b6688b54f7ea58ce740e36a8c4d0c379e08bebfa4901647788966378af884ea5d846433f9902f73948faadfe75e1a9b654cca3b507f81ceb3348d6ad2bfe8e08c97e6d4a1ebb61226003d3a7fcab4d92b3eb46fc574af41d77d5a8a76335d96630eee9216e59c3e9e40a2cbcfe7008b2bdca989aabe86c30ef3c7df4f4f8c45d765b2d943279fe30ff1323ff533d347eaed80a5601f5e20cb5677cdcaa9235da891a6003cf54832a739c2df665939766fd1618e87e3a01046f8e4e7454d29b487bb1a53988ca9e67085cd6f9c89c5edbc8606861fd5d6c15de5bcbd360fac0692201b8218db186d3468a46af5a61c363bd4158c827df6ccb8f312a218679504794cabe0a9e544e99fc5411102f254c8a881e5cc89a90ec8586f493addc90f70d5e55145820e10c78cc570e38027ddd50b2fd7e44e6cd7646ab5c38c800c2f5eda1052fd757d12d4de3aa821f30212f3c5bf8f8690e536e52a242f3a171d3e36e334345d9d9e7702c6201ef162175b308f4ad0d34313530a89e5e87d9f3f85d425860d07503125012f082af6980258dd996508ca757e5cff6e1fb979b0b767facc8889cbb9a870dc9066f44196ec48469b8e3fdd8f16f15bd8c62bbc553eaf26ebd459af67097b9ab48e31ecc5aaf91c60be59b73b6b305880eed6b7f5d01f8f6b4817c2dd35354a8cac0d28603d6b6210061588ac075574c712574179238e461a44a6891c88f8a5107283f8c3ebf77d08efc81a1e9a0f1e7ec628727d7f6e70cab48c8e1697f8528aea786fb5a19c608b5d7a656644e447da6e787ed1478e128fc45746105f0d6e5fc4e59812d4f4e4cde4cc4bb5c2bd21d30aaa67b1831c39c6237239cf89f0dadedb1a1b189ae61e447c447ec44cc1277cfc59fe461dddd0d36a01db71d7dc7d24b648e11c85fdd798b3f901267f3a2a22c6d144405e5d6770f7b68fdffa0aaede1d3e5696d231077e889e327bd1cb5e97f4a75f529f5aa630b8626ee0b0d41f645ea6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1c4c5438f56914042448bf0f707d4a7be4107931942e1bff7a8d07f5e148b51e4038e87189af1de710416dffde532d2fb32a4b4f8364d6c06fd0594d814b70f81eca0e4e82944a9c973aacda18eb10c668154567106ebde065a223aa33d07d7d4efe927fac365cc8d3e031ac360760eb98bc062dfba03854c39e6257dddf3f04fa791d36df8db24186891523cbbba5a9dfd80f78daa30d783f2ed6652957ca80b688bbf1b50f1ebc9fc2c7da52e11e92198acd0e61db8f93670df2aeb4df7122aff909e639168f37aa9c40f5e419740aac0e856bb54d69fa860effdf6cd6257960d0151781cc4365c2f1e1e80001b29e95ab4eac2ae07d11c0f6190050a1db5e031692badf4c46156d40d561440a480566fa64162140ecada5d66a6729e600b045e011c03fe8f8fc48627d2a7e813e9f28fea54c228944b2ed6f34375f3012d60437b148d01021ac3ded0455cc286143f6f51d7b720dcc1dd3f8a5234eed7a7b38adb3d454e99457797b13a748d39d3fbb9c033d1eba255223798e5d3a68bff88231168debf6b5cda2f4f7c33ef3a3b96685fc9ce34c449895948131bef0c750afb2e2f1c804cfa63bfc58c93fd593e3ddc3d43953758c86bc641a9ed4164443c3115a90eed238717d10b36c6d794b1ff09e71338c84f0ecbd3f4c671f0ed6be740e50fe1ee1aec47241722eb9ec0e83ce48a440cc560f5ee1cfb0856aee297aab1f9d977131915aaef0735cb817d15957b0d9dbc77e029682823de3891eb33585480c0ddc681436ccf549cb6821882bbf7f21b2514aecd10c2a76048715b3e37ae4479e32f4fcf930c1002268690c814a970374ea659d85338d3cf0a10c21b53f5e8cf70e89d6cd179b0fe3c86c68e162d8fae55a7f6f96e2db3b74ff94103e4398b3e12f7110d97436884162d1366b3caa72a42d32a49be62d930dfa28b5f7335846964b53d50e5bdf0eb82ff445bad0729daf70bacebde7287f4c2c89f9ec320f4aa436c55d9504548cc34a5c03545be80356091e538fa696b7818c9f628fa5ee10befe9b8d38f7f953d30c76fb979e25ae1a8c95d42a66c50b8cfcfb3b6c74d18087b69091401e7c36dba4d0cb9020f5c92309fddbb20e41794d0f6824145346955bd0d73c1b1b646a1a28eee6aed029b36a3438b3f2b6a2f6837a7733b34f23169352f55ff69ea8efcb5ee830240056e5f7a6ebd818a27e87ed411498e4cfa7efec534a6e54b157da2443c1b7bb67ccc3cbca48f3de0ecb665ac60752aa8ed4ecdedfe0d527442965cbde738d83509d4de548e6b775f6142b21770ea9692b36365c50588333eb832ceceb3f4432e9537c57e807521daa0e2101134c3abbdbc5aef14324c2c0bcbe3f235ed33bb2a51616327d3fcfcc2024efeec5b59e66b8b084292b899149de3e255d55c092c31f95ea21ac913a4e1d0d131c0e67dd12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe47de131dc778c0ff6f455684f9acd5ed62f3f66b24f1f526378b8135b896165619f98644681e8c331e20845fd74cffc907b785e8667b558d6edb3cc64e50d84f3a2239b85df930f0c6087bb88968c07fe5c74e8c318b73f471b32f354f4104f5dfca250d559158c6706cbb4a76d25a0c5df927a8641c03e765ab5a00310eac494f3e5fae83c07c9f0f7e361ba1cb8c7ca9cd55457e8f1a3f8b06fc8e7f258753c4860b500038a3f55250f762f414b8cef4b271493a0b7cb2e4ac8cb5c2b2ac0b3ee0dba476df06097aaee2b64f80fbe37d47d0d815ff871116fa1864ee8e286e09a06b88c18ad74139475e3ba3e4ea994e33b1ea12fae5dbc25a2a7e7562d46ea1c3ea0e15ded1822c078c5a1b70fc374442c5db2e07ec69ffe51906b74242c46447a653af1d071698afe2a018bfa0867ec3ac2de14f6481d78e0ea007a5c19419405e2ce91d2e1060ff4deffa85b88eaf0fbdc6796aafd8b50246089563437e879abe8674ce9bdf071c8efe2c53ea60a1710e1381bdfa95839e01e81f2031cedf0e8e4f64bea317ad2866cfd03288743641a5ab41e041a6fe878df69ae481a2373c7228f737070a0f9df7734a9e1812c8bdcccbe425e95d555c38c85db71ccdbcb947a06ee9c56b64d39c7408c68625c85f4a7182a6c81e63642bd75eff388496043543b826470f3728a9608dbf6e10ace2fbf7d84dff3eb26ae3e00e1e70a2226791f7933b2d17ff0d0884902368522cf880de2b7283d577109d398b6e4084f2ac112a7cee7d80c5321ddc5e3ee16636bc6335506dc7087d514d27a3f8816ecd4c1af6dc514d19880b031eb446dea23a1ded518fcae76b63484b4d3af63f74ef879d92625c1333f8fe4d1972a98c341e55e64a7bd3aad8b2a28f9ce8c020f18d997d92e92bd34b7161bc54954ae7c3fb00cf24e5a0722da142c50e1880433e19bfc8214498a6638f98f187e2c339f2b4daed2a34734beaa03e7525f4283667530e2f43aec859895f171501c907d0709d1313415e259b4bcf2e79db0f5eff1f353d91e927e3606711fbe832de42e16830a0d81991290b6dbd670c242d8f8b7f9c58c51ef98165fcafbc41df08aa37af42b1fcd948b51f0d48fe844ca3ffe899fc9716ca8be0ce42db78ff1efde3c5319ad48654609914aa6e6af4ade0daeb71fa5d739381da16363e79ef34e0f215ea7ae95273cb259d34ffb879695ec81dda94994e3d0d2a53c86953c78b6d656378564eaa2c5011f4cb3a4e6c20d19fa22a189e8616e3adc5b03e7257f01cf0219203d57ba6bd3a010cf1fbb4c8357f48211968271c831d4c03f72d46ba4afa34e66fcf997aa3f25c34f0f8c1f65031eef7b6333797a4f1f2cb3e6cedc054fa4e3cf2f4a95e86bf020eaacae09a8da856b8fc4779e35ac9028bf02570e6f8a708e3ced49f2f1b42d8c61a476765ff6e90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbd2539d3fabdbc42d6e8063e9c885e5d8a52d2197423726c9460cfca1f49dfa7fe40a7b4fd07801d9bd089cfa5be3a05e0c4a546391ec57587d6b1d580f91bee3a6b9f5cbb3379d8bb460a276028887ca8738e45b4bdc111557410671410d06a650ebd4d3a42a075eca413aafb283240c41a29e7542f271d37261479867cf64248db47ce19a8b90cb3dfc6c381ea27a2eb73ad20dbfd2dba5b91ad006344111ad99842a2a2963c943dd1c2477257864110059f45f0234714d644640a94265906f625c674bae2f3a71f492beeb97248528aaa2e9be0cb77af4809e58c0f1835b8d10fff985beae90b63575b270226d477904f5202f3a6fdb3dd3549de04e479afaa569735eaf906ba7faf180a3b642d0c1e8ac66451248d8618fbc26af7bf426fc250ff0ac45571c243a00f689ee63603f984027f730430c607412fbe4eb4ff94121dde2316a017b9e1214498987ce20a4d3b76c28bae56c1b8156136459b67b016fae63ea52c5465b2ce64a6984a6d2edd7ca10a7f82c0cd9108be76caed749637a20dc73ab9b3914880f6e75b68acd073b866b35eba1d703f70e434385a4a12280728be13861c283316d5d42677eb51e312a0fcfa728bbb09364de2b586ced57fe59d0bda5568ecd9424f49e95f31e797d2b014aa21ba80ddaa54a40508d93edd0aa48501ed300f6d7643c94968f52e6042d0abbef12f26a50e0227795cbf8d2434c97fa5eb08d4452ce50fda0d789fb6e667e3809706f4e832bdd94b61076357376870a42147906a355c39afe60675c6d276d016e51026427e09fb8d3f724fce36e1c897e7532ebe7d39791feff472320d2e651da50ca9c987693fce08625057ade69cfe25babefd32d5febd5f48f88ec907021d62dfed5c79b530da54b1c164d3634189067f410e6717c7096ec7878a32abfba5cf500dd05f6df9ebbc6873f2020cd431a705a2871da9c82917c71b009a6394d609ae4907a7d4a3a09a7fa01a961b4548c6a85578c6fb431b29b5fefb67959eed33a1252f830b4665d10ed5eef021810195465d88427fa6fbd2dfa3371533c6b68a0e870b0b0a006ddb998ac198aaf97066042085569d92029af7ee1dc60e99bf77b021019644cbdfcc95cbceb529c2b3ebb166509b5d018bdc5517930d9b0636d08dbd90895b3a606ce92fa469d83b971684bad3ee9758eee661077e2e82b7c1c8112d5224b0c4bee9bbd0105965a7c9f4c65c63901270c4c00b7b0a7952a1693f7385767321a7b273825164b1647665c5f3c5207e4c859594e025f27dfd622b04519c724961ec4f000d813cd0c69edf21cb348df4337a7ba3834d3de019613ead47ce63e183493d85839b5e8601ac129702bf4319d5c26208f4958560fa17ac0bf2d0249994f28150274ff991152e011e9c5375b90afbdbb4b4326e4466fd921751490c2464db996e45ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4c4033507370a5c9552617b675256c916e158b2a90326e25c9b378dbde527c6b11730c0c27c554e39a5481d1d18de2bcbbbf4594171790a86a9d57f95ecbfa2eaf834e3cf82989755446c592108e3338bb021801ebc77effbe1e73cc4bd4ad8cf49311eddfe200c28c15803501888938df29b1ee7904a5704762ab7045e06dab2ca3d96c497d434016b4a09d8fea7a4306f734dbba978820b2c93da6f05d3473779c7c9e3e6c64310e62455ebb2dd463941d89a2bfc6b4f1abdb4d919119922b82517cb158b1c4cbf1ec7a66a01e53369e8508262f2fea5ca5265226032b1a77313b55e1f1540800f91736060a4af923125e9dd5f2572fc1a525c8d875c2c13680a6877e6b970a13cdd9c4eff92727787e80e49dacbc3d8c7d0c80d642481b70fdc799a420ddf96f1882f133402136731775d092bc9fab3ee395f1b31fe5b28c75dadf3d59e6f686b53b1776ea551e19f0a6c94399a78922fd1b326edce08cdff4c24e24c95a388af7948d948d68c2f423c98657dd9c1edc19cb802639be661b05bc4188a69a13848ab90a280a58da9f967423327f30427c0a9c0ea648e94a0b3601223ecbe77d29bf44bf239793d39fb4c3d5d66122c496618f0d1b86e1c37f44ac8dc2720bce46390ec584da8a0888d94c4557bc8db7908018795ccff9eaed6d7e66547aaf5c9a856d60ecc591b3706955c11e66f8858e384e4def7ae98d4d705e33aac89a7adb50de74d7fe970696da5146f87580abbcb9d4886e74603d5bbc087fcbe14f3bf3cec4a4fa4457c1118a1660c055479423335139b4ee090acd84876c7e0cea2bbaed4399cec7faf8225c08d648b6b882dd262bb34b5d1d2ed7d9ef7bdc562bd48804637ba98b75c86800447618931ac4447137d9e1f03e02b96bd685949f3234be8b0d77e0720738e8f2171950f034bca5d830af74be8b4b4e4b38285f420681bcaa53efb24507e4cc341c969aeb281ae00ea8e76a2fa18f64b7977574478c9032805dc27625291264a6d379520155372f8cf1da6e4ff2f36d0bd0281bd057e203c34e78043caddd5ccb33a86541f1ab7481cb630ef32d21509488eb992673a0425319352b76dd8388156e928ed2c3ff2527886c54f5807d0eefb5e2f85bb925168cf33c3c8c212fae1a581cc9a598be70778d101fdf7cb36625bd8089601d04219afb73e1ca5d2be37147154bbf864c4a784e8f04f0925282dca8b75146dbf5cdf37e8d9eb39ddcf2ca443e647d8df4fd2d1b2f4766b2ef1dbdd86caea72998466f784205a229920b4c4ea3b9c7709166e84ed39642ef957b7334964f52b452d8f33d8565f528404eea9f4fe52820d1fbf84abe45c143483f48909eb286751b6c2d0e74fe1d677ac16c263a58dd0a1d71f31948115d63b2bd6ad7c700315f403a3da0e6d4d2990fe2d0e9e1e00c0818a34fdd6032df5ffb02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbb9260c28167181dc2b7e2134e93eaeba51c1229434cc494dc0a13a4afbc74fc80bb960f630ff217541903cbf9a94bc824654b3c33ecadfd2d72a49f7ec3dbc7e9dda8c394b30a55bab46e5bd9a4c86499a5b3b2fb60e2ef77ad7bb11378621fa6cc4056ec799e0ab1441ba9905c06eb4d62407d18d305c38c9fa1e8801f36e940a60890ea991ecc991a5e69d21ff3856d2a2a1f0e1dfa8bdc8353bdd52d15e3e8bc688b3606f638cc40d14bf333f8934a6525d5ed9c8f22b3426652f57934790d60b2c15d4c2d96d792c0c624be18123698ea24aab5df3208a1390f370c0382ff257dc6a8d3a350524d4bb0808896395cccacf7051d98533d48bb705d43ce5f7b65f38572c1ff2c0cc4a95d4b6ec2aec20165a6135df7c31625f06a49bb08eef0418fa2c082b612fc42856c203e66183f05c7bad840166f595d4f190d696e7cfcafd4adbe69e04ae3f5eb04273b759ff01cb27d834b75cc81ce5278ae92b64c33a4631d32f72992590b0755dc5690b660d08722684c0b06f260d83f6885513c0389973fb5ea1a8e19141dabd0a0b25b2ced6c98b8e0e982a3c45bb280f207b3c93ba032139594b1edfee9cc3010a1cc0e4f989539129b7bbb77143a5d9772456646e7ccb52d6e53e9140909a13eb860a9692a61d8338b260330417830e66e12df19df59501316950f5bb2130b21f26fb45c683da81d6bb0b3793ee2297e1f318de4968dd8a66fb811e8f828ec7599a28113abc8db54cd669a625aedd9abb094468f1938bac0632103379f66873fed7d19388d75ce181fcb373bc588e43a8c7ce833ef64c1639c52a21617fa4a22ddacc2fbf9a5bfa405628b72e3d19491f9201f80dec937a3622bbaef35f6ea9d6262b2e74c0c873d053aeb0b339ec0ab95d2335b0a9d18aa9bf6249ae9f03067faa02eace88b0f2fa1db2c3c842a8ffc6ee7e7614f08c63008779fc75b243db8c8be90dd6b373a92d7adfc6be05f4e979fcfa7537a52b5132e5c526dc919619218479d0f0a84e8d3834a844848461a5fad6e1dcd7c74cfee726501d1623bba369c4ad68185f1fdcbca1c2e85ead1c4c4d048846645dc0dcbb24bba586619b8dd4138001aed74e45c02367f8d8b65ec8b24ab8839ec26094f739fad38fabdeaab35c97539a973ac8a621d6117af5cb9388f57a702b9d0b41fbb10a74bae90e3f2142b9a4cf6290a508ce61f088a276a86630a7ef335e1047c77721d3f3bd5e853792b471bb16c2749e9bf2670564cbeb9716a1fca7bc69dafcb13feec96dabe5a52e39890a53e4b6e09f6fc353bbb79a7633279f447bfb08434160ccd6ed012837a8594ac5ad17035aeb7afed467a4f090194ab6757dc916c706bde3c9b6571d92a0f1c28b188a24e4c0892c2a604e2a15424c8cf852631231d5507d55699f52bd38762e5ab070d0727ed6ee71f92d55cf53e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6276220f28cb8c5a74e6cf5b3e4cc8ae0b47397c5658238068b4e507a65dfb3846aa16e790272fb414675b5e6197d77a0ee1a520dd9cf61d487dfc144c2f1ececd7d75631b152b40300b87848962313861c7dfee8b2b1e4e4a649110c6983dced228998bec008f823c2fb84361d354accb0af70c2e4e0cc220977a48a772d4b3ef6fa01599acc8dd09de0537fec03898ab5aef79d2c09f6ce5564bd3767bc76f2c3336b841a97da134ddb7daefe075ed309f03e5e34c4dbcf07856b05e99239b436ed5a5f9299ed8794db95388a61ca712f837dd9b215711a7c03f28e2d75a0b21d9829368fdfd36e919375c58f6d98bf5be4f370d506be088bc8110bd07d6ec21c668cb6ddc4b5c51741307efffbfb2064171a59423ccd0e2fc7b45bd86452bc039c0219435497bcd9fa56aae1f9375a003594008213a8470c4ac1a92c00e2889484af4f151049e86f7d97b9c386c4547d05ef52ba9cd1deba34f71b37e6e588cb3dc8587be1de6fd55bd2606e811641f37835a6cb00da32e0e490c9b2d28f17865ba7e8b97096e5124da3af9d870119eff80866b0bdf2de96858520fef45c4cd79f0372fec48a7ccafe58303ff8934f9d4a9c60166459f40dbf3b3176cd13170745fab81b13b3409d1fb16a08b28d051dc0af36358fd13452d76f69e00727ab3e74133d6e2a799aa37077bc18444b5fca010bcee41c4d8be9112b2317dd18a9cc5d8afb470de84f6100a99cfff978e62d8eacd8155a00d00b19dd57c853ed44ca5f843cbe1309b7ce8dac77ee6291c90cc54ebef48472cd096d3932215d5f022adab3e4d76be999e51d48553bcc772334137e015b1bf71d85ca64aae10686a6b740757383cc55317bdd46510014184997a71704ccd59ba46ed4a5b64b9118aa5623338f89b60c929cf14a60681c6b26b8edff5b4a7455d1ad921d646b1098604b278eb7c89fd4639511e3bb9613122cf55a814be90d4e43c941b85ee85b16ee12ec64d2bf85951abd68336fc10fe6896b3325d45b11e12c8d013071ee21f97a4cb848145ef6015ae3cefc85ffd672f3d71d82ba8e37cd1364254cb5389a41d782cb736ce7ee8e10b6d58bf9aff9b68caaec8790cfd902176caf07ca9cff446590c40cebd6a0a04630718cff853e1a283ad9bcad2f49b6feb1cb438445290ba55ce57b966bd2da1c174735a885157e88766ab14f22008739bb2865b0beed2865ac2b0d593785e77acdeb9056ebe3101037d36a9c704b05a96842ea46044cd75754a9b1b09045a8dd5f156b99a2047f570804cf4d958d1de7d8f5b2304543793da93e1d831a4319fdd754839b6353f1014eaa3e32a6209dfc47d750c9eadd92292c0dd98e8901025e9787fb7af2f2fef79976f1edfadfd1f5ee25e46f5aa168276ec294f5bf1652c103e7c18476207fe6e9ed8e8524f833a36e779451a152a9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfffdff18b9b0e62fb1b6109a1f06eea89e574ad2661afd5987b0a62d36eb8134900a449de0be26d75716d69b012f930ca2ed8993a89d88667203392138a02f9336c0c07311618ef9ddde18ffaf6a2b9f57653a561b0afa5d8a7ef8f9fe5384c551f8b127cbc964923f5580448029f8864d95dd5e0027fce60b70cae9d09a9bf1b13dbd8082d1134715a1a6533ccf1caefe5d305153a53a5cf6f6d2ea170354e7fc9d43592d0ace22b744e99752e53768831dd78208b19c4cceb467c12973fe88db2c365a9216972bd993ba464a723815e2c10c71dff66523eddb80ccdd3ed54a08fac79b4b332a55d429d2bc3939e5b1a5b99b65083d8343110b1f8e5c0c2d6de7bb747ed7f40e16b328861d2033ebe25e9444968a22095523bfc777c325325766a575ba262db4278bfc77a3476b9fe4f40cbf0f7b8c0364003effd85108d5d2421f350958088a2187ef578e220abb4067852b82d12d6f0a02d6ee2a0c743cdc1bc7a6282ce37f2adcdf41fb7e69252bc3bc01d263711884415e840e01ea216e74ada4fb17b9d34d6b40ae55a240b0a639c6761078b2741124cbba91f6eaaaedea3f3451d02b8fd37c7896a1baa8294b331382f34cb2d309c3a05ef874d985eb88a9bb89152f27af7f781f351e6b3913459296bc1d89a036dcf2cd03cd30aca2896bbb99d5bb3f11b9acc2999b05e785c6b1e5cfb08c677d4680ec3a3b6ec75d117fdb65465c2c83706abb65678d4c038f8c9856bdbfc45eb4b8fe782571012a065c89ea676ebc95742ad5dc3c4ec572c897485c4420e49ac452e8f8937d9038fb7034bc3b1b5e1809726f2270af9ef38dd9ae6e887373bd890d3ade5dc0aec4b5277d3a5fba44d3df0758afaf0f3f8ba22c78ed5ea46acfb6a2a168b28a419453ceb2e1f44880f214a4ab3a80cddd690178ab7f84c96392d004be26269f42d4bb22101a12a8380f3540825a85c320de2e717af262751fed4827875aaf38b3918b7aedadb29b0ca67d138016efcb5d4f669a599f1d9fe741aa1d9bffb47ea7ff5a88930889a9ddea553fc2022d3b3575d46f21acd9dd3128cd17d4546657193bfdf2697ec668dd9b2197922e395f2c04bee547b6a9354de3331eaef575e58d745f481fbf1ba30722507903c44da92f72573f3e22c48f16538d6c5304038b78f3852a0067cb7455cd00a8db5d6e7bd359e18158d84a1f3da30c7ab1ccc293e1d8217a62d55d010923a71a72e42da22de2dcfe1d34c6ac1f4cfef2f372a40845f385e29b36e58533426ce1e929d4ed87a2f91f9cd6505713ea03cc1230c9751cd24782f49507f178292b862bae91bc392443d2729ae556060e80e5088f9764020b219d46c9c6d0580e9efb4493da6d42ea44fa91be8726901edca78fe4d6aabdbc62a1c6f96e3f07fdb43011ccc98dcddde413834ae6af32a9be59c431cf847e67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4a3be159c72edc8d98422c5838cca17b530fd707d14d1b51b4f2a0bd07efa036bfab8c02536fb70f1cc6a0d88fc010112aa4bcc6b6e1ea290c70d6f31c916bd45203748f2ca8eb895f8bb18e3dc933d6be4a8866b1c8a78745026a6f4ac0d1b0b50ed0b7add4d57b7897138a3bd0cb3763fcde19b611adb763afe0c829026170859399b21600a913f85e2b42321ee61267be9bb774a8161c819c5cc1d1b9971601d7ecab4e1d4a6e4fe0d46bf659e3daf6d8bf1bea76c66feb984c254e9463796947a09416807f13d9653ff4d14ab4c19207c30ac353ac73563100f97ae396db32f1f3c6ddc3087747d83173c93c0aa2cc2d4b72cedfa4edd2ef430161056f693d9c5c1dfe8d6163443b5a297e6ec20d249458060afdc8446ec6829b8413b5937ed0ae070280411e3769da73ed2340038ad7c5814771a8519da4cba85515230d3c20079e80224e08db603baff9ef3d1dd9dbd03460ee819d4aae993d2243052ff9b0e7aa7aa189e30d571f395cb134c158b895b391079ef018343fca65efe44bb2138c01f7eb594d5c711f3904e99a8e5a95b78f05cdd459bdf3e2cefbb22f426327b042a8f8b1c3fb5d7a349c4680b7fbef3e85038159a15f0f877d5bf20df5d8606e84665383552637502681f305d3776dbee8b6403a91206ac37e9a04232fabc0d7e765e64443fe4c4f1a8b7decafa98aa9baf53d3ddeb4f5d87bbe7226bab9eab308c878b1883a214b69ec28c5dbd72ab678cddd14539b6bdabbd14139ffad495cc95d426e605ff0cf2c4ef39f021033fb3377dbffde48182cfc2ead829dc3359c98ee0fb2e89e95257471c71646eba557e58007ee59fdfcf66fcceddf8ae6937de8d24da6d4dfe2623b53f31e46716ef60b2900c6e794b88985d7c93e9dfc232b326882bdff1d3d648ba7e11967e01c12fab336a6b633f254e5b36c4427ea3a2a167ae2c830b7e3d28cc0785972e12e4d902f71add80dbbc28ed74c1c0a9e3e89f486eebf8844b212b183ae3d85200d91c76ee6fc15fbf388db96c5c9b7783901e0c9a021d82eea86cd1cfbf0ecffd98dc59d6f0b35dd5f276f68dcb79b91aa2163ba2d6864167866fc88423489141c711425b0fe9fbfcdc45752a7bd952aaebcb45ba205e4d17cc8bb963d2512b1f5293aca3ac4c3b03b6da5cc8a40059c75e88696d12a1ea24c3251159f6fe04b496c99d4e895aa45549320b06bb677c81347ece29750d2a0c75360f1a6f7fa44aea01c7cb3dea141c7c8e2b0cda45da0a1bbe7fd9eb94b35a1d1dfc05c5fdb077f0ad86829c96cf145c241b2b69252dd06d5bf336d1e5ee42d7a63d14211128d6e0519060d901d62b7b76d4eae1d3b2c79867678c37a7dd9365d05098dc70a63aee2050a6074fe14889a9b676be5a43a08ab08e773454acb963436157f61734dfdd15af768a9ce995e4fa3983d3687;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd7171895f15d3c5ae89703ecad80115e9b9cb5af62dd6ba5af026548da28d24274a71e17ab4a034717fe2da8cc6442ad98d10e38a068f6286fd7173741480f1e295613ade7ff879b5a2ef96d648c469400e5e0b2fa5b994d3bf7fc535df6a51cb4f6666a8d5d206dda2d044eac796c04f75349f0e970a225b525ad3852625d58c32853a704e96c6d8e0bf6e61d4b90ac635910604b59b171331030953e9c69397f3251c8b09cc0100c8a666787352bef048f9964760eceea2cb7b4e57e3e604b97e9b258082a79c4f439e556ba914933c42bcce5c118cdad7317b909daeb7ac3b525f6b989cc42914eadc74ea3eb436cbf17aea74b98aa4a222381204ddf5d39bcc61a2648a98c5377157b01a2808ac62afbbf141a400c2d80960b06e85ebfe77bebe2ecdc556d66a70804961060f491d625e191f5b4813e9508295c62d05bcde9203d0823fe8182f3d75c8bf6ac59955a48cbcfdc1c8741e8ec64cf7b54eb2e5d0c896926877fea9a3bb168d1ea608857c7486639b29514ce04519ce23762e503049c3bcb20281147ecd3425062e09d5bcc94c03350e13b80368b06829335ad3227ae80abace52ad3b71748bad5007c7d6293e7a87d7901c7aef3b0af85243b95acd3f167cd1429304a4f870cddc2021ee6041e61cdfee47c17ab012924a9cc7df444d102b7c719033b0bb5714a2f0819f378134e61ae03bf17084d51689e718683695edad564011203600b1f8e640b3584ca7b10fac98cf0187d0edfb155c8bad637229ff2c2bbb9a6dd236ee800361be3bff6a358089836f5d0d459ede6e5d8b4fe484933f935ccfc80f3aaee27f6bc52c88a9fbe76a0db631d3d5dcf46bd6f3b796dfda596b6d252a4ec120c369cf50dfd8a97931fbe6c9cb27a5b81f85c6de0134441c1da8810835d02ece14001fd51f5149afbe601568bc0b4d0667c4bd921389fb3360eb59bffad7383d3be7dd5d02d62ffc6d0befe99107b6e185fab2d39c2424e902b6d15adf474e71220fe592b467d957ed99e7ba032b050189f86f4284be3589953cf966d18e96cdfc38a0536db10b9f41fa2946f97cb1843b12e170539ae900c16e55b570f1e770258d18f407fc1f829b3e87f8614a15771d6507e34bf903766785a858a30ade0d81b3907c83ec950e470a524f0ec5582bac3ebe1811771299986ae5433702e393c381d6d806f8f1c5dae248e75a99104ef4fb54c7b0e7955d277414b88231d501f49efb04baee3c0d92a4c80d68fdb8f7fafafaa5709f1bf78a30d084b896393a7029b1ea4ca03f9d1f1996cd42b50c0e0df1cdd79bf0282a1fdd5eb414d182e2ab26705cb51bc28b812c966bb5c5320c396825510af1101b42b8f355a0d71520734d24d1c39daf9ef4787892dd9e8e4d010d882318ae49170f791429ce5c8393bf1a829276035d0c9e0b93cd295e498e2fba4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbbad346907e561fc23db47566df3b0682af1634d0dc1366a457d62bfca2c2bb5b154d45262c46336220b62ad8c70d2379650f61bcdd3331c7f5c0f8895752d307240392eff41d567de0d0472074c38ce7de3fb2ed553d4e82935ce69417fb8c0260145afc849b60687a7a3426a1c4020f804fb884aceb16a6c030308a5e7c046c19c8a2d335497fd91c9f170bdeee7f148f50b2cb243cc830ed3ba499b4cfbaf93ba862b9f7e1d9a59678b4ac628afb76145d387f917536636c78a9ddab6f5c0803e898df841a15fd5ebe4f5a93d3f10ccf3d7b31da25992fbf6c6018c4a5cbdcb99f24faa4ebc66756c3798e2169f74463e61daa3e4dad8ca694047456ba69a75d4ecf8956aebeff3fe519c78d4b4d768b4c3cefc94e4da48d3d715c051a0e8ac3ff3de9bda8f5ac08ba1f73a4bb1a517ecb243ec4650dedba8e9933e58b3b9d978b4a071b6a223b39031a411a7df170f9d5d20924f94c88c4f17a759fdc14ab5843759f112b611278eb51b7975244acee382a33971b4838e399d597c83efef693a5d5ba92ce5fd8401519d4189243fd330723184dadddc2fb6197413cd94b59c2a444aa6852e5c5125aa048556f2436510dd21606fca693b97e96d6868a1ebe747031dcd5bb2a12505b254b4bd17966f002e9472403ca14567c86906052bc302f12d146cd9918e92c3c3e7419b79a7e247d2ead579b4baf39c18d09b9a15c9ff7968dc58fa97a0a63f1fe8a7d07849cbf80200ef8358a41d6b45de77939cd29f301c17efe12e8465778406efde7775cc3c702c8ab8214f988846a700d4e04166071fbc7eb8eec16e940f42901b5dff96b04b8d8cf51d85b590faf9b538bddb5fa52929190e0fd3424f619d537d9998addfa62a711ee3596bb9a6d34fb429f29860249ead7b10105f7657c53cba6e8c96740a449cd2871d73e3d621b0001dac9289be909dffbf85876d1804982639addece68fd725ec0cb7387ed35b52392d3ed4c621f425a4ed152cb4224c3b6615e82f0d3f6f14d818a3eaeb6c195257111c379004d01f13bddc53f0739851ff9f603223e1aea02f5157efe20c25f372613e84c266a9de02fa6dcd176f57b25f2c9c92f5456d580c734a6d9f21306dd1244d46755ad42a1fc2609d47aba5626ea3dcc7b10786304432961c88840841d80101037715e1721a49898ffea539b64c01b44645716f0c39e51170b6baef76825ae2eebae0e37b97f3aeda5f56210588b0be7cfe103dfedc3a2f6ca191e80680b2a12880cb85709d71876351228fe29a3902a0d92efdd89595eb155c30f5b8e93b030d2d8c02debf0f5ed9885e2dca80eee31ca167d5058a80833f9a0cbbbb1bee472b3b4465a43edbf0aa1627ad54880e804ce4b1969aa4d3080480a09983984b710882450570485876081d7da324789c85b65d7a1682e12a97133079c6e63ee09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha04850ea49febb789d4c6091d10d207ebcdeb2b9e25ea1631c5af575c0b63215c59263ab5bfd148e517f3701bdfdaa027c4c2183ff12f0263396b1d41bcf6dcd8ca1acf2f8b1684c0bd4b237c5b86b784e998d89ddce16c61e495e13750648e13021f97cbd098c617b86cf4302d70a38f88c582ed1d70a4910827acda1f643e5daa34849c3a173c01cb97162211d85bf2f38693f5bdfa1f1a3372a3164fc07f02a02538562ca9936be5a04bf6b26fd9806bb9541e2401e255b78d476d8aa1a5ff2d6eaa2f1a4448567523ff08cc4920ab9731b2e9c2207bfb58782256060f4831cf0723622b0e73f37acb1fe1535dfb693edb14a3a49497cb4d1e690594d0858ff05248ce90b467eeb1681e591cfd4157643ff9d1103884748b1531c16c069a62ec7da8944695bf0c99e26d63ea10683ca4e1992fa242d3ef20aad1f62857107610f042694455ed594c45bea08cf0481061894085fd7ee85cd2ad242b9c5ffa10028e9deac8a0dc0122e3568f0185f50957cf819efa3a86feea6443d24f67729b454d17cb16aca1437e9274d87f2eaac9e2fcaa5ca97d2ef26a3f636de89e591e730f0e851cc187c797bfcf54e5f7ebd58aa5a71212c17e2085459696662a7e0311732777ea6198533f8477491ac1e27eaa801dc3532e10314929d06cbcd0549785f1382de1c2a007cd5c947ad83ce08e433965a0833f920ad232e43a2d1d1ede466af5866dce78c03f878ee7147bb2c02b12df0c28023fe86bfa5261e6540ce71c537a11e1167a462bd6d5f179a0f32aa062d649d3f3a90aba2a18d2bb531d649571c1e32f40e7caf625d7bc4699ccf8a9069916a2a5f0731cbbbcdb9ee4c166442ef667a033c418233830edaf3f087746a634c8f67fa6fceec406c9567d2d8b2bbcb39017df1d6c380a146c678feda99a3ae55b703fdff9dc65a4ba62f20f3086b29ccbcbeeb4f1f0bd36d53e08b99acbd10d1b378e3db13b9bd3b69697057b73b05f6787897af6d28091b7595b6ef56a17c84b9995b0dfcb05df5fc2c7aecae29c7e3b0432681cea633774869082d944f6489afc350f0ab3781ca8614e4f6f2629019f5cfbd4dab7ef967f4c60c5f484e6098100355e182aaf5cd663689f59069413d258d3605559d4f997987e0f6854d2272e4f769c868d979124e23b357159a8bd6d7e642ad955e609d5a00186427e2ab086e63e5c3515ad393bb28c33dbcdf95cc35a909b64824ee7dd8700a5c96e03537dcc0afaf1d5e7481296876b31f0e2ffc526346d1bf70829f4aa80e8c0d5c687f33ea23dea4eae550464eaacf457df42e3145182469c8182fd762a10fd116b1136039ea13caaa1180e623c680cff3baa31861c9b674dace73f0f6b423fdea93a80b53025076300d3ba497cf8495e37828c27c1cbfae7e3ea0ed1d89bff6d30d6cdf13b175c87a7ac710b4a2ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf32d27ed440f8a27381c642030c8e2ac5c27eab685d790efb7ac69f181519972ea36398ddb2a3e1292b7b2f1b1b5433b51a447fd01a13a8e16b13959f1e2b406104bcdf65a53e6b8999a806337970bc7bccebac5a8511ef355dc00cba654fac5c75814e03b3bdcc5243091a118a78989c0bd3b289ddc72e53dfa40daa83edd87b8a1c85dfe3fd19922e1f0d992fc4e1ad073a3388626d28e9d0f9c9c208ca12bf481731031cc6ed67881933e276caa6b5a9ca9d3d4dd25748b5b3578d3f15658d6cd24778d5dc0841ef0eb277c6765ed9c6cdc89d21188b38130c8a7ec2a0f8ceea25ebbb6b6f1fe5efd23a01302266e2bbaef60412393c48310653e2ec8de7672020907b44aa3297c46ba937313aa098031f49928b866ff9a2785a16c65ab92fe117583de7aa13009c9dcad43895825e39d086cddbec6369a94d534a8436bf2d5e49882d7f35d695a4e372b2ccfd092c574b9e5e9a98b521f69a045e4014ca963d1cafc85729202b8f6a7f4d94561fc6d939d7263900f42bbc803166718c7d0af95bec83675f72c2ef04b1585707dc13e2c024d90460ad7721a7209ca4ac9a8687a2604c69722a1775f0e018d8828470fb364ce3c5aebacfa97a1dede163b87940606378dbfbf43e490ae96fc33bc3e3b7506325e471b93dae45b3c475c8f344a29326e0310a619ec4ea0b424eaf330d0b1b4a3361a53a7ad085775ef55a7c1e7e5f571f42e921f1681e5319b1337e51c9df33bf3e70d0119dc7bf6f72e2378211cfb072a59d296e012a878d52d60ecb302ae5721eb708b4da9279cfff80d4cf993f2edd43014c3373cbc163ecd041d1051fed96ec4d45c96e71e10583210d28d4c5793c1b419f3540cc5fa6ed8936c2c5465ecaac6e3586a1f3ef6aa9dc02ca492ac292fb43553a662fd5bbdf0ca7e3ca11097a9d64a568d515001429bf270bc92c78519441fa7c2e4922f4c39aaa4cf3ee9f40b7298c1b06677d00581d279f9a0d2ea0768d6405e3396015c66e4e8f30526cbe0e4f57a411076144c0e2684bcc2a797e7c0d389b7959e8f2f1540ba2a2c1fb23e49938631b15b4c041ecf44ead510aae520aee1a51fb5c1180d063e4691052ebe6c0e6ecf5ed6e0e6c73595e5d3120c4dd13a8d5c51e88f72e2d16cad140b8214d42f20992e340c08e6e0cac2c253d9b4ec3f21fd466fd083c1f19c469f1e079f1aed28477c680c96fd90f7d6b606400366dd012036a552b59256a97def44d9f078785e9cdafc57d345c644b25d859584309cd5e91cdf30a5c8cbdbed9e89b9f8157711bf15742a7cd91381bdfff9669d2e7cc83eec9412b1851f90c0c6c4bad846ff2f9fec26de472ea4cb165ef6facc2906b5c87e329b0b8b218eb2925738460f8ceda4542afffcbc9cfd09088ab595c28ea36c51bd768a3e863276113e393a1acf14a3018deca84e2e74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf6f222e05341040f267ef899f939a5e3e2b76fa493f8d3cb3760a309a8dbf5fd94b6744bb73fdeaa8d3715115c9e6b00d164713f53a07684e1e633ea0a484aed3544f200bd6cea619740e56eb738320c763689aa2d138951451a8d8a9faf9dc5bd34746ee4300dac6879cf98a53d0932844b22cbb5426fbedba2873d57d100c3aae2feb99796c5bdc30d50665739c9fb9cd31f18a28f119921d62ff64852acdd49facf82bd7a44d8ca8393077713a1f217a547d8fd7ca3cb809b36d8e3c362350752c1471058599a434310c07ae930e130d91fbdc6c4fde7cd139938b8b7803da6b7bef9a951d9842257fe5cab4f195d791d9139408aa57f2fbddbfbf8d3ad858d3a92aba1b086fe5412cdf2051d08789df5a89a35fdccfba7232ce3ba555a596b55821fb97e8063a4f6cfeb2f16aa20f18fa66f5c1b4cb4bcb40545529e1872fb790eeb35196c3a8f080c52d9f874b2c8c72231f509e9d4264ff9bff33dbefe803fbe0e0ec37c5b1ffdbd792205d5221032c87ccb6887be9a88cbeb915b13b3fab10d84d27b6766ad0520f6a47221c101b423dc89949556bfd4d1288df54a318ab5ba1d022bb6949115ed0e4f32d178df9b9c15c07234eda46e81efb785f34e5426c2c239fa24f09d8dfe1d2e55aece16162b0d498af8cf4f2f7b3908a45f1b268f8cd2a93053ed3409d019d53abf39687b98137f807d9fc4f9317795d511af7d39276b4b0c7c98e0e93a71b5a4cf711353a7beee99e132e0cd30fe9ec4d05315b289eb7e4d56029677440b41ad6b08c7f1930e7baab449affb1cd753a05fbcc0ac4fa7935037a5b02629010baf89d881c4f5960e552d552d468f6b55c64e7ef8384ab8852d5ca670b2c7432a3eedeb1b4e21bb43f9401cd9bb6ea6ad26913f039f89ed63944d74458316293abe1568bfe0e100a36b3f4e74f5c748afe9d886b7575730a0e0bef97dbd72841840fad42226bc303b015298fd01b2f2c4780606babea3ec93119060384510f0e8ca02fa69720cc63a7cc82cc952e578b50c3cebb943b831b6e2f03e8dff211a10ae5117c25636cfb2353da73a35bf789fa5e26ab3c180f303ba8d4f361e6be6ef761df791b6b4a17ba47e5c19f8d6ad2ff918ab39cbe8206b05ca7b992858a5a7e91f78002ae7604d43edc3810d7d1afbf44bdc52b46d992192479e0362d32b39bbdcc7768cbfc80cbc650d8b39decd7104c0af5625ed0cb599894b604e64300bf1a7a86b522ca4d45e8571dfd720d792a95f59498c581885abb09bd4a6233df31b7d4781fc83dd77203f069affe109d9547303e9733f79a99509adfe0a7dfe6b57cd3222768c7aa0db49db972c25d747e912b2434476ae3f6179cef759b42efdc3c771b2affa4a34c506852f57071a5e114460e8474c0cd2949df0cbdc77d7a673964354ec5f1b399f0d31c08339fd1055ebcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h79f081a5fd9a7ce1a64485287bbfbee5a484dd3c6bceaed02327fe9bb396a1353706d5d8369ee03330835d42837e066cbc41cc78d6780f2ba0f0f6589068de1d7713b10cb82fbb99e8ffa9158d7fecf3744e4dc7cd9d22360cdbc72202b4b2afb3fc8c0a3a0eac12d7a08788c961d4444753cbc4272f6ac845abca47327e45fdc9d350226cdb02c7e35c31c3441091c90d626685c6b870f0cb5af5b84b8717d7b2998bb25e4334c6189585c7e05808534641edfa27892ba986409e9920dd07265c6d09869e53bd38d454c2b42796868fdd867880214df8af3862957151bc36a3e37a6cecd5c783ecc2afefdec45e0b3c0e19c67e09f0ce99e2bc4d645ae5910c22a0e9a1db4efe808547285d6a33aab5d78db8c9743441fd59818bc41cca1496b3bee7275a2b0c729104171d284cd068f5d2abadbfb90c666590c2300f54c032a48593e2e8798df1ce87478a92cf98bc5c5fd7b09c2715c7357a489d86163ae736d7fa7957d3826e00e752b5023e9b6cfa68225fc4dde225df71bf30447d637fc822e0ab66b2a92f5dd7bfc8ebd03859aab68890587fc813ae36308067c3c0d83fbe7e9c4f798e64c8048cece57eff000e2a7480eaad1826573c03332a768e9d0e48adadb3a0b08b3c3c43205235c2bc1ddf708267c4dcc22e5b3a168f8973dfce1e49d3f853125c56cd2ce386d0ada4c47568786d4e1ad6eed29232188e72ff01226f52f3d8ad5ff66cf0877e429feea3383e7fb2dbba5219c4d65b1a9ddb18dcdf3906db3363461cd11e9e4c6bc97a93113e671da0c3c6e2241e21c004344c7db05382dc764348828bf223d21a37d331533a5a6d7b670fb776dfb59ebc4af25b298eb6d794ce09dd3239dd803f5db386662b61605e69af4d7041c9b98a746df5370cc9113b7aac9eb29aae008daa0512dd2145e5a2124e7e526a307ce1262f86564db3dadbabcf312bba0b9f8a3ba7a82839ca8d943b541b75101028c450b74497eeeff1913694287745987012c422ec76274515bbab8973a769009a7e99a787b7998c6d6f3fd3987a3c0448c1e749c21b2621cc246ed23223eb8f6c0ad2d2baada574cab8c3998cf53d14e88cbfd0ec20a411b26e44597f60d6696c34755cd629ebcdc68a5b5cb9d6631e60590192f9a8aa4b88eb4dd09403b8a4bc192d3d0233f2f44778b7921b50f01cc912ec84f7e139f6a7eec81332ff053dd436f9416e9af9c04770e1608b47a0e258050717d27e06c3574d08acc0155d143b3f3aa4a0fc5e5aa5300262abc705cbbc8171aa6da53dc8e51f011680f3c3e90108c40a27ef0503f23a4c771a29f092c36152bf37b469567445764f31974110e07a84c495d7266ba6aebce9a00e73540fe25f5fa928b4bf9162452a1e1f1df104c29cac992fddb0888a7beb646a3ca05a59287e0f25e0c8f5f15747e36fe2c24bae90f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hed27ca2ab162e603bb935fc0f381813e948d6b1a780f3bb8a71b60ba50d2b62dabc054b13cb7d22a994ed0447d59be0ce4d9930dd3830ddace8cdb336052b5af2b910c8485bbc48168ddb0eeac7b8a28c40082445f82f2378aa14ef4a99baaba2335c031a31a9a04e8dbc277d491766ed07f8a0528504397ae58b3a85bdb6b67b5d85d880968c4fde854a9e8853bf5ea169797bcc041ab6d37c5c43dd1f1e31fe1f00d8e535941846c828d6f723f72c80385dbbe0fcd97e38acad6524154cf965942a07409c29aea0b763da1b6f5cd7a8e6e2fc3f596545960cd2245a2641a7c02fedd5f8eff5c01cb7ee2a9ea046435dee285696cd5ebc89a7faa0022dffe550ce8b5a2891df64c6862fd9182b0b44ebac5e71343d1467c10a2076e61808bf380f0ad0bd45a42e3e65d52de1367249c3f99f48497c9e34416a6ad58f7cbc98c5255110d072738d123d37b09cd05dc427a19c1b23eefa4383b6bea2bbe08e17eeacb796c25e5e7d33dcb934483af23e6f529ae094dd4f9ffcbf10888002e325ae42e6222d93d51674f814c24b3ef53f6f6f96e3952c081e36a83702313b58db8613e8d81570996fd8a54c9baf5f7d1b5c74e9f2f86bbe18ca6ad9770908183d532cabe950f62c891d999c556720d1661eb27fa179714976f2cf80fba35e6b97f749e4380c996622d3c883e134bce1eebbdea36fbb50497b4cb4f839766ccdb632a76cc24b05304a1a2698ddb6e6823c6ace7974c0c212382c2a5d4c8b065fba82800de6eac4e52b24f1a8985ba9272c6d0257bc2a058236e033eefb7c5c23c1ac9749c7dfeee7e07984dcb9935d9f1654070fe28ce3256cfda82dd0ac55b8b2e99fe7eb4739fe04e7b67fc43eb24820b49a2b4ed5c047fbe5b3231d916dc7e825f2c315aaa6a55b9287931ae2370b05734787d363a75075c24532c86bc55676367fce30aca3611b24549a961a1829f5ede9b6d3c85f0eb459526c1d7e23cc2124dcce18b554bca04c4a2cb1903deaf3f5d441d695964b6fb1c32e124049ac69c0514cb95cf31674259701f366d6400387ffe34f8da304a8690c3b1620af5c70a1f4415dfe2c44ce7f161d5ab5fdd4d3f7e15458c53a39650a770860f5fafb42d3a5fd63917790e2f3dc460a551182f18207603160fc719fd4bc27003bdf672b1e20524b287fe4859a4d2be898feae0a995ae73e55b5a591fccfd3cc5666e121ee3a6d095aa725cbc9ce4b533a40fb5aa13c009550c25d3c46aa3382432b1033210261937dcfb5ca1bfd20c1fc65050f1b85e077bc597d708944d375bc42709c1775a37ba63ba4383151794afb94e5e4b4322350f3518ab46725640acc87a1e014aebe3289ec28d2810fca93f8000b2abe1963d805ca867d46cab1c58a47b4f87c583f73992fac014ec23bccc34c937bc5117135bfe55b18252ff29e4a4998830;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5f2a69830d2f9baa2a17f8a678a33ef8237bd590250e8617be630bf4e1d46e59ec1b99e1ea30c6302504c33253797848f9bf71bc644bc1baba10632e436c1567a264ea1712efe02c70caa3eacd74142b681b0ed4ada3aaf5fb7df2bf96d877341a365b73d5c51c004ee899827e67246db1a3213d8933212e9ebef27972fcd6857bd8d4331adf09597489e4656b1434a1c9ce3e210472255293c5fa633abe50649cbd5869c8cf708ba7d4b36dedd90c25dd56887dce5ecff1f3b00a2e9277d3a234330badceed71fec6e2a9855c8a9a716b4b01f130a863bb0dbae7fc4c9314a0d3c3cce99fb6b6788456f23b9b5985106e3a419ad4649fc1b3800cdb3877b1d0f18cd41888461a51946b3cb6f880217da490e60148c9565546e3717a06812cceebefc93e3e16ddc9d33762d52586a48720f954dbeff2a5cdeca6af76c47ddf6ca421185f3b359488059fcdcf36c295f5af9159d38c227c79fc0f4f30585804445c16136451d72f2f4820e93b0e758cd7aa2d7a9486bad20cf6d1aea35e41d7e020bab4662a534b567d04eb47d1582537fdd6b069618e313a7bf346c74b24848f847271d257c38320ef29e994683da29e3200f85a5cc259d59807226a03b8303eb15ee7587a0fa482e1bdfcbe6f05427d80a516a771ee2596ddf434260ab4abcf9b86a60070e0770f0844753231c0007b6f8ee1c692e58f34f76296e7c5b49d32e2f01c95aaadd19d1ab0f89b0806427b76743c8e23bf9e780af7baea6594a1f3d36fdba8b32010a2a56582cf87debda15152e5e7afa3eb4ccc226a5df1e9da6d3725c1959ef66f57835ad0af16919bf2fc0e202b69dace732ab20e17baa9ae67c870892ae1d146bd398df84b12518c89c16ac952550cc459cee70531849fc34265e6c0c5087b2a58f1acf62c33e9a5fa69b618682539a5ff14088530a1e50a472a908d8d49df67b4a86a57926a6a4863e7524edf85417932268ce6b36bfc7804fa523a16e719c1dd54067fe3ffd7268742218ac05a987c66d8572f5488968faa34f45d40b525e0a4bb6167231c02a0a4aa539b0b35a7673ed2a17e014e5745d40f23decd0973ce7bf3f5a658609227640942adcc8d705a354a510eb88c80ca63ffa72d2361216a08c4878b0681801f76dad021fabacddf69503c740d56292a405635a4095c3dc7f50c6263056b8ce1920ed520109f4c65c9723c13d90f0b7659ed4b69649d502e4d662d955ef6ec2163e696b9137f5e6b1cf3c36250011bf0a43c9b6cb001a67e2c4b7da535d5cf5ab11de7b042b645d9293b4b91e0fd7a1e21f8ad6d25f76d7b2bbaa482cada91acd02220e09d77cbef73b0d7b84046b4b87354cd9dac346fb6080a927c1584e31a882c3c65644bf741f980c21152662cb2f4fb9505f8498360cfe34059b35f7e6386be279c35cbc44a7b9fb8a9af62a925da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd6c1ee75b78f62c3327570ad8cc2fa285cb8e943cd4adfab6d646cbfe4993f475dfc6e6b1939a5a7d176021fb28c845a7463f89a78a94e25acf35fde5d88abd9d2f09d69ae86fc4ec3e08a240d98888728afc706d29b5be899f9e385bf5f0a3138efbb4c042208a1897e388d604c7b3d20eda8075e125eed652e84fa36d0b7394035bb927015c2207f589caddf9ee7a333b9655ce82f2f2bc30e9da4c737b76b084a5f4910f275ff4fbc9d00b146c85cb6da43412413d97505acaf04eabf8c3a2928594434e789ccb1edbd3adf11a151bb1d60bf5545634285cc20087a7ed2b3bff8716642badd1323debc19aada49eee9ef46bbb7b9c244c0fcece5337c8afc88c8476051d5b8970950a34172907d961297601cc7413e43c457bcfeb763667c8036c244fc787359064864aec6d29cbaadd6433984858a2bc0049619f156df1a4f37603cd690f39721fb690fd7d487aa071a1fb6417dbfe2df9087d073be003e428cfb98ebaf9a040ca32c16a01f9241171afc45aa2d02e581d055699330ac80000b95a83302eb6dff5f7a5d3f9de9590760e9004dfaedc780f6c6910ab70f6f042820b652199754b565353ef1011e068f9851e062f06a031b3b24c495f6f0aac99c07e960b5e56740b680559969ef7dae85ab9d9ecea99d1d3f4adc7c7b69f206dde5bbe2c4fb965f8ceb98299cf5f33d87c880168da0ef081657083f230d29a9a88d6cd162f22cbbab47707a3fab9f8493dd1af970be9a913235179ca1ea4afa873c4934a46a81c31ea658df387b0e48ba4c9073af4b90ddd695f4b449511cf277cfce0f3b65563a84ad2490f7a45f95c4d12d17fdca793e53e045ef633d7b634821987062017a98646e45fab544174d5760d478a3222805a004e89fa2458959da9f981b8e2ac881cc26f44a81115f9c1c14067ec2c35dc88b102d786f9394d7261e0b8b49c9a2bf4386be18db8aa86da8b2e99cca5f2214744f9c0dc2c4acdc82a4632e2acc8f3f642343eef5e89bd1abb46f31424431afe53ee6ae6514ab353e11efba31bfdb1784a54d6557c583059d8b214e5dada4e4c0efe37c4c58fcccf9d05316d436a66039a2517546babd3af16d8141479059aed8c4e1aaa964e05c4b3e5082189e0dd1dd5026c886630cd021c335445f4d74dffbe7c7eed3f97fa30ad80f07efdab778fb24a8604c2f889f917753aa07c0e34cf5d3c3722dd8d26455c20f218e1bd6efa25003ae6fd65e4205181937d325f11a615980341ce0b29bd248f1d24bf52fd5e6dafdc16c030f0d0852860a30f0064b5ebb1c89341c8d9dba7e0fcc18f911a5582f9174b9c0a64d7493f6eefb8336b0a7770ace30ee2ab466dc875c9a61c8e6d7c98ee4e2059ec41fba036d8af4d672a02d1c7d294b7df59ff0c9b8cae2e7c50c22969d18f7bdc8c724a1d8cf5e306d350bd4cc78e7b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h701a90ca598270475354ae7bc55bf8ed2d45dfdb1ebbe204a9962f97452bb288ca00712b43dd61ccc05b21397e4374f6359e6eb63de20a97975e614c400294dfb762ab1df4b15510c30e6ce182de1f1b38db735e8c07277b67ace6fa44470d08162452ed47ab9c7e2cefe6537ecae699a4e028544d3b26ffcfc9b39c9b6588a95db27747d354b4276c2133aef770f742c7628f82a0986a3b21447ea7be2b1ebe253a744e7231bae872362829e7f679e90a29d94c9b7e69703370910e6689f2c9df1aa117a45b19b3c1dee0616978a187ca0772d91dea767fda31177bcfffcf5dba7b3b1d282425be52c5fd5bd2fd834bcaa69070e4d8083696236e62ac7cae7f70aa2be00e79351b6eac8aed11fe339e2ee47e136bde91a049679f3b415f69f9a1daa3f9d968fbfeb5cd81cab464e816cab2f63c4b795c76632fa45e729cd014b9f13fd68ee4cd7153bec1f72177f18cfc0924e3038f08dd52acd0da12132ebefffb1aad1ff9e3b09ec55f106c0d9805e2744d6759cc64831bd8ece63d632cd4e67a14e641d641c649f999a22ddd686f5c929b7bbadf705d45d6f2c42aac4b3773258931ed14112945a787280862d8c0022d1316a0d8cd1ac1e0acac8a915c05343393918500c1063bc00538c94a9ced09c0bc267058a3b2e01ec1149ba0315a498deb01485c2b481e7a9362662ad9e3a14ac2378c10c5b9d8fba6e73d35b9aa62b5716ebc4b3ed6136dcd6ce2d307829aa0ac047ed7f426537811f3914da874899007c8bb3f99f1dff96d87762597f8760b8f1f021e9d2120a733cb7ba4823444a148dcdd878926004097ddd1a22fb120d3109f54b3e764e3852d7f6f53739c86c456962f7f2a562a02e196e150e854a06ba73e939ba9442aeaf377243d9e1f2d264e4787af91af6bdbb680a597b3be8afaa8d57fad79be8fe7e03de6eb164003379ef092244f62216220818060574485435aaf0f83c346b927c433582b81b749556a5db5adc908d287816281ae1565f1d2d65a4111a93d47f0e9410ae909c329047a189e3d3882d5290664bc3b807f9324473066c550b01ef521fd705ab6def969a0b2e0d4208b0ff1728de43adac2861484d102cf30b8a11a413a3bf5d16721f2b33ea510090dc9811b583646a0fa151e8c7f8dcde3b9ce570024dd0ff21cea068e7af015df54d95b75dcb7e5a669628d72f0801400bb8208daef5da62186463be83a579f42752105d2244ed9a08c2f5823175843e20ce642ca508af6b0cc3618c7a1e8e7530e9bbbd8a281c8928ca5c620ea7e235c074080089518f82ff4a7713a5efd3bfb62a59fe52b955c234a537b1088d9f4fe2a680829541a3ee84cd488639ce5738e4be96eead693133687cd68b670a2ab1767a8b62fd5af6533e35a38402ffb73fd708029485a143e9ce068b0ab1ac272a43f4b0cb5d803a5d279;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h55144465df31567da6c188fb5bf2dd8222fbd46f0e1c9d24c63f06a31295fc6b1633b341c5d1bd36be75103a34b03b829180008745b18ce0c049d20eaa245c3c2c71f2346b392471f3a9a12c12baca7f8d9ee591f075e33b4d94e11da5b544c64dfc86f99b7dd47a89414f27fdae370d73595fb784dd52737fbe29fa071d0d125231fa4520363664b8a853435913fb28f0a17442ca9bf8ff355ec70f11266b14545f7237fd90868fab75f2deb41c26a599a676e648aa8ac0bcff181fc1e341658d41f2bfbc9b92b4ee8238393b38656f8b4da6afaad3ba8c37c3de484350fb6b327259de3de7c52e1991d2bb4c0eda3a405332c42b276e1db3622fa5acf986f300ad77bc759e495040a0d1410ed00cf0d22565626d1e5a3a6f6f02f9e0ee8c623cee92cec1eb08aed7580bc97d3e739beb5bc30816e0915a33e1b06b270fec5ab2e29c60d6438fbda391590df16ed5b503837f2d7fdefa12a41666f40fe698f626a33706cadfde90bb70590e95340b2b86908224d20c78ecfb94d577fec60dfa66a061f968a6b4cd969ac6fdb7bfbde2381f56fc398f5d491cf18e20a55107e641b5f024c07c1d9642b0e7eb475fc779fd5dbd245ec0f28d2486bff3e95d2f4e6dccde12db1ec6d436c0247637fb5560c462027fbba0e6eedde0af206f643b02e5d7194774cf3c41e56b4950b05ec65e31db443594307271e66dcd2bb0409d4fe2c8ed562983a43a9271a7b059fcd1c50b4bbd520e6cd7ebb165d4b02318cf6aca7eeec58a556e85c6b9493cb2047b5e506d22c5d7450e34e0184d6b966422df2de169924a173bb40ccaa79577b3858d86ac21b95a0144bcb926687c88b78d8248ab0ec6d8a87a16eb60d2709bf2aca3bccdf505a2276d524d6d6f62b59b165ad8382f438fab3cc15074a2e35f3e055a784f68db6cb552bd479d205b30c9be80779fd33edad56fa00d2587c32964c3219e616ac3eaf3ec6f572cb32bcd1cbcaa0831f75bd5d16c60e7871847a84960df9e339f303007822de7ec2f5d94e35b90a5df453455ebc608bb4b59cb48f7c81eb82d9115f619d7a8fdd95b5f2ce17655a950c416cb6eb7a755a63e7415aa7585883991003f3e29f02a5983afa8f4ebc8fb883c3a7ef414137ae10a58e74bf7a806becf4203c175d3e4303edcb5955f68201481a5992522c980d5ce2db99e06c057445cf5324ecdd9acbee75a092378bfc2af1f13fd6f9b1ce3996474c47b32c92f6966fcccffaeb82e7c1aaadbc9dc9d4cb542c8c9cc823529701584d2de8b484841dd82142cc6192bf3dec5b40a907001513e5a2c5566a60312b2a1ff936ab20b3896c57f4e9264dc9370f2fc6ea7da0311ea36506b7b3b01bdefe167649eef765f2a4dfc7260693905f1f8bf0210d4cf9445d8433230affef63e400c41279f07d098876f0b4c2f3cc0a9c9022bd5f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf7d904ed6ef623c536716ef2f57ee15986a04d518e4c8316b126965f57b618e671e7e7f372ab9d6de2e8f2d134df7e077c65ac72da2a7d2d61ca091a3c86670438893950055d17aff58170a4fcb180ae2c7220242df0c9d82b7456033a57c24bcfe90d795ef035393bf719e45651f22751dc8c859d1a30f3a88897ff5a2e96423728fe3e20bdb4f1dc7a3d34fa50e54df1180b8083e43a52ac13b23559632f930366f991411f59910b03a65a40b9fd9fa3cc9f659479e5af82a9dd544beeb7e7528e6f91d7e9b9b7df31ca253dd6c8258e4e100a967b9d7787737de20e7276d7908d118b12971fcf40dbc1108d9648fc95b0553a93803a256cd9c52702c0d23d0d193d4b2e8986b13ce8658bc8f9db8eaf7230b6c885cf76b4ba382a2333b0ad6ac3975e616be69253788142258ac93c22a9dbd6220d2d29f382f3b440ce4fe99fe1fccef385959eb5504c4c0de41ef1d057913e96238ba9a40800b206748e01973057eeec2bc5fae8c1da724a91aa7c29d4c69a3af267c63db1853fad54df7210a9e8ff5d8e65fa5b433510074aa0fd89fb90d8c25c17be2492afc09077aeaa59eb950f08ac9b0b994c2d7fe6f8afdef91f270c25c8b06650f7782e9f1eac40dcfd131fbc9081f4ec9b2da53916da1c0079ab1550f873343da860c5e1c417badcaf3b572c6b0e9f63d6acd21b58158d2fd5b188248128a9abe09c4bd8652ce7e740dd424f5d4b869b59ecd4efaec1a05ae5ec3d803c6a42221dd01211817082c862662e9a82d835bb48497137c76d8efb41f8788b8160654169ce3a1b4a9a48ad3c4f3c492e6c01bb0f391f472ad87954ff98837da2615c750c76be33845f3ffd2abce15ed3a2901eb84a6075a2bffc84f6e0cbf4519d1f8db758c72d70aaddf49e0e8ada7309a73e757799eeca3e5224262f3c3df98fbb2baf749d05bae38f058d5609707c290ecc23cf2b57d2bc2e925168075ed55fc2781312a2538e2521f305b7187d39f06258651396115df2d8c1d04d33e351b2089919f2cd1fd84331ccfb99dd8d656371e41fc7b854de67d4d615a4bca91749d3758fecf925920b217d5ad761327e32498fb36d2f02daeb3fbaf7e855265919f9b10b42c48d5a629df8596df748f965d0b332590954abc0b477eda7a04056833e01860ea76153fe0906a62fa9ce7155cb5934469bd07ee0af8fb033ee0c8d5045237158299c828e3eacb7555415118d16b1fc548f5914baee205356a79aca4730445ec649bf8329edc98b8b039a4740a16fff9d8187669588b28eaf4860b94238482b9b032ff5260a028c8dfe2cd0f1c44c7c7c563973d86dddef0748cd146b4e80a7578eb18a5bb6a219e5b0be422f6c655c88f6d61302dd7bf9ccc945045e3196ba84b98c76c80ba6155e654e2973662193987bccd6c4e98c878d3e7334dff419c293030f9d2e26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h42559ddda9b38ea05276a8ec994a44fe544e7178f0f6d6dd14a6cf9c013531fc306ba31eac0b4e8732d38a7edf8c14a2f9c00766abf1e82ea5b24eac476d40f980f9c94bbbb78eff9766d9578901183821df15dda9c650447e2adc36cdf61b01333dc8a50bd2087f086b1a493954743d3f7316b13c5c9bdf403f0df2a2db801ca1a187a132ff8f2f537bcf90b388e3c8a60c92a89592c26df8125b240f6b8a1d76f162fba1a1c95b5ec9dba4e17c836d739f400f2818c1669feab68b602b42d134e33f6ca3ff37d7acefafb124c1520f8f9991e5025b376221373c9554191062a530709517c0447afa3a97a4f6fc0a9c0181ceb2408b828d2efe7d36f07f05788d77fc80d4b696317fad7d00156a18a99b7d9b602138c9815324101a8193266b32ac717a94ac70f60a706602d1eb95a1b75e7e5a73ccfb9d7ef59fc7cc9c5ac08849bc94227ef3b6e2d3f3cb5a3e5a1bd11badff80ffc0df9c91fa130aa41fec81af55fdab45fea2e309907aa4f7910f179c8bf95c9e1c1711c162dc8945f63cc8363ad310e67dcc5ef43fe24a0da1fc9be98b2a74625731f6e93373c9ce000776d5b2a355157e6a4b7c6cf003fef0b9e5185ea6347347198acf716ce7d69bf8f0794c1fd3194f25532311c352d7c66d152115d865c9ba55da5cc8bea0f7ec92a3f478ad71f95fe1f1df03f98b5d346d8137fdfda7813a8218c704ceb9e98961d2018e27cbf645170cc8d202a3d7b7d93e8250751e2e54eece9dbec00923de22509bece375a759d107b6a43764dc0917afd0b041eb7332e4c049170bdacbc8ecec6741394f994f9b79f9962c2203a5a0c7fa6cfae9b9b1cee9179c61d35b683fb32b11ac56d82c59e21c3d174460e9c641704125a77a7e5140e2a20a64b4e8ea82f417eaec998ea08d3d31b43d1c186dcee7bcd7a405cf0d062e30994a3671944de5ed0974e70a4b313512b0a2e7437359104ad5e071e9d611daedb370497c5da9cfd07c20f0e65b364f21a2b02acd7607b41601e7637ac2215b720d7a00c1280e1971976246caf58afea77d68cc02c9742f2e16e5fbe8663892e1405fab3ed3c67754bb2b99e1659013928bd7d1b59bfd34b92ddf07dad72ed86e77f32f9bc7c6fca4b436d834c583252d659f39f2aff90a0a55286ab492760724f1b4d0cef58ce4a00427bd8d1db2fd761c76e251bda10d8698f2e17ac0bc758fa571099b47405890ec5ed2f07be75591ec714690ff89dae9b457d4af67ea5646df62a489d489fd28728ae63c9a888fa550eb9eae257199ff2a15a5685294ab08dfd9183145965b44f7ee1e7a17c1ec61c60dd80a3e2033c6d7a753e83b84c34c06b3c3032d83eb91fb134a1e7fbd274b5cab9113155a9434678ab4bb95a0ed448a32e05c33671886721c1f895e04182071ac28fb06a65c1f5f7e5c507c612f90f181329662;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h379a3c91a82aec9540832b8c0efc2b03a49629d3ef43057a05d0ca0e632c8050246bffbf56bd6a3c34ce27ff585bb7bf3b8b317983f68d81cb57b2b2d3e0ce1e1fe1ee8b71b4c8ee8718fc90ca31a37a79d9a5bf7d07d47fc3548d76aa15763a9fb00482e61bc3444fb0867b4066a4718d008a635cd8c056e0913163eabe187556a3cf5513fe93d2a3e9b1e030915487136095a0e51d99ab3f58b12a268b300f2d697ccbabbbea61055c4680ee3fcc546a3b32479991087a0bd503eeae2e8832324cf04832891847bcaf106b912b520aca81a1e19d2e704fa70da6b445dd52105c1e1adf66eed615f61eea4435f8c1bacaab1e3fd0597eb69e9a7f05526a79b05310e30b46044089ecb65a379a4473172f755aa436df0ecb2c2b52090f9c4e72b575a4f610b5b512cd848392a48d5c92d01b9b4afc330883d24653fc0192165043de9036591b772f4b049f48327afec1a3d5a1459d51fd1cc225602f2fbf56412c8eb23c43fcccb5c28cd177a4d75e3b916f0008d796c2fa1724254dd413313a32ffe9cb71e2f45fc450098ea1c685fa26e8fa05bc30b9f1218bf36d84f01401a00f3e3190b1566264492c36d8d3660ea77ee434848d69254bad39ef3f8ff95667241b34099ac04f96e4e56910e6065f3290fea9d7456b5b6bd9d028d483735f178cdb588a91afc5b1f122f1ff71cca0257092c3fdcc089913ac79b431cbe064e027375a730994706aa4cc94a9791bad4c8f2c2842fb66725aa8a4f951eb3bdcb23c2b02467b11e864883c04df0827b0bf26a18bb76cbbb95da792cbd665600987bd1af4f6acd5871441602d2213f81ea579fa73c002f493250a646c8fbd0ff30c2ec3f03ded9d8a6bd44a872d887e45616152ab7e7529a5d5880779c69a669d468261e5d5a6131f4f70c9f41ee6498e729d56f9c3b15bfa47703efbb4add6d2e909c604e02d60799992737757001b5eaed7932d030d3bd6010895aea2721eb1e3d615179c23ccb25b2e95289e2efc0f2c117c93d45282120ddc3384d3e634ba5076aea780f0dd77f0cfcd926d2980e062eb862c68d43a99e23e2c5cd944ec0637862151dbab18916bfc16ee43c0343bed20ae0a016e416db8f0a3b1ff2fca58a229beb2af50842a5c7ee81140888b8d5d3bd916aa574aa615cc8b26371a4764a8c22baadc5e1d000c690af70b85fcb42bc4ceec4c326eed0b5b49dfc7a3ae1de58de9947ce18ca98ef35b23f1d8091e99bfa335c103035408d648dd60a98606bc722d2d0438ae7d05dd60f47e197cb44257d54faf9225974dd727bb2d8f899dd1fe83861f9a2dd7d03878c132d845b9e5cf3192c74b116b4263a64dd6e35926fd4c1a470f4527e9b4a3721aed2a2ee14fa18533d17a8e5749497348e486e7b9ad7173b62878fd64b39d581e5b2864c3bc1eefb7be476f3530584a8d592d8e11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hadce5dcaf260d45d69b904cdc8aee15387d58cf6ae57857d08cd28e18bbcc1cee86fe60009067a77abd4041121f2e3b4ddbddc27beb6d78ee4b6a28da8e46b0f1ec8d3d6901f3038e99e371649f56a0237f42fea3d660c24e4fa917aeee2670222e589c15fc18270b0e4f0e873a2a1dc66ff3c71c4a9058b1c2dd45c02bd6a6df09e0f8959e8b273ea1ff7824a5cce933a59d31ed40825ec19b497a1e6534d6a419bdd9756abf00f04495b692806f60c73a902b96229db3f327c377237af48f7f6132e084b413d8126518091211929e3f0ee2c414aa764916aac48812b6de48e35294089651aae1c728037a7f6835e0c3abc8f711a5f5b929c43b66f33aefe9ea49d3bb490e0493db2bb46fc6b38e9c482800481408c19039e9cac79d904b3f1a2c36e55fe2a517cb27bd92f7037f1fe0f8cad1a4760f47e1b05c18c060e2f271681ae1c27dbb20a2d8c5568339affbcc87df99921fc9b8b9b949698b44ddf53f5f5ac89c06f03c5cffa86c003aca25a85cd1494c71367afc409e123c35b6bb2f0eab07ceac034f1ccbb1bb9ee38097f8aa69d0440d0aab27a4ba36b550cf9728e0dbf6767b66f7fef19d855ff125ba7552854e443129429a60af8fae075238bc7ce86e44a05a3e22fecf79b58b8a296cde5ec2f1055b5c398ad6ab335d4e0354782940a6745d2d37cb2db09562f4582dc68be34963b7ceacf3e68d6c71bed812d04e7841fbb332f113f307a39ac64acd42925ffbcfabeb5020a98118c37754d3aa97e606024723f01a4db26a5dc53ea09e6ca524159172b5c2cfa0fa79f6c0c8eafc3fe87ec7878307ca3c5bdad60fe62069892f3de7634340281b8b2be5d04cfcbab5cac5d8cc14f4b1f8481f1400dad8f0c312d0e3602420eb7827c31fd35dc015f1a0ac1f9642663602881006226e1b2671cc4236367d2455eeeee8a85f55e6b14a1e6ed96742e1b0a7952355334e1e7a9375f87fb29f5ccef36ae17e40ae25db8b22c4296b6851e25ef0477a281b38bf79146e2ab411d8fe265a8468dfc28850081b1e212c86efc4c48328f5a3ecfa3bbd2e8c664f190c42a56445f1467da4f6b7c153e74b92b3108dee3e665224f1ea82111594e8328079d8388963f9c490c5f428801ff2a1cf8d6adff87fb386f581a38d610cf98db7dab7add6606500646ddd89df0c98ea6eb77061285acf02119c264edd2aaacc83da1a0bd30e1596391e77143c1e926fc50be2163f5df1ab2d0f2eb2d5f592305a245fc513025aafc88be9260eb9547df6b8bc8874427a20722e8c67be3f641a719e680a82f1b157e21e508e5e0de50774a73fc6e389d19de324a1ca6cf4ce1d1f56961f3cf694ba66d57be02a4eafe5a1b5fbf825e97862a8655f13884f0db13308fdad926fc87248e99492abdb39ba5778aa216390e904e7e3ebfcb7dc514989dd99525906458;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h778e4f5b78a77c7f5db0e86beb00c3f06a8b086813377166eef38e5bec133ac70b4ca18029b7427a06cc5e0c54d674d1cbf25d02692da547ff17a6327fd0e72e265bf0703b337c622adbf40668acb4309b5a87673020f31927a9d3c42af423371677617087e9f038e8e5712307328a712bb9799544d10a51b1687d4823e0317e6cbb2e1d4bd6ca5c76188d506a768cb557fe4c0e92b45859e79061002471360d0d0c94f6838f475c38b3dbc065061fbda2ee0c97e694e9307de84b556e0426cfd38b5c95d1da5e4d253dc1a9bf78adb6f2eb8a64292c4e1e29d06e8cef9d22a27b27aa94009a6e7e95b84cc7e4ec13a9f57d725db2fa24c454446edd6c296d233fd627efa581be76c106e4c5f07697fef7016bc2774ef50c07f6f35aa7ea428a25061389a757c246782bf27c1cf1eaf523d77a458799b698e590cb66172f07fb5ec3aad43b3a294f386f869926e7b5215b0b96165552aa91a6600735cceab3f84c48235cb6be659f934a211469ecd21dd819e7a7fb7ef3669575609c7d0b70b858338c3cd87122174b81443ef047e8b3d04a73bd0bf42a5392315e708cb8ae8d12701dd1fe2089e6651a725f6a2d4fbb4a8cff56c01e20cefe8bdf16164be4cc2a723cd15777c0baeee0823ef758fe62e45b124d4ed7b9b74a8a3d9ff9ef447792cfa9b061f62d0e5d7f92fadd9a6a962d0f21f9a142ba44aee6ad1f9339d8eefe0bdac3b69bb9d9cca40e0e459538c176219158ea995f7c8cb73b8b73b5443ca8ac006f4675e25b7394ad1ce9b3bdb02b8e25c304e6034c31efab5affbe4283161c97c580881b9908672a96841fe0509b08e94fc3914aaa61960528b0b091a5462718a3c6ed6bf574172472ec08c1451d270db39ab312cc3dab28e86b94ae670e0eab64545aa9905bc6f714081dc34bd76622811d1ab9d467b0da25600058e9bbb6ef36672e490f0778bae430f8464b182156a6fed09e178ab8eb419d5c371d20176554ba493adda7de4ebed5772d8e829aba7b44739bc393763b62153c6d5e2fbf0e6676e20ab1c89f8de82517edbd3ea2f9ecd4bbb530311e2ebbe1305b7bdf0259b1aa40ea2f9b214659d53b323a42bd7e7022ecb9cc6ff16a18e0dd6ebf3e6161eb736f86741cab9bc8ca40419534f0c05699818e8b4f1c3e43968a91ab396b1ceef19fa37dd80baceee0cc5c82bd732601e1ada01a523696422cf8d85ee1b3d89ac1b458f8fadffb5ec55127ae7628da9d2031d4f2accc0a0a04dee355e5733d12e732dca229c284b3d78b143993b48d79f092930e6aa24727845da0594f7145765309907f44c9b2499c35d2e8be3d4351eb4ccf6e3c381d2cb67b52770fd51d4faf1062ebdaa25f0e87c9d7a53a26a0e5ccb7f3aca8c5229d2c814890c9f72c5b24064d8b096eb877445aa13e02238d4970dea5216d07ca304697fff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfdaad64baabfce3f62b8a3d018bc0197445a25fb1891260d0ba0fe9a39343a0ae8828a6166fcc81a69bb56999bf1c8934e3055c09c05be86baef4ea55f9a067d73e9617c190f5800df7c6d448fdd00916f07450a0c040de57fdb859260618e9b78fd9cf79656fb1a8dee1f600835524124225050fe0cc976f13c02651a035965c28ad0438288bf5a75a8544ed52f4f3a3aa80966ac065966ab36fb0b60c03a64f3ba107b3b7ff8166474186167278cfb643635d163766399925fe95915f449bf1d093d2356c4e46c59719080f0dd8ebed38ec1bdfc69d8815f9051f2c5ab06671bed2923519c02c142c78784f98bdd286de5494d0d5096187dee643dfb000c5affafc263225a9692d15b4a7f73246a036c6937220ad5f7fc29c546b09f5a4c8a0e7a5a3ec88b0795c03059804c936c3c617122b9a69b5a49156ba1dba80f2e402ba7db71b8633b828f1bb697fd98620db2bead798cccf2794483cc15cbf4e5b8f7a0b9c9882c04cbd1d10a7a548ee28f7b0bb323b452f6ac828958bedbfd1ed3322677c9f27e8bea0cd9b599e1a6b2187f1f7c6f88d6e45e914063c3cbebb2da2a9d66dda1e2e5fb339189f62620a5bab27a748bf90cc89dd25e77803a4de152c2b7ca5f9ac1a0524468626921e84e38c963d71545a891eeb8aaefc0a16fb824cbbfafb12f8029002477ecec470fe2d09b6d7e70801fd142b3c75b37dcb1fc99007592efefbf405000e7259dda5c0977cb67b854a54b1edcb8ff2548fbe910327e7e03a91d1ec35cf886ffd7dbb2c711ef07742ff21c6ad749d5ae0dd86ecf8b40c48f49b90f7444e8bf768e3508fe7880647cbf93bd8a6d2405bf09defc615464d8ba6483ff971d9c57b91e9c75e6a583a8470419f0416cc6ae4cc461857d8b3fb918d1a3e016b395a31c7585112f4bb301cb31c17e3b4490d3ac68a9451ddbb3967f31a8b55eae2766ae092b46b162d4d7b6b2a6034c96f105834df0e16d50c50884add0354208065cc44d3f0da1861a30ea4638cf57af57c6f6a1d97380fac0f00c2665227a52198e8e631967bee03216e10cc57de185c015823f8ee5c737373ed8381388646c8363291b3e9b47c130542da6fa211827433f28598edf0729ee5b4dd1f8c01d8b168c1d3c44e3140133d2bf020cbcc9068612171221db84ad41e1222a7a644d9f99fd02ad82a2a5367c15ff77febf73a554efa983af822b95e94e2ab63c8ac8b4e1fb1375ee424800b65ea0c3c2e11070a2ce4185b8f6594617edb18700aa8f0eeb1783875d92e221f1a0a3a883e0a027306a2938990fdec42d28f38e714f0f99e62f916ac8190ce1251652677faa54c557114ab971c3809902909b70eada8241a16405d5942c0c3e02bd1720f02a5b156f3e59020f2b687b49e20df9b9f1ae997ac1287d26ab7a3db3d91197e0e5349fc58fa02e7dade685;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h18fdf75062afa52473c712febab80bd1de50644186d61c9460426e2f5821aa2a0a57002f5924656b60d63cde9726a44d9cbe43ddbb006cee4ae09201c701ca14a0f845023b895769b5ffbca8b9f54e240f4e7bf4c418f4172f8c14294b8f82c01388d418bb73d20feb113310a0e1a80b2abd8b5e5a1355ea45c2d34ea972fcd16001476c4e110f1f8cacb41a3e63da96089f333ddc488eddac0f1f65ba16c8e26b058a955b1b6581396d2edd6cc20944ba5c85881741348d506b0e58e9a00cadf24173b2577bb03d6820a784550e44c9a192ce9f28cb973915884516a1b8eb16ce9e40825ec0d893d3d09cd7a4270277e1d7fc2693f54aba483e007a9fb243eee3c20aae17c0989b41d0c1e49f537361dd9daad92d639b9e615cf5ab654a631d032ec3fcfc9a7134efd7c67596aee092e2c302b81c1e5f7eaecf5b42132352c94ce6dabeacd14484a6465c82d9f508ac57b12362836b9194845c94c39464a681ebdd7ff4425fab09f25823aace980d65c3883f9b5640a321e997a7fb52a91a48e728e5210b2b93f58eb8c714f0aa65a6e6be535adcf264c2d3a49a1a002ee07ef81bf87c16c02132d13167f7d17d6a4d777cc5211613856ce81f822e7dd34dc18cde2f818002c5be615a9d64f34a96b6e1938fb2db0124e41bc8687e3da35e8686c6b1b892cc55bd07c3b7df8bcd32d2ad3ab53c97fff078e2a68838fea031b966d38b19ed3af8099206d0ae2b85802324d7984d0fef6c439f6e5df6a0305cf45cf4fd34a5291eacb4acac9464b43740b313984988f7abe527779648851027f206f872623c09a693f3d67f9470affdbe6eac210d4f45bd03063b1c487026cf861f9c65dd22e6092d038144bbe5eeb37ae4e8596c611117ba40e5255148523d4a9da34669bc02420d8a4df2a82f1ae3fa43b5ab952db838099fcda5ebc973016af0e1e6cd48d199ea623f71d068fa25d95c265af07a369895c10745016ff1ad8faf3c3c551302ed3bf5ce7599313533f9379d6905f0dc95a15fe378794f5462e79b131b7f2515799566fb7ac614f7f5b4322570e6eb297e1441b56a9f954317dcf27187ef092b9810752d83f73ba8d00c973ec60235bd951bdda5890b0f1e0f08729c99253061f7bf8566738ce96eded959912d614628fe0bb33ee26cac7173b8d0527b241eeda30dc916a20a2fab134cf54f2e05bb43a2fa9996145f4c331c602971ea71e1fdb3550cd748c0df852245fc1f25c9fefa85ebdfea8c2f8347b2ace6de8065df35d357817e0b6296973bf21fa13f60e84a3a4ad7f12b7b81811e6cd22b27b5ca5941361971c782bcd49f97eefb39366af8fdeadb90c39a38466870d864927ff8288cd89fd98cd8cefb2be4e562b9bdffaf4ba74d1a09dc54039556de0505bf2a6ae629f7272edc2fa2508b6b74960072593b06ed6806f1f79797f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfa396bb0c04702ac71d39c4d1b399410192f2f6c72184e2b6c1d7189630c944177db3fac484d74f8054b4e521d82025bd4fb922bc1465c5ac3f995159587ccf0aeda6e6858323217e4e64f00ff884fb3b170f5451650ed4a78ff1f73fc8661597f4d6b6b782dae3fd523b122304b25cd4a177d985a9a15afad40f9bba6f2545206c023d115fa7eb11ebeb0a1ae8081466a107751bca7ddd311a0bc7f7e23d53f60715a3845e76b62ced88a3254a320ea76bb81a7f69b2bc6b088b13599fe39eaa6e5275c2a859028cd4fb58d856093b2f1a1df8d8fe0ce10d133f33102ad6c12481e417d21f60dcd0086062dc5097752afb9aa559aee21d125170a1202ae835962c5f234112fecbc23e95611dba05c74f6f4b10de2f79ca8ec6b4f549102b9bdfe9565cca6d879e6e1ba2d6beebae56534b5cecace02680d4168f2bf25f71fe9bb948c4a89f8012a65c771216f96286a275dd9162720b78746eaf769d4297d81cd3c1a5ae7bcb44178c013c26e3d2e74de58748b89e952e3b115b69ffa55465032308b42159de412895787506b6d2733cc51734431727a6a2ac2e236f00525a050022d823450e0280a7a27c23747c4a058210c8a65a7d9a7140a7330cd10772656c019dae3c78144c140c91a865d56fb08af4e2cd8502bc9af21a43d86287fc5c0f899888f410bdf0da2eed7b444138708a8a48f370de68062a6836fb0191e6c11a6359ddd215bae783416aeaa6b622791ce5a44e36bc6a820364689fc7ecda667a4201eedca4ad6ab72770e8093091b90bfbd8a6531e9a906815cbc702c1362fde9a83ed712112a946c91f76d0fe86813c9119cf2fba7ad2071cbd8e6b9b04bee385d49a10c65388f3a4af1f90c9134e9663588c151640fa7dbc804a7618640a777f531b1980d39a7d4fb1a6dd001c0bbaeff0c98dbe8e268456701f0c99e992dd14ef6174de5277f743faa1f7c12635db2686510d4abcd639238432b50741183a50e50fbceb4e59cd06ba564561717b1f1bc8ef3dc369e42ca25e8a1532e50b86dc2f9b690be95ae7b6c0495415473e87c361bb678efb4646d5410220b40401a8041dbd8c04be760d1d4e860ca3e9904688d169673af4bb88364127a70e58c3707b62ce9bbb620a58d319eead5034fc616057b956cc2c42374d31ff2bf527fe3b0778415669e9b8384a264f92782ea915fef8e18032f1311e7038b2598f3b8e27126e57cf879118328ae0ed7e73468076c4ca8e2409a77a7c963839e43e71833182b5635b0fd6df7664ce8143f7d0c7bf2d815a718d8ac253665014e7cf0aececeba4ec41b17ba1987f1c15e5ab5de251daca388ec69050c516e6b4f5b188ddf5ea90b150700fa346362792e6b300e70ed6428d8a06359b3ff49f1039b1cd5bd2d410bb167d8f4eede243a3d8b754f4686608afc80687fa98c83b1d4656d3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9b945ea26717a94592041ecae5aa15b8f920a964f01519892e8e7a3e4c5a56e8d946d4cec7bf263289dbfa34ef766d1eee6074f80916f2aa1ea4370306602485cdd96539e1a0f46a66c3ac392f4a1b6fd6b5967bc986ec236ba6a7d954eea03bae3b7e47fbb32241530d487ce47e74d4ebd5c984c69d3b869f04e9d9f1ecea46d810cacd98f6c0286c60fc699aa48f770bf06922a2d3d489913eb6a65eeb26efa216e2728af5078eb3adac45e65766aec64b645c5d15bda46fbc35bc2b8ce68998e6c0dbe480a884ab2d9982af1f533a55d28d656dbf066fc132cbea8dfaeac490026448e229c11aeac64cb5f0971335993e790569aba792e39f9d70006c161c0df7cf5af03026cbeead3c997bdcc77edc25433565cbab6ff798dd14b5c14ac4073601f950c5d2665961a52ae16dcee71289f3c1a007e91438c43be4a9f62be36f02bd51f0bc29fb5b0f44dc709b8b46a67cac124fba97e0bba75ac8a14cc9dce66741be57e99d1bebe697c5196801a34c6af189f3858acce3ece0edf1684177d7581cf6139008f6427ddbdc9191cba2696e1d5f8b8f3024df0fdaa3f86297d1403d637cec49505e7a2e3f13a603bcaae34db2dfa293cde2ea4a67198fbc59ddad96d0f727174564727ce12130052cd6d0a7cb3292f9f92e02fe9105adae9555511f7bb7ea5b4bb2c18d80100396b5ed5c8cd54a4098a392ee21d18c2f20d740de19c21f6738c9029c3b124caae61cc48c22ecfeffb9ec1b351d5d535bd7374e28337f4d0514c1de5dc70d89a86d530d8632b62f860e2cecb79db8c1193856788b8ae8bd8ff8817984265e8f84c6b428adf06c238de8baca4986acf0da76bf6242c7e32713333dbe1dfb73e59a8125d1536be4d373da481fdec967df7f5020441790d5bb8b1df630e700b2cc9921d1a65ccf6425803bdfe0f54b522633998d449ee4cd8e018e8550d80d7216ed1ed37106579f56cc1af9df19420fd62190834ec11fab5a12eb815ba1a3d1e4d00ab708d706144b7a4ebb69e01f6adf01fe7cd24c1c3b743e862b760e5da927835f9d389d40af122313958287fb151874fc0fb4d6793d96269e5630ecc872cb57ea66fafe8d41e2d68c25532dd4c67969106da5350ad3405c54e93ee46122e26d1174cc18d765c294027061ff5858b1756259260973d9232f465234909d7e1bafb518f8428d117126f28c03c33f83f799f760bb17afe3cf32422500f1831fbd33f377021552eed834e420fd98df8f9550dc177d7e84cc76dd9cd2420bac1ee11f117b2d71ce9b6a2adc0a4d9480174722440e27f2cf351a71265a2b9ec6e58c99419f6193bf7cc11684c3049ec29d610b042d2f1d8f19daf666e2b15a3569826435ca232a20fae979872a5deabb9aa0bf4e03f61d6900c0ec2c2f256e5169061a70b0ec2b0b102d0b31fe261f54de6ca7918b47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6fb50861fe16daa90a3448721c8d70f87d1c9b7eecdb8410861f581f25828af9439594aca7714ffdc579475c808a8470b6ca026d099aca1c47defcb125aa88704baaac4d27c910ae2dfd82436beb19af481fc4f5aff390ef3fe2341163c00920cc2e17bd543da1e95dc78acbe6b063ad7e7e2b4ef79872a345dee53c41c4853ebdfb24c32c746c09eb1d469db35dc0c1ab81847c84c4417ba297f3add1da046a49c5b53ac1eb87a5b93384702213cf45a6c2365d5539a1a7a7ff0f3deb44491ebfe2470ca1b29a9c175cd37784f5277fe623bc2d620c06b266e1533d764a0a7bf639d98b1e4fb7d20cd42fe99a646755205196d3f2f2fca80362b6a6e33b988f40cd75a299ee9572b6980fa3e1d4102b7d524d336fcb85b2ef2623596fe3e2168029e3f4be4f7a4a2f77aac981a51c91f836003f442d769972f512a6509f7aa6a93f39968f00046a3101b80e069e5f1372679d5b278977fb1d45cdab601ddd9e771a14a260e51b0bcdceaec59e66984dc1985be0801dbbd91f4493d4d1ef646b38d91b63a2a70fb9cc4bd49e6b8679c0309d7f48ad10f119a8fd5b36986dee5b9b697e7dce5d3dbeeaf065eeb0f05b420546c0e48b10938a2579430dff57910452fd4c68d2494c42aeceed9fbf10226f1c7c28dc8a75c0ec27d8ae3e9d727465f2222b34639504ce0d8bee8b8c07871cc6dd6b22586276f6611d648ecc9373372960b570dd2723f47fc625a9b095eb57ba3fe0168ca21f2a11e051b3c9f30ab7f2983d13de6e644ede7b256f01dec4639692ab58a0cc2e49148883938c89912cb9711a8624f19ca4b5b64afb692cfcd88ab754087db7e004b84aadbe42054803a1c1655079a38b76e1e96ed46744cca47a97a44521e9aa0ebf2e3dd2f6b256740efb80363d18fab732099c08a57b9f6a5b95119ec285f29e10c4662c564b0c28dfc6f08c0f9dee577e5b8cda5d44fc4bd417367fe803bf2caaf33a56f33a5f66daa29be030842db51897e58614ed0eb5d8f6a1dca478ccc62571e0cd5328414b7153de2cbc893ce7d2c4bd73338365dbd27f19a96afa69aae77001082d23e0971cef62736cec7fe523f450a02a6bbffe281afb400b4e9b3c349e11ff4666f55f02ccec1422733b1769f4cf0978edbbb781995cdd50d7f1c745d5886ea4730bf5013b75dfdf2a3abc54c71599fe52725e8d6e8581f5297d1507929e225d7123c5cbae274ae99970c3943bd3a22f8a505325b3a8fe171bfe2cfcaa89a92786fc9a1dcbf6b868c7d0fef4b7fe1701cabec82e579e0e677effddc17f4e75d176927194401383f8f23f5355e9c46d46fb351331d91adbf7e756d022fa7cf12c3494d5deb4295f0ae258e84759e9e94deb3be7d9e9626cda8328d5eeb56e4b9e593dbb63285a765b008eec676f72ddc25b0c8b4b24c72a62c32064f0ab7d1a5006bc95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4fcd2a356caa848e85b0941773a305041acbb038e1b42f6255b3df54ba1174deefe776ce66202e8a71b47e63d1523b520c7505523808942432fc8efcce0a53953099c6f01a84c155996b834e715eb6e1414231e98df7e39f9e2879dc6b14ad1a3316c4426b70bedefd65072f0b04115ec346c994e76ef48ec18b31b0c93e86bcfce96592d3e4fc426f1bda1c75dbb6cdd9eed27de2ebbbf173ddc910e5bf6bfac59313c97ec45e6ccf7a734bb82ba345ff6612e55abe12c8ceb86dad860ea913d5ec46963e16493e951338623ba91ddb0beef75f173b74549b73e81a25cb768a8c3001dd3d689a0fe1242f8447409f5b81c5e5831d4a7a725340dc826ed204e367527a9297055609f9f5728ba1e20b06caa112c395f87080b96b078bd3cc3a59506154db892ca9d9ab2b41ac5b6f3c6b60463357c7b3f2e5038a2121c7e4e278169f1eacfd9fc6079e8a74e1c8cf0d17d7b6b39097a53dd261a44b05b768f45c3196c380bebfa41ae8067181b65be06af5a80f540c54a77e97651a452bd2f673e1bf73f6af7af3d92f3ec3085a972387ce5370580d49ab25f9c108a644cf11a20c8606f4d73b12ff65a57ba4a9c0fe992e6b221cd73d2125b4d3ec8936be06b0feddfe7fdaffedff67e1b6cc53dd67f2673b5f7bba4bcd5b69d46dee0cd053df23967316877d7545238af33393940fbd9cffd51967e22afeac5d152db6b03a8da47869defbeeb7eeb3a6c003909b1020896d17009be7200cd0ed90f1ca0d48e4bf20c5772e787035955ccd093d557cd2f8a9d52dad9249074f275de107e0182d49f4caabf5f817dc6a14483ba2eedb2d9b64197fe32367bdc8cbb8dcdc35bf74c7e54d42674785881f5f247c3e173c93931df4edf4ebeb3c90f437c77b5d90cda46543948b4ff925fc9a4f3f6115c4d32af6efceec713697ac8993326db7f181a755c11a07ed4f434cc8326f953c28549d32276345d6666bd7a59510a69598847326266923fc96e6474b7ba9c381dd37112b7e14212020c452ebe58eed0e09c42fe4dbc6da097bd65e797f7054b5ffe71ef481a2df43a785ddc15921bdc8d5d5d4f1cfd465ba1b23455246afc4a1344c96965d964c0b09977dabd05c1cb8df078fcc1503094f0691d4c9fab20cd1b2dfd97e0ee67edd127ecd0efcc1edb650c248710f08d2a161e12f194362910596df3a783d301c2082e97f1398ae56dab0d4d67893c4b5d74ee12e9006abdf0229873f693629b3712c76b018466642f9baada6318a23acc5e6aa9901411621dc23cb3a7d5b31176f422043395394531e705635ac6f9b62e8274a7f56b792ae08b13d6962d310e262875cd26ac2e1057faa4bb40d48f7106e662bdb9116568d19b6e4a8325b25784ea300b87c7deac228a0df6b26c8e18d400e9e4af741314358a4d6fa8b6c609c5e553ffd90f558621dfff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb13bce30595b71be67c405744acc49009b8c7f6a623d5b418210854f3979b258f06b6820dad4f3fafb4fbe8fa73ee669633aee8e7b300deb8be267d28fac4d496bfa210f1949ecac4c56d9e5a09403c909b888c3764146f20282132e581cba1ba5eb16dad4c55e5c45d3e0402f36feb162cf61696ba7f551f4d0e56936fee5a769daf4ad66d1adb0a6a0029e01b57531ccde7ccf5eb4a8e89e6c121917285f028e90f3050df542a0ff4975571bddcfe075b9dce0f72733d382b488a89281becb132222bab88e11c8944a31a70078aea416e69f03a8e8a963ecbbcb81bbb9592cabb6e23f02136f046a76fa59d8f4314724bdb888a05cebefe2e77ad8ea6ce5cc15bf56f7e01259e1786fbc184a899ac6e3aaba008f6397260bf1bb02a0ae5effdbb1b3d9ff9d44aa88f38c7cffb35bdd097d4c56ee1d583a6627224c11b06eb794b288e145d81d0eeeb691c7518618da038c1bb046eab2c4fdea54b36aa3d0360380df66345c831fa4fa410f63f99935a475966d65bdd9a35551801530c5948300ee1b4695b986de2bcb0a12eef9399495b86998d9cf275fac8438b341396a7eca74a5c0e3ca2f182fd0f508b22c2bf054a56906d06f8617c37046da3c734baa0534848b05956d19553b01eb20fe0de6ff28544d8375f8dd7f8727a8a38237887a7aa328332409fb9a1003cf69d97459fa46117283c3b88c9bebf368cda3eedb6aa98a6be7edc7f035ed1f8e6bcaadc67870bcdd7e3ff699182907d36d8b19c8bcad2b43f64f5065e7073c5843e46815c8a01efdb81c5008913981d93b66d34dfce09d7c66a5dc090e036590bd9ca48a49e9448ce5773fc504c3b779c0451275541515adb0bff489f16e2fb533330e707da8d3a486db8f94ce34ed49ef17adfdd0b020cd19ad14df0d8af714ba8f5ac14d8f7af535430758ea2badbfff8750b18e09fbb743450fe954d1c630030d6e0d37878f91d7a606ce673517545b0db52980ad8e613ae19b63fbb103f3e4a10bb8a4d66d054a7bd9dad0310c23b3adaea50e2a23fe3b44b80ca55f809856b1548b199dd43d4a1a8d0130ef63c4b5257356600bfdb54f8db01ee6a0f81e178b90540e0158325e09d11d42d3096881db9a75355408d28c43fc992f989fe61a47eb1da6d059b010feb74db8f8abb3e32484ce7f1f6fc3dd6bbdc499d91e258ba8054b66eb95681e97e549ed3c8347ca0dbff9578f8b9eaf04aa4d52c268991059652d081249d704d0a17b0bc6499cd1b72635fc1fd0a8c9a71c3f19da2771b8a2e5c8d9e14b2747a4027763150c0d3374f2cb09a72af02907821310e4d706f7f753ad80417c13a57a53b45820f9cb5c11ddf39956e29cd249dfd46f34cfb514367412f188dffe5bba5330d0cb3c91ff81d54006711072335f595d0f8054bbdd33f76675ce2646ec8cc39f82457582bb7ecd70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbecada2b7b3a9c73b606e702de468decc5a4d629127db40569e60a879c5124833a1a0e3aa6200f062e8fcb0679670d39994be70f96e8af86b4dc0abf7270d135b6a579209149dbfc1161d74dc753aea7c7ae391d727b04413ce32bbf97e7babe0b03854437959ac67f4a006b41076f1a1db126a7afd082f5ec52f9bf2095dddca67660c21dc0857bcd81f82e9b564dd4aafaa5e9ddfe8c65214784fe6a7c4de4832e2ce5d8239679182845c9dd608213517eed9e37b5539bae0eddaa33a94e151f53d19402412b6a397a7ec305ca4344b510d09c8bc8372e7fdbc0f2a6c0137f8f99a7f7cacd11066a43f19dcf21857ff3358225c2386f9540e514ca626fe157601f2f8092c94b296eb4bd5cee5200cd89766c266f511f8fe83c37c9f460b51e776fab5315bcff31a2ebcca08c05b61315fc2b19df369e2879b36b01cbf19f677da1721f5928758b04c563975d2bad0deba0ce1cee5370600054cb6c28405bd8761ce1d71b42985a9315fe6a09de02b15701edce574b6fb0490b589c039c1b4eac098d26a3e5f6e1b72332ff9b119fdbebe1ccac6e8e85b240a60181973718d496dd9a586f04ec4b5e3950652a8a48244d85b7f810f0d88f5fe6108f5fe4198e29e53a96f55dd73fe013ea47b7151526842fa3a77974f6b9094fe901e6eecad7eaac176519c2b5a8af5a8a8bac64784bc3167af2761605750841c4316e45916bd9675e4724993d7fc7058e2f7e9f932d0ce5457ad3b7f1183befd8c22a4fc270da9b36bb799543089092bc80dfe6e5e481276021832d5ba8199bc14924f5af9e00367af02be54af86f5fb2abbb4154cb232eb82d5b10ad74251c56de8b7966e5e903d88f84d8c8b2d6960100d758b2f8e8532d2d2320cf6fa36a83740ab7c8035d9cb9f68ae5b9af13057aa7a890fc3a94e0ac25bdee38249b93afa336876ea9101cfd48c2a8c9fdb2e0df5547c531f44b553814291788bd7c22bd1826077c6c063e5bab9cc4aa57bf540da02b35d20bbd8fe3ee4943af1969a3a2917e556097a31104caf5d7f0ed4c828bec216b7a969372ff118ffe5147a080caf878a0df8d206558bddcde03baab4958864e06e84ce4362958072bda020ac8da7eb41333efcca4c7cd26162284e513e2f0353919bbfa0539f75b04e1b6ab297024f539dc3e53c98fc9d22be1f5efba80e07a2dd19cffd6c6056b6d66d28443df4db42e0bddac3a81b015276603d9e4a684a1f52a533bbf1370faa5de4417b53daee2175170441038461b869c71fc8b96f8031581327155fb6cd3b8c53c5a8747d22261b74b54317f66b4448277a505196a65e55ddb0a60edea63aa0748da9b10903a458c617d6c50b055e84da1fa655e21b489e37a56794701368fcdc68a46b1adb3e54807f090eb557fda6198149e53c3a7827adaf83618416fc4d152a01c50c9b98b7bbd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd6b5936419b1839e43533c54b261265acb7354bc43d3e082ca0e2acaec11a8b06274cb27f3ed7f42ab06f4616ec14b1526404df6bc3046d5ffabe7560f4a910acdec2b0f6d50f01a24b3aa4abdb26f9589c81361995e1c18584ed844b619fdb9ea265edb052a19ceaf35f9111d5b9868983ce951edc487afcfddc1a2f10537abe5273a0a8b907eaebd64a6c7586838386955b04d4e38825e4547bb27064ad05d3d50ad9ca1f5e1cda0f8f42adce533a455d4edd497f0e993081d9d8ad1c386ed6694d8f025fa82f12b3452f51f82c931ad163e30a71e7c7401746b700ea1cfe7e9d2bc8bc1c20a73b998d12e49261f3422b724606424b8288db0466a0b17aa93608f09d5f2064c78b49981f72ad74f715741c3a0d406a90e0159ba5c4f75d9963c73e897088de077fb3823940362ffc837ec77e0dd04e26e8af2a65e9d68daed6dd2c1c26bd8803cc1d64c73c4c4489fddc5dc0b90931b2fcb6e51896f21ff2341649a975a0bf6f6428a5369cf9f0dee5f0aadba1ea9d843b7add485d132d733e9cb1a2bbba213e9a34c43a0dcfeef1ffdb2197510ea96541fdf72dd8ad9f79bc0e25253ca347ee6f84ba0fe4e07ac8646963ada089b5406eb0fccca7aeda8f4c186ae409898200005336e05f69f4e12534b8b99e0387a8ff8ddae8e68e61ff5a5ba662eab74e2bc00202056f35ef7e782615ba3d16ad2168c2adf5a0bfec450f0b06ac5eecf1871ecf7fe05d289be317e11ca31b49e6c85e95be5168bf84767d97a5b77b457a7592d280557a876862a63f78f6033390c54b7c94baef1460d8fea4f3eda127529d0afef484f9480c7ea8ea72eb6b46766418fe44f524de31d8a90af1f63d3490edb1db14a77ec54fb60d61a435e5f138133d27efb73df9072c0570ca545277485bb52471e46f12d68bf4ec765e0602e33b0e4a470d52474abfcd70fd555a8cbf2c7be865f9c04410304575cef343e4c59d7ad91c8aab655fc8127c07b260def6fd9f5ec56c085035514cc6791114d76dd8190b1d0dead327b08c292b3fe6886e7a1c186bea8ed44ed772eb769fae87d84d9f7629306f08e19b3625c3a812135f03cf19e8743f5e61b903dbb63a25f7d395bda4c9ee0e6a7e8a76a6febd5bf32a1bd8e304239f90517ea903b7a190118c55b264d7a0ee24ca3d678025ebb479033cf90d0d888fad8972a71a2196c3680440b39b36361d68f24a5f4bfeacc8fc1917c3a3c548224210dcb5e2d29cd7fe3e22b024e43354f7e65738b2e532b5ef792789de49fca499bd636b11822c64e61d0aa98657825b4e7a66d13a5f837bb79676f4008bea93652461517b4e77dc05f1b48ace41cfb8f354a471a204abf7a526e48fa06a482ec59131aaf500bca645896c49aded7c1e60f73b54b8f8edbb4d305a63d234c96aa60f170dc79e8c6e6c017dd4b1cfdfe99f53ed5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h76ee37f1db40108480a06e5f41920819d482324e2db4ed4ecd7ffadb2805522e77dd45c26a894e8ee288703d5b629e291401f9fda74068e920acf2554b676d2db5cd067ec1b211bc05c008fbbedebd0aee80bd510d31e6714fd5e88986fee528b3a5e724b50dab66559397825790ac97c421a38c8e37a1963ad64f9e758712cad354eebc39c6a1471bc3cee49bc3f2481873cd80ed8f36e7fb58cb535fe197c6e1fc25ba5761b9a669413bbddf0e8acaea9c902774c3d0dfc8744e1147b8a0e41a3c90c8949cd53d98e8f07941044f295f7d508802b93ad4f556831dd1aad25dc9fd196444adc2ef801ed86cd37b3d1086815df1054fdcd444910ae9352a11915f93c57b66040d5c422126be7135dc6b702952a4925fa0c544f52c976dd6c46a590101c26fe451e490473db58b464491eb2281f2d19e4e95a291eac13d2ebf194f0789406a07b633248bbcc4e1165b7c4f9efe1d25860d98f5e926a15b947d0365630603e27c375c719e48e4938956a3a132c70a464436dcf96ea3474f5932210d1cbbb1e80d48278fb5a239880702ee64218cf14fab2aef4686d0932c26e1eca1658b8443f5657969983655d58dd006314f6e0da73ac758e75ccc071d5a95f35a62f90277118c3860bd19d907f20370c0fcfa6ab3685bdc9280a2c48620eaf65bb47cdb9546612e1f6d2d7ba44ebe5020db68c67a35e86027ea105a25f6e1fde8e400fc49c7ae6b84fce8073519266a046ff5a2948efc61a667da443d25eea65b4243b7012a6e5578bfc2a1762642d10bd6d2eafea58dbfe02a3b92e50bd056622ce18dc6cd1dac612f67b6efc33fbaa2b353d086f6686f44f4eeb5a977570bd3ca370c703c2bf2bc6f61dfc3b0c7e2bc0d2b443f002ee1266eb66095630263c9f762abcbd2f079ce4795e0bbb441dbf43148480788276575e7fc9a9297c8d9d40002e61bac33734ff0c2abf8a655997c4e0ec4316b4b9c75445a844338f6eed05f978680cd237091c995b10a39ff6acd87dbec167b6aa9b483770608ffb8bfcfac99d27945c7294572a8134261d1126cb50e1f89aa5e7f7560dcffbabc88acca6214ef8e3f10893df7ff31368f9aa7df2a505f7bb580382a900275526c35bc40086ad3ea90475e490246216f47413210f6d4f20289d86540d5236cf03a8637996caa94d2510b8d9fe6ce0177558ba61d5f29a69c288443a0c4e45395ae644e366c4de681b840a520da1d02432eeb8e4045458bd7b8ad98404a11c0825b56eeeb238f5f9261da8a4e7469ee50cba8bb95db467eac039baef7645444905c4685837ad3588d1c075f47a883482e18967fb5e2e184d3a815238a4c53f6088e11eb1bb4d29fd2af388619c893997efbc6c8639eaff8864bdb9888f91786ae3e204c356e6c35d5d85afd305187cf9de62066ee6bfe0bac2393a88d4aa98733cc5cbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha9f0c9525de544c7486378d59256e75fe3c5de7235ea0eebf71622db5f4623ba3eeaeb42d5d3713927e2892fe9cac764e4554a94a8f43b58fb8bfca646b241cdf02f488cd7187dc5e480d490186454c55eade9a4c1e8d2bb32507042ba3cbb4af60b2b936921b1e8af48c5809ddeed7458b455142de33e7d40bd94f770a161bbf2d7034661f4736788d44834c60b65c5cbc9c9d9c05fb4e28242ec090e0db4e0132dbdf843eaa69e8191b229b00a75d62f859992b7f990474aca64c5d784ce147084c31110fd5d3d7351f1b7c17979e9c20c944c653a4d727c8996dc57ea1cb724fd078d8cedc3b66f84151c96e2a721372cbdda4adedd0bf9eeb5518432eb8b376b2aa5d2d5b523dcfb8461ae022aef1fd2b9e91a69ffb937e8bf15576dbde82aeaac70ef8d955aa29cbb053e6ed759d2b55661806e137cd7781443ae9d8a1f5612f86d82f5c873a011ccd2d44dceabf7ea43ca3d5128b80b31f7aa98db7294df04aca192bc90d1032bd59c2a1eab6ed6be551a5a0777c0a2ecf378b9d6b063c917d6f4a6b9c04fc7ab96ef2fa2a32716f2d48a85267841f6edcebef3bc3570d3e294006f14aa4321a47a50c019f9c5ea6000bb753ba15ac577397d3bcdf9abaaa4356651d83f1c3280f30cb92ebf0b498c4f531f203cb7591aff356dca33f14c4d3fc09ca4f77681e65f95ced9df1453e4617d0988a9492787d497d244c6b424dabdc4790555cfcad17308d3f40623ae0ae7de53d793d10d42358bf18789234c75d90ec38825f56a08050ef9ccc7b0885cb24792b1b72f49cf3d541dbcd8363f59f51f595a0f0637a3b6a0cae44879ec3746a49be114a00aae524dffdaaf2336ff607565dfc397071935538dfd156c0da2807894a9d7193034ee097a23e4687ac0eeacfbb3eb5d1aac33ce3eacc417b727bff4f996856af393cda03893d53356209ab1717d160637a79b8009999314467af8571d9a975f874555d60d1b30e99a2a3a58bab57b23191fd321e67e6fa2ed7feabc0460623c74b407bb85c9d837c23da038538069289858e379c8f6232f0a1ed6c8671496b5356b9a1f2cdc5a6a580ff59f5c7853470fc505fa7c4288bac83c21e7a31ec073c50a99d11cd57b53fd0df497355972d1cd0e880791a5d89bcbf3b5370c12d340ea3d8f42e6656f7e1d6fdbc31af623c09d444400e56a9534248da4661a4a73b0a20ad68733a7a9a3d6436ab36237021dad1aa5a33295952031001b5e2b0fdcc7be49c4d6cd3cf8ef74205f2a2be10a10ac3ebd37bb2d6ef50e5d5e24a164a873f22f9811efc0d7e003f1c48925ece2ff708642660cc6c6c9532e41d3bb20ddf93e12507bc552cbec2fa11f22a09ac3fa175b51a3a1bceb873c24f86b0b3950a0ad0c4aab4e3a0ce02db0927830cd642563212a97f33bb7c73036180d291747d2237e49415b3c81d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdcb36a6a20440ec4023721323d2d656298ae73be9604b2184b769158c4dbdb582fa11b54fb78c807cad4009228e4865d38d96216f414cfc918485b67db5949933d04fe1bc613fc3c96192c355bcedadd7afa0a33d524ca234c3c5c642de5ac4c103de840407980e44f3ac5ef8029922ecfe5ce261a1fb72681c57077acfcc6910de2744f3e609ad6165913c8442c95089a835fd71ec3211689bce2191d38328e8eed763bb79204e18bda5d2fd55a67a0ca025610e05f5b46109dbd255e17864648d88524779f6df259cfeffce16e39994c44e2bdf26101eeff24013a8dc90f393f1810068552b9dbadf3a76d8a2a3411d90aff38b0eab482b6c141ea7b0162ced9033a0626f15ea4fdae7855fd5872a4ace6c85146bda14b8669a182aab9a59cc34439e1c03401fa4f7dada5318974a78764062221d78b1815c0b04430a0aaab0d784ddb04f3b045b4af206c4767e98fcbb9e68b176437e16512450c2cd68483ff16652bc1095b61fab618160567c2b1cced12314cafb422312c3c381e1e5427fa60134429d2eddeadb1c8075b7cf79226bb6b9c91be1ffc603c3254fa3ecf0ca6ea325ebb4fce69c22b6f7baf5a7d4eaa040c8b106d7a784556b951aa4ba2d7a169ce1f242aed0544a055af74b09a6cbe31689bb413ee0e98faa63d6e12e2bbf44fef18afd9c14652003724c458ebb02c6a3d9a6dca79af351af5671a09fbe14445c3bd3afee02f143bb56d4f5527cdbbbecac7bdcb22c38ffd389ea21ff21d0d469fb30d44c29287111df008afcd72bbc8b2ed3bdafdb552cea29fa2b25e9862545b52e4e9250e73062259b9c8b18a3e134edb0dd462cbef8ccb5bf9c43f4d44338c9bcbbf70eaaa83e6a3231b19a89c6dec2ec61f20ee95f1aa4e4def218229743eebc8db59eed982979f61ea6fb846880193f7d2bc7796f77185c97b9d9491a078e931f157bd21c786537cfe5bb8601ca7e64c8d2b22d7f56c53e7c554d19cca4a4e6db01bd995834684a7d5456570fe34351f6997cef483d2625105ad71b7d4f0ad66b1bc860a4b17c9a2e49a41771bbef8a0790e60d77c531c56862f2687b6e8f834f646f17faa295d11011a927c12226c64085b4bb61393cfa3238b2ea273b4a00296f30c1ccfa623a237ef921d135f925842d34c42cfa61852c760d937dec6f43810887ccdcbf180eb2821ec7a6610790700be87a6d099bcb531bc08321a95617bda8dc80b243b37144bdce81284d4fd452fa6e1e285b4fb2236c45a0b7e4f179e06ce92ba3343c1131a38f5a7a8ea33d78e87ddb822fd33b075bf69706a69a83fa49c96888f56fac8556620168fdd81f72c9e3ce1dabcf64fe27b62a96c6a60422fb1ff76bd55cdf782ad34aadfa7ad0d504c8cb0628eefc313bd974900426e824de1295bb32b305137d2fad63e281d8d4878332d14c6f63b8ddc3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcfd3ebe608fb635a594db8532704bc5526cbdbaac7f3c6819bf7042b7b93db3e60774bb1250793c4487b3ed8d80a29ee1defa986518e280c85a2fe232937520582db45b3c97e5187ed16414b1736dbbb524b70bd20c4c2c828cd886bcdb86f7fd2d0bb7c6d8fd0c6b2559a5c52b8405dc37bb13b305ec93273b053434e10ac8bbd1897805f2282f54dfd0d45b1f3b11cf00fa6bc09901cb0a114fe2fc7c43bbef81de4061e61f57b31f7b8c62d5aa2f2df9858273d41ccea25965df597e24abbd8882ff480f5299d398e359601e769bb3c09df44377fae359a2531e1aea512a1f47307232efc8881b1174587eb0536ec84ed754073d71307ba9a749f3262b515e47c8ea1abe04221803f2099900302aaf308544ec16195bd5f10a0654d70ccdcd9f576aa3c6544ce1c5014f3cd6f396263250920866038fa15c7239e73ba1202b62ab9b977c5a238160c4fabfcf87028784e144b5592ff5724df084597ee99473033333f925e88c632a0293b1c601ddbf381de5418a19d75c3b3af3dd823b8fc3f2b1a5d20a0339cd07e2cd217fd69700d4c71736fd4c4d25cb06640d11369e4224a956a3bcc04703dd3525b410113d5cffb3e00eef07ee8ce64152429070f13f0f7c1115479a3c0991d28ea5fca5aa8b0b431449690777c13070e6235533109e55573d1c74264c72159cf1aebfee3048d7f625e0c9170efc13909c1aa5912d3569c0b7f94ad475044abc9af69b58376d8265cd33a09d6afbc5873e1c93778b58ee4f2a31c1ae7e069df933b53a0072f0f310556aeb688dc878b9931a6dae5e664fd2cf48921a4ee198f35f1113bdf3ebd9c520f39a6fbf7447dddc512c3e240a9a7d576916e10f2cc76a391592d0b91ddb56cd60abad367daa52d836cc5922c721ca807650b7cc100c140404a37ebac144387f0c05669db3dfc9fce51f06a8d2bfd1198d7d9ecf6f32d85dcbc633584cfdc5d9120667bed4dd473d27527e4d94c30156c6b6bfe486e937c18ec90f9639b6dec60569bbf7c32de9fcb894a965fe5bad0919347b3eb62fd6fe38ca9e1034ee26d13c39b4e67b509f2ba8b35fa26a260b12f6cdd34acd8e8f1b5a3a12f7e4298e355e5971b22df73f50f7de79b5f6400dcb630dd1fc8eff526ebb86291cce839868f3ff2ad32292be784fa1cc3dafc829e0dcf24e2e3e149304404bb5bd6f1ba1de89bc12f0e234b0c34c73d8d79a580a3f22c7cbe8f8ed347557f3bacd704c6f4fab8cbbf1a98cf5a92183ed66a1d0ccd265d22bbdd9062cdf4465a2004cb405b8db4e31bb7a7dba616303ca462b4adbdeac9161f8ecb217a4f8095d87d35fd684e696a3648fe0f14635fcb492c1c011274ad8b30bf7bf542d9a443bade2845d5f9a5ca6b6baec520952668dec83aefae20907c25c4a94bcbcd7a02b42be1ff27a7d5c245d01d82e86292936f1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd813313e76ff3fde1d72f1520e9753f784967f15cc84563a004e3f53a9e57fe42728e6759a76411644f113511a2ae38be20ce713c722ad45637dbdfdb392712d14580e36e91ca41f9c957bdb361e082a01f761b6c5bea9d61ef2a8aa8a194284fceab0e932c6520a0e8ae8d414eccc1a3c9d856b4f32a0c1a9cec71a62f73f40df802b056e8bc77efd849063d3ad2875af782370c2900a3bf1d9f24be8220ca200799c0e42de83f2f8362e44ae4a6b19792c19e5328319aa8369650d99b7cbae58f63f2aa643743c363944f67020a2385b6584d190bf0165a3d1f388fb391a903a223998fb29453a986f205c96194f109805697edb3c96f564a6b23a2b9ff2969c4d6eeb690178b2bf557797bd37c9fc3da7b242cdc7a2fd04476023ce9d1bfb00c8b99c22e371907228c126a9b8e00f736331a55c471fd440eb809709cf81dfeea387e9a9d68ddd994610d28ec5567234225fe23ac85419255c4ebd1b661490587d834df0bf2e9dee64a591b74550216cea62d1b114ed6ef84b37f6da63e39bce0cb2ab56291f4cbac85e38bcc8a6ef25b1521e17aebe8be59b7b3be7f0117b30a990489431cfea7e3d08e33f32574ea0c1fcf5564bb41dc25a8aba28e3b23af46085150b7a16372176466cbcd66d01001d050f39d494e53d6e114424cdc65afc66c18daddef91d3e8d039b2b2bd2fc2f69bcda5ebd28aaeacdfd0848917dd59e4db946eedd836323678c524577534e791582e2680c466bd28501192477d2f7aa09c91a5991bab5e548704c03c66c9eae72e9126980c0181bc9f64f05cfdf1d392d38d839c917d8385b3a1c1d29ad5b5d7b418fe8d243573f8610ea624777c9802df4f83781088c2f17d8cd9aca7cb5fcd7d75c12054978581452b35bb9b5157ccfb8e083cc642cf7ea5f31b30d4f5e0001efa42c04b0ccb6d863bb500e751d111fa57b793167959ce94470fb789ae95096dcb45ad88be2e17a62f80d9cc8edd1cebc39e889497a33c3fbdece83be962451a7a0fb592bc8a927627bc919f05e69a163dddae20f4f0a4b18869404ab333536b7498f24153565b273cb6baf1d49bf8df3b2155b570fa38b7cabc8bec1dcb7d66b071b6d36eb992f53c18389769d168b665a4949be40bcf317ba0fd14b02ca9092b053a1f6d37853d2ada0931e1d87da13edfebc6d61d50320bcdcacffd08005bbaa15370337b32a08f54cfa03f84fbdd2bac90879ed8761192a80434ffa38aae6b3878bd9eabd26bfbeacdf2ea8271129bcfda0a547cced62c82afa9101bfbac7d1748eae5042c124eef908e8bcc0fc7981603105efd9d4c83f130f1fabae912f0f47095e22ccc625b9d2e39ba7197c6901fe7873ffa7531313ac03297636a0d92716db4062ae6506783d4602f5696181c3cb46134a55e33adbb2c574ab807956b83ae41c6e5f85c3cbe7b22ab0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h535870803f5431290df308b3e6762a6b00a3e4748fd19f03f9760941b355e1e623806edf957ecda5b3770e252229e1a840ed0b29efe2726301fc507d20bff547fb1403a99067abed749cebab5b94ad107feeb2e919a62b34b5cc003b32f8a366246633c21dbfea9f56b80461f60c50e748c469f868dc456985cf84b4fe571f4d130e10eba96699394aa7cee179053c1d46437965b9721938150018d3331d95eff6d9eed4c5f9305893bdee231c71963a08cbe1077913a6b0b1012360380bf18d1d6d58b1db779d3e036af5891b7735a12e099d3296030bcbdc57e0bd5dbf8816c6b79ba3326a6fb097a030ae123f3083759d8196ccf57653f27b522fae6cc5ca8c32f72b66d82fb8980faa30f8a4864fada7e894bfd28c4b4a5b8d442d266652ae5afd9a021605bc770e1628c37438cc3209d5168f25c4a7b2bb4982645ae0a8295964a25d2e3091f44e899df8f80f12a785a723b64db5a06a561ff14aa395b83f4473fc1c81a03233c5c03e3ea6d82dd71b20ca8c4642aadf5d2861a70acfd4c9b355f4eb73feb10d6a3e926ef04dfc026dfc15c43da7c2bc473fccdf21eba13a68a4cd809231f9d0a4d543d16ae328bfbf565960d8879a6fc10cc525b187a848c416a4863ea9c547baeb24a809beb517df57f33867ded2bcae651eacfee433a8c5af82fb17371bf378c2221b1766a69831d2c17108b3ceb5d59c600838667da0f4611197bf3c9ca3ed1e92e1b4114764703d7c641abf9f07bfb2e72113b0bb64a8db9e5f7a38baf7107a3b9b1286d70dc94c011cb0e5b6cdd4c2b0b9c1e911eddf1365936860ff0a988fc414cb051be995868af2368654d1733a0767c385970f2edc49a73505a59c34dd8e0f403f09babbf9a0441d5c084441c0530f51920a69bc3786c91263f3f4d3918747f6eb9188c202812dd29f04fa4fa420076fedf1f1d21de63fb9ef63c55376dff9bd093b079bd91c4cd861ab3da6ed28431c2d12db7baab6b19b09def869e43578bdbf367f9bdb5bda6f103f33bee27f4cb7271730e3cac5eb3511e6a1214bc4ca32194519f0dcddf915147c6b48291562f5a65cbd25c088910e08be21e3ddddc10bae9dd2a06b4468b53b501c6f8f9cb9ba7148af470cb12049183bad064983feb6fb95c31f2f438ce074053370cb983cbb1ea2ab13cd4c39caa3fed07f06dd71072bf7eb8466c1d20af6ea49978bc7aaabea4da081fb42e0783d974726f9c63d4bb0f7ec3d30cc1c69875fc1a8878596f23cc45d9ba502e3414abab6dd80b67d904551ccc403e6393acdaa76296a5342f7c1c889c461aebbf35b85a8b09ac24b7d7952e4c6c186ea962b5e5e5567d4a9b41fd2ef3b28129094cd2bfc7f2f33ab97952dcbb487369813ea4ef21ac3fbaa591cd22d1acc380ef7ac18203a39c244fa7c26230e5671148574032d3db27269da7afe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6252d2b3a09ad77d4322935ce9b3b5a396f4c8e728ca8d644c10bbe337094ad53672ac656d2656d3b15c09506bd9237ffe8056f79e4c3ede4cc769102627e9eee696ac4cfc224d0fc4ee47a59fdbfd3720ac92b06ed81bc649efbb112b2f6aee4765232a686d3dc6e263b992c3ae3bf654ce3fd107e95437b1f8d0e8d1090a2332df77ed6d41b9ca0a58a2d372bdb0f801a8f1ce364c9df37c423931ebe4550d1927d159ef5276b547938cac5522a16131a922767e2301c4dd47433260151a4c2b0679d60f60e3117a96ec040c19529805c766eafa3c56288315eb0b7f4b958a0035d2abf035a4900757bc710fd0b94698ae6a5cbb146bd01c16a4feaf7332b1ac8a46f096a485680c30455b8f678f66380d7e6e497424304ba4ae53c51bedf45eb4aaf729325cd32e4dab13b69de0a049a8e79e4455acbe2e9d3c577b30a2c12b657cd68b2ba8b510c878148fc8af1b1d9d05b0a86ab8ff44490d0ea9490bb192f15ad28e89063455bfaaddd038d55777349a307a57f507ae32156649c419a4e115f7cec3bd7ac24350037905bdc9cfbb844d437ba352fce3560afd486c00120aad294b9f6643bd49160c543e412b9d54b5338932d43d97b83ec3067c18432391d2e6b5c628e88ed2612284d30876d1d1f671c4dbdd46ef8a73fb6ed9f96df59a3358433beb3ba4e2644f8319cb9bf4df83b967b780f8f7eba95102e97d2c5eb1d58551a24f26c985da315688f348a637a8029f069513bff81aa7f5c6d8f50ac5ab334920f45031c11a152fa26e49d3ce042be63bdf5511e7cdb623dc6f9dc7d9ceddbb95c00a40834a677281a63b3168bd49294bf63ef6599663100d48b06af944a533aef9490a88b12a46c0f0dc91de9060fae3b2e08ec88d95a310a37d048542b0130d7044595e6297d2ce1908967155a5686e6b5d7219bd470c0ac9f844eb66acabe09e2c4f4e4f9ab6d5f12d50a83a5d2c43d68394eacb17ee1016375f5895e8c582ac2728ce8a7f0b6b083637e002cd92051f77fdcc1ec6d1d0369ad0e282d30cb9b0ca8aded2e46552e7ca0336b7fc030d35ee167e728d43058ccc57e88d18cd2c9f5459d00a9e24be8d2853c33150a2726a76055f508393d8bec29212e26671afb53f21f394e213e31502b0c720329ba481b0c92efaf169f941a4da9d6daac0bdd82aee504fc5c2f472870892c83a4fccde931e7dc5dcebc8278ed0ddfa1271554eb50621222bd8f5e1b0a4b42ae9b31d1237aeab3ed3c1242fef5182ea963dfe5b99c9e6051f50cd2a44b8e37b0bcc5460361f3167a557970dd5b9a9c722db2059010e416556ce4604da6bc70225faf32180a713845d521a2fe0ef9ae10848591609968d28fbc6b7e1fb568a927c098de367c52313aef8b67468d43b76bbf08ec41b00c559487beaf022de27ee236c765569b75ff8866e0220e744;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9b0c699ee8c156466d0a0744d98d19e1db96a309dca7cda68c89997d6bab1830843bf345842ad239acfe8c8a661db579dc33c3e9ff8c0527613aea337ffcd7c1757076a475ddcc7f401fdd4523b6396326a25b6fe27071faec2ae364300b5de17d87fba819ea2d2cd7bfb52b7e9f38b5fe05811431661613b5e9eb3ec4ab680fda91eb3cfbf02a7280efa9c56719437924755af975d2f2b319f7a4844c21442150635030d8d75e069ae47942c2e71db5266324873db2d13f707a1afccd636738f60be7c108b34c15518c254763fb2e371a5a034f4228f3717153c7d1027e66b7ff55061f9dcc58a5f117238211d4c54a98374d31a97a4a8be50651ab593bca61d68a39bcd971b3cc4ebc24df36c0141009cc7c013a316e9c0755e3723066084cde9c021e08e71f969e05a57c1ef4a569759ef64195ed1cf932556d6cff24ca44e411ff0a562b8bde83d65eb8c1dfad0615c7bbda9bf9b98b77c3404a4a1fb9f7a6903cc76f6ec167f0fa6ac73cca0c2884fe7b383256388f9f76deb603fc5f8c796c903f34f0777cd5b5a4134563c3b217af1d3708bbae2074133401451948d62af9430cf37d8de9e9b4d7754a5b74307617ef1712b621ff7426a1d12541386df9a294b62e2b68b207aff0fe50cbe34bc835ce254991f456d4aad921f44a74ef49edfacabacfed5ea86d125c43536ddba037122dd68f82c719953346bc84e7be1e68282a72778fe77ff5bd5272210ed283c0c1e1a2856e7a1855bba6aa2559e8bb022cb3835352aed314cfbf1a29a31f4edf6aa9121193343844daa6ead01c0f5a6c20afa809ed40750142e674f072386ba4ace2dde10f060c4e99cfbb19195ed8a35cfd45eb8a83f7d40e6912e048b8f2091eba3f0d59cbab574b5cd9045bff080d8362f423f0f05c2d2f60d4b7b2b29ddeb9d6b74392fbf083b7a761a01477ba4e69c3510e00a4622939f7003a329e68de41988ddaed2fd18115e2a7e442e25ef9ec293d76b46219f77f5ca0a699701120d6e02cdf889a8474db06c6aeab0c8a31372eeca2f6e780e72e6a20735d709d7e89f0a99536336032bb858bcac585304d67a626cdfce2095db7c0bb377b1eabe9f523c173fee651d804e907cbfc78c9d6a04bd521967378d867ff874da55083880950f3b20ddef707e84a875b340da381830b04831841c498abaa12be7724297d376dd0b99fb23f9f51d4797eaf824ea7093d37af6e463e6fce66137b26a6f9cb4e456589abdf70e3ca5e8da4d52b7698b1e8e32dbf2ce65eeb1102190d185ec54ec179256d43f5bc01ac5c1f793eb7777fdb2469ee881825582ddc4203ec73a230f4b02fc2518c7f0d7367bd0f8e02c25c89fc9a59259f6de68ef07ade0698aa916ab46bd6e624157f61559ec09bf482be108ee8170d4d49b23c0daf74c3552bfc97d92624cf4601d5f03b2b9c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfa5223c7fbd5300533e25ac0d0a1ff75e853a5e50df7db5450f1db6a5506223aa20ff4598f384fd2cf93a28e0428505b7625c97fe8cffd984e13db0b09249fc06b84653da269df005079bb262485dcdca66261ce685e9409835aa866a687f3043a599ce6dcac00fe3edfe4e43f7d54671ea420e7d2d87dd374c94ef1d09f7ee6f53079aed949dfc914739a32f77da4767bac9da9ad2d148a43c5e7cdd8ac552d2660eebd972423b1c1a40a073da5a623e004588ea2840158d11634182ddd51b541c7cf6cdb1c3af6460f06c848d7d96626f1b21ff55dcee7ad6ddd3bd629727871376ed33aff536ed5424dd919d8e48a0c53c8534a940fd63c8c72f46c4b18f547e2f1d13047eceda8e142a6e8c3b62074257344b347bbcf7632747bd70f04bd7784b9e0ce5aa13f273ed8fb324319bf108903baa95cd6a71fb1fa2711540dca5fc8845293ebea1a8b61bbe5fdb843b7cc21342a009967b9ecfbc890b57c9f6fa8397fba7fdfdab02a4410b675c3a5921f27be04a03ccf8958689f900489a82d078ca51772c3b64b12ab83fcb496d1a46d6e1619dbe58342dd01a99fe3f74410c35b14fa52644e5fb6be90297ebc875264c526d0486dc75942a261960f6a3cc062619a16fb3a9ecdb389265779f91543d604dbc835ddfd388e260d623efe4f33907e8189e0996a380fc9799d541fb5af47128ff15389e168c95d8bac800dd1a8b34c5befe98deafa3e0d9febd0b45adb5afb3685d3da22a54acfe7f989269f0d35be6e4d080af14dfa5a4848533a3ca711727db0c632d8c0684d10e19ec29271aa11f65b95dae568ff8768b56988d3fea69fe5c6250fdd10fd292bea335015982c1e8c70434a3b337f0ebe26f19c4562334e4f7483b0e621d57ed457f39e56f31be9357adccc4c0f71505988441caf0ff4290b8f2a13f866957b34adbb9ffcd7852e715aabe998dc3c97f44c365ed0647f7d3a4bdab6877f7b08fe1d1d1ef00bd28668a03733e6d53d2b64ada7e6b3ee62178e602709621218258a2929b9c4e485dc88eadc5e791bfdb626b6bead0a83ffa78804d6f29721eae397350221aaa5fb5f4998a05c35630e5e4277826746ff2c111d6f548030dad97f5d3a3e4225975bfe0395395032b84abe798b7f925e727152293b4b1cfdec6f7749cb378bc86517da446d690be45b38a2c0170e893f7faf5fb4f11057be0a1ccdbfeab7dd65cabea3e11be2810d4563c146b168426dafd65c2b6b8f0f65bc51a86b322eceef83c46d2098a942b2ff475388c785eca545cbba6d3303a617e5786aca46ab57e326d84c3ca53e5056425ff351f3c33d9636ba2e820dceb2e36faa98927a6dff4c91d584d38777735ec77e8716a14d5d017ba49cc7d8a7a7715b69c48b537b17626e4688bb214ffddd4384962ae4cf292d6126981544e90444ce17dcf35f06e6cd5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he604f679ac7ded0a738b5d11557fd5371c9dbeb48db06cf899739a891500edfcc88ff79422986c4584258f0e25a21ed8331f7ad91088c658b7592c41ce95c34ba3c4090ca4fd4f888297a2d208458dfb998ef2a3e962f9c03e1ba9e1fa4ef5a7ec7b3f8a583566a35dd60e72778b78b048acba6ff5a723e1422f9aec575d9fb6d2929d7a4c13c3bae74a8f853d9ae20274e295db4c29398fe36c80f1380ad4bffd7ebaa84e1c3e716dfdaf1f58ecf86df59e17928bbf70c70c0de687b27c2410cf28cf67c6b1a6fdcff13584a493aad7cd8737cf4d3c11d3869c72ec2a6b035387507156dcdb007e24ad71bc982370b0b7034025ace0c2a3f38b277fb20a457780caa434a4330ce1af645199014dddb700bd8ed7ef0b04f05868d797be88e1ce9a2491e53e8f5541a3acac5676b9cf3fecef54723afa1f1aa4148e70ecc7b20f972d3a57d79a460a640584e1b113a076bdca765e31b589ebf611cd95d877d9561f456948dbaa108cf272cece7dc7184eeabf2d3a69dcbc3b0a4d50504396ac245f435f8b0a528efcc2bbbc0b9be35bf12a73fc4aca4b2fda642b02c3be5b6b92496516d0a329489ac9a2bada47e3a0bffbd1d3dffeb220d760133cd0835d35b12cba8934da7486241c40d3d8da8e27ee68b5c8f8aa67e7c57c47cd0861b94456129bd8e50a04da0756e14d5878ac2606838d719490edf373121311c5e5ec2a046740eb4a7c2983fdc87354690712bdc3cc6334ea0042555e9b18c1c79f179de29445b3b90fa365a9f96dfb096bed29f966b3a3d275282263bf820d8135807c8bb3fe9c8a5a3dfdd6b1fcd598886acb4ec73c715c1ac3e6512da2d47fb683ac84451f7633c49025b38e342fdb7b7f7b1de55a64cd8fb671da8f38daed52e4f134f061a3b45e88b34a2277cc2280ffc5ca7c1554eea70d4bb563b0afd36a7fbf9eabd909dc788682a51e25d34cbe3502b11de84f2ac8ece703994d4a4105413e990fb624264e644c29829d072e631406f56a6a7cb0ae164559a5dd720976321c0f8f5e6667eec115613a31cfe045fc6ce2fe1d00cd0539dd6da41115cc202eea1f24b431513f14c0bddc2c8045a46a066a7afa1972c2eb2027b05bdd098f8dfdfa5f90039519f464b75c67a9f0958176e538a93e2b864082f7e7d5ab4e8fd86388db864d1ab9a3b5a8be46a69b13f488a9e353ee2464bbd567d21db268e72a3f9474a98838be91d8b4db872f95f444e08a4fe797ea7b06ec7e39d2d266729c1d2d057127a2a1379da89fca0785c522a2eee6250ef9e6d157eaf4adc8449fe78ea071a63cd94e08ffea894dd676226325fa43e230a98834c95c04fd77ab4595452d945a69bf902386deca36099c2da925100c51312f7ee270d6832c3ecd11e21dd694670d16b7c2faa80703405addc648b7a47d0e4604ee2d629ccf069e022dee73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc204b48412b336f1ca645d5196b8348be83cac837babe922c7bd448940d7f393c501a5ef8d02406598bf925d5dedef266037d836bc582e00bb2b1246c426c37bdb66c3845abe95da18146ae69587224eef8e0f557ecf4bd580d01a8c8657fb5962cca3e37d4bc8fd0ae00db2f8df479ddee8e5246d0bf6968f0bc04e2ef85d141ab6b7b1d1b898b60beb6480aa704bee6cfc172c535602c31844c268ad7591ce73d1b95337996d4f54bc3e9717e52cb1f35670f2049bf87a270975fdf63ce6624e56e3c436d56792864910114cae2973b96af8a3bdcbb3a8bdc0a1a97e00f52cf688301d2b4d6ef140d75d69da23f101b725a274fcbc30ba356b96bd9e9800d2055a4e210143889bcad490f0f7e8193fc6531872fdf3dcbb84e5194c669ee663df57425d2c4bfe1d6300f5f024564ab3e5b9faeccfdeb61cbc7609248deb369d9192a35bbd613b2d86a4d951105accedeebd3b5e50e445003b2521b1f9146fb14506d2e26a8855a1cb66beb6c1485eb55187fdc39559e578a3713cd82d4b4dc8f38859f70dbca74979a933912b858497724b06533236883eb1d8c57d5fc3cb0148e7bb023fd9154b4e9120fa5ae239cc217d6c9828b2c93ba26694538b1cb61cc3d0e6a291461686df8ec59e8c74bbd3a27b9d1834bf9f64b541d91f2e5f8216d1208c9c34d0a06cc7ca9e5e7d1a44989295fa4429a6346f6cd99c510996f9ceef32cfc8d8b82249e6651d38195784a73c56d1911f0d520e035551034ca7cc8fd89f3e4cf8f65a22b537a3babc23b0bb2a75315ec32ba545a3dbf830d64ab3dadd2e084dcf6871c3cf9a6b89729d6dc316bb1ad61e15fce02d7b5b861f161303e50ee7221e9d07e12beff8e3236b4c679046717fb0537dfc4afe67cc714de4b666a44a5c5dc9237f6ce6000135e36669da5a9ae760cfbe43da08c0c408ddc663913c839c9ba89e7d5c831f495f0a401253fe3f4c6f5ea2a8c6c0d3bada502960ab74132f5283761b633fdf2dacb368019b2e2a01ff31b3745a9c8e52511a3e08978b308d8574b36665abf5bbbbb10cb1e4f1a845fb4c61412eddcde467c5a0825ac151207e4f0b38b38274c7649c6b7ad4b1de9ad88a3a252e82a84088765cc10dea3f6546685385083f7769016c7b404e2fe0c1e903a2086c6e61b78acd1304bbaf94ff449c778cddcff7166c334f1f6d1fbbea2bd8dffbee9d3ff751c3e28419f9afb72f8645ebc5fe1af1a795012c7f2ab29ad9ec7bbdcfd67e896add8492e17afef269ff61e0c2c5522ef5ddd61ac837754f371f3902a6d9d85461ce2b77cfd7996ef3c174013ef7ab7f5f864aa9e76480005169a16ef807f117832e4c7f03605070b32b3d5be018a82e2175b20c1f56049d764ac1649aa38250d95ceeedefe9bfa8a8ed1a78f4f65b2cd1f5b0c44643b9531647d0701fd8074d119b0bd6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9a46f70599a0f5854d8cb3874f787bd1746a5363d01933df1d84bd89d725d042d64d9a58b58a5152d350eb89c8cbf0069bec019442aa2642554932f212e5d811f3a0cf1a7d7a25b0125996503db57ba66a6324eb63cf0502ac317609e7f44d8f7bc8129b444dcf077a1a5c781061b6a22c053ebd9fcdb61ff2beb2b403ed2f00c11727c664b03280c1b01f73d81262cb2c6f4936f86da12678a98b27d94b3ee5e9a29faa234c5bffd5a0ecfdbb9322ffd9cb93de67a0028f166acec6406e2c9255e2e766e45596edb594307e36c26cc92733d1db9e22f9d45a0014ec2dc561440f5d74417194c2bdae3206e26623c22d0527a90d39c5cd1d5b3558bb1eb0acbb7d4911aafaa76e3f2b0b99b55dc6ee68f2be07868e87dd683278296b25546227473b612fa9560e5365df44760a6422521903bc2503be3790f437521bf029ba962296a9b1f5976ebe7f1d5f7061e674113be2953f9adc980af6e4d18d68e9356782d927dd3d375614f10448ae09d2b4443143874134eac3314e9a7f2392a9c1c6fc6f7f54a985754ccaab456d308c0a2b39e6aa764ca707b2f6264de1e33ebf61a1776565a382ddcd47fdbf00abe45a1feacf412be6f46f9b27d9c8014166020265374b09bcd29985eee3cc924df5c5803ad7593960b72d7fd9dc539afc0c0cdb5ff85b785f913548d55b1abaf910186ca0ee59e6ec69ba6aca62d0b0e0afdf0791a841e96f30c8547b2658a5b0f21dae1174996ddf4c974e8b5c7174095272966aac683167133e9f80785dd9352d8554950ef229e1d7aa1060d4dd88c37dc799ceaef4493c8909c5d9c2c5eccb12c5894f47c674bc4016d6a1eaac3106f3f0e72409bb836ef221ceb442fa2fef72414c62d3d37570d42cd8567d2c2cae07680d4056617d2752d9352d55587f9b02dd3a75b05578b6262e6a4587773e30519797cd38f888d66b37b1d11f4bdd1c903e5c0134bbbce04e38314e0f74eb5a37b2660db5886ad7efb0889ee36cc0faeb604358e097e9705d6f6cff917caba94cf7073e05c606b8da02541bbc78206dc688b837fc909f471066e1aa14f27ac8c22b03a8dc75bcbde06aebfb56c432a49321c6d0cab7c1186898e8a7bfec8445e374be9ea7a8728f87d929df51893c25a3e0f2a47e741e61272a328e1f338a0fd4713d8d36af0341b10396f6a2f88fc28f20214f9d99f3dd836e2f59fef598e807e6a05140b8db9f84bddb9f80a9957ef0741108113038342e182595b8e1756521800d9cbf9d53f126abf64f9fead3218e60d4e6d518022b834d5a0a1815d8090cfd7c5e56d7e160a05f8c539c51fc1655da767f5257284f1e03638520cfd1d280af47ca54bb0cc7b15b7df96c52ea897a98403014e22062455fc394e96bd085a7713759e90f33258923e2dfb3c8d3fa02d17c1fa034b377a146d5eda86d792b4544ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8e6bebde722cce1d9bbb8e96812a5ab7c6b6c56af2a1fd89d17d4deb24dd218b58287e0fd9c0adc856bddbbee830f3df07cf184f562e22552d87e2410f01259d01bd43be0d24e1e2d43c70f438efe6aace06743a35821a3286b450ac6447533106c3a7c61ed5a55b3fd4e8c5ed2e9a7a4b668e0799d6806b29d29292aa37cffab2641a22f8f4605c7a0e4dc438dc63f8dd201f52930e48630c07e2adc91b9a3dceb436eac77e417f71928811cab655517f80dc611c8275b7e96753ddb2849a97dad090d40b757afff20db211e94e37394d5897c30b2b0021ebea049b3fd5397fb44de954a5b0965e865af35a7394f5f34904abdb8e9a139aedf97ed101bb1a9566e7762fa86e188352ec5a14267bfae556a582c228a7ac30cb20ef74e404931a87dae6e9e2e17a24c8884d74f943fcacb5eea6dd3ac57c1a5477a09764f3216fe7be5f189a630577c0b6411581fdd75b62ed9dee55f80eb2bfb82d503126c2e75115bfa539539e381f94fc4ce88827fb4c38ce149c3a85618772d3458f488d3f07a21cc36667f105369c3dbac9216fb51dbf923376b8a6a0ef861a1cb41dfa7b68782bc91e0591ec9d63e5848ab19f032440ee22489695554f746893967ee196648fc207c1d6181eca77a013be2d4bc2f7a4ab90a90cc58e875d6af4615146867b7c527bc8510f7597dfa075a86167b0e4d986e3de42a1471b0c0fc9cb915697052b25ebd4fed18127b87275810ca5f04e1d731b76d87efa844c6e0832f8926e922db548d386417981610ebf5afe18ff3c07345942f1125fdb5a2310328ca133507213f99f89436d1d080b0dcfb1959c381f27f934932b9b2b6438a83ad4a97733c55c4de4d66e7e2a740f8fb3a6fde36cf493fbfc987c8fda3531f78436439840f0786fc39060ad0c94be1ec6b970d3fb9468d16d716a8a5d9c3597c15eafcc214a2c9f86a2cbf9be6647e2ef8d08d68561aba4165ae5939118571386e56083e273744c89220ed7b0db40cb6e21b1e04e6d7e845aa2468133e2f880e00f7fe355787a4ec36eadc2b1e3b404696739a9798625d37b89f5495c1d414bbfa06a0bad90ae89cfff0856e39ac0843b9c29433f3a4182da0f2ac199372748cfb93d6b186de7b77ccb2b043e6ae9cb8a1e97eb5fa4ec8a8e14bb749ad43d248cb855d67e28b4d35ea83629fdb34ab250b048b3e61b6f4e5a3514e2f104b4f0588ccfd34986c7f0d8beec2512431505808162b31e9da8cebc7bfd29fbb702c9a24406b10e88612c7d1c47278e3d363a86d71e2ba10292a463dc8d62a820e8d72ccc7da5d6bf92d257054f024b17f0bf4db7b5413b882ba5a4105fb0aa3831d789a956c922a704c8de07c5b5d754ab6ff33236ec993a68b81cdaf85b9a43bc00a60db6bd168028c4723911c69adb6e0e9fff01ce56940313ed9dd4b6a88b439765a4b793;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'haa506a07d903364259a47f4b05bee4949f21c6119a631223f34e66be3c2984dbacbd429939a71a2e04aa998e7035bdd86d918f6dc29a8ea413f78c664c5e8257f085abc1351b34bce717a2824181f64c70833296913eb933a2c95e2f7208689ecd847c0d98bc95cc10e3849d74435d79506e08d7af32809c1286f6728c1de861837f7ad133a67821d69b2fffd4721a8121f2224e2e35c1b709e9474b127536de11cb05185223c1ab73a7522b295e5d9c659fbea5498d742052bead4b6b8caf6a06138e075376f4071a46da16f705b5a46abf1a86eb5e1ee9ef92ed7dbdc6416690f5d524e4dc133a298c13d3da749bce473394e9edf24a73c11248a2f50d0eac3958b9db20cf8b833ff5007cd3bad83f9b9170e7b0a909a6d11a9f86d83bd6f018dd38cf16baf4dd4fbfc761a18273cc76ac837e079929cbddd1f6db5fb1361bb149a3c2218630e942f42ddbacbb03c3aa091853dbabe3baadf91e36a35430ebff184e67044e14eba65ee9ce5e9adaeba0cf71139a6d52bc34de069e49d285902755ef052104efc3ddf97b9775f9d22acb4d5c5fb4bc5d55a9134526677fa9b7dd33c36976f3209f0729fe8d51ba6607204fa99ade6d073e7497e5c5385bcb2e78f220e2a8044fb88d3e361fdd0641e900b1ddf97ee706b5056dad22c3a438f9e7ee193dd10d0beb1ba875c26fe823e55dbfd1d7164cdc3c34a9dbab9bb42e2214102eeaabcafd753d5d7834acbadb184844ff6462a7fdae5d1d2f0bf8723070ddffc515ec10f78ae92525561cc71c90a2d2f4665c228d05ec94f66f39f4bb398b99da10c5eb67299fa9f4df5b3494cf415925c7b7d60ef9ada436bb47500dc84a37a649357b64fe316b5a9f05848a39c30009f9f7e7b153c49f95339d6b79784fc0827adbf99b132fb5068ad7c7e262c2616c0458f7fc8045b893be90e9776324129bd916d0a13326682bc6d76c4f5689fe602ac1b9da903f0087bc5c7b62df7c27bc1b6d1b54bf1f56f8dbbf501d01f0d4b00713084be125d58a65208637b3ab7a36f220ea9e3d82622bf7e6c6dc014c77ba1209bbc3b75f8f1fbe37e5b12e823bf1f5c9b763aeef1a03a6727e135a1ddaab25e1c6bdb4eb704b3d2340a6ad1d6f99d5351dcd4da7dde9463c9e0ac207f721493d877d95e3da4486918d884df70a5b14596a4e0f1de1befe5dd010c957ddb36eec89c1354388eea912dc39ea11a8479677c809c0bac1dc5696440551dff8b0146bd724ae76c0944c7aa37bedf42a375b1d3bd58919db4d33e7b766c6d9ea5a5fd03b1f68fbd5aad596873dc47981c21c04cf0c73f350153065b7833464d4156a17fbd3fa273f72014234b73d2aa516ea0f7290da1d3d1ca56dfe077d2548a1e42804caf65fbc6bd3c0394167d60b04ba150b7dc6e3bc0cf42b66f05a814305b7f8161081c01de84f6f968cac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h921f48cf268701edb5936ca2ae94a977448ea019d011f4ddaa2f9b819acd13f5dc502e909888f64077090a6159f11a8c4e9f6b9995778d7b9a10706e6688559f44aba611dfa745c22fe42bde48d11a5a96abf04ffac5245e07309e027fa44c095b59ad08c19119116b6ee25a89f58c694f663782dbba6e32c3279a9587be6cb8af0feb8e7ccab88064b1d4d191bc631a85e3fdd9531cd361f967de8343716ae68d6e40842372d4863ac5e8c6bf9c79fefe747b04685fbb0ef4a2596850479675f5cafa6d5bf0919ac45f7d5ed81b8fc5989708ff06f43c4eaa803ced2576c8a2803f9bd4b6fd1146c4d72f275af92405b8d70e9a944c65f1cf77759aaffa69c2412618140216fcf1ce7b50cc3dd3e6225937393fa2e01322f304abea2001a8d226dc3ab62f8084db45afb9dfcc4f42f24babfd0000342ba92a08ec98f5d73106663dfe2d875a12b2f3e231da5a14fdc44e4e9e0d01beacfcbc7e48261eab70f54f186628d92e49116d06913b13759c4372b5ebab2ded417171b86da1eecd2b0cb1b56e0efb7b4591cf0e4f2b106bef14adeaf3f8e601414890c3b279ed69e3064ef94548b6942cd1f1487a80fb8408185cf9ca56d912e21ab6a747f0682344be36e2990a33a9723545b765de35660748d5323b844db7fe54fec7a8f248545923de8a3366be1ae9107c439ef8ff332a522c867af802966b3d2c4eefe82679a76eb89b658c04d4e6dff2a0774d15e75525e52515e2eb1905666a1dee0e6dc97f7a4dcc2a270e5902a641409cdeab866aa4a6e4679fab63dd0eb1b56c67945ad2ba012339ce43289e3a241fe9923654d401c9eb6b210760904a160238336bb0d0333f2217435e0f720577b9dfc57182a9d8c3b6f32e6bdde6ad2b60e27e4e1b216161925b900bc749e15aa292041ca5910930ffc1dbb4b05ad55d9d9b306cf127ba2ad27ab66ec25f38a417785eac9b1c3b0187d6d974cf408003d012d3e25787570d5a7ec573a51d2da2fcbd9429b77353446dce1d4db7cd48706625f71e66091eaf2ab8cbc0a9a522511561e315946132f00b3e3ce17c762d0323337124983f7cf46d11fc917bcf4630ee502ccad08e92806f3cb21d01e0880d4272441bbdfc5dfe568f8a8f19c0fe910e942fd42b64312e47500e1b52b545e68bc2d6d4319eb7428ad7e131982bad4dcea11f31a407bed6d6b1a7ba052c5f53772666523307f67fdf72a406bec61acbe8982b74cfad27798f107111b83cf76fbf75f6ec9bb69b2ba1cb924df378655d390158b8fed65a9f52788e3307bfc2c7a0dbfaa0458fc02b967dbe44cebd79f1c9e550e6df0594b942ffd02e12a3d5ef45bdda2d97dcd5771c5b05a8a3902bb36f22076f26afe8a083b03e44f72867fa649562c3f8023b5ebb7ae67be4f7775c96dd7149e49a9c5e06061f430f52b9e516e77a5abf8636;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h97f58bdd14546685540b100350f107c7c63247590f032d6d5024933cac7129365914f7d0dfdecfc9846ca41948eaa8d81cd046218932dacc3661f6547454c03a5f25ae8922b5529d1d5a47b986f99ced9f94a5a675b6eab42c05782d3f247f563214ca5670d32a4185c8bd72c94f827f1ff952a76e04a6f57cd6b6ed14b782c1d9311bccdb33577295ca4aa3d49a3404821e0e641ba3623d70aa442fe897e1862ef499d1f7554b4cb9385d7e5d628155c3906f975c13345293d85728503916f92d5210efe73be6aa9fcc55877a7d2c358acf32cbc62d9d183ff9ce60ca1945f41a8a063d09a20c5d6c16e2b2903620ffba9902307b1082f4d98aca2931b0bfb4862a24887c8cd42161f9fb3682eb72155fcbd9dd67215df52874b0a18b76b41e420bb9a424cd0febd6c90a622f69add5702e128811322f163f2dd60cbaa7c9c12d1ef3a27a43163d032ae5bb80925ce321a3e604abe63a7f97abc89357799e87a322f03161e69f3b83dfbf6fa1b75301c3819622919f5f0ae2c86b5d88586338298238018da8e804a6050c2d271fe1ff6aa141a07b3dd61793868c37b6fda0c1a8845a5eb9e9107e4f4d429e1952a447ff370a07f8f6f2bdac27eccb81fe286ead4858d4f3f43b0bbd01b475f23da174ba32b116c75247208d0991f9c2cf85f29e47b4918120af8ff16d7e2fb585411c4d55b43a0ac1aab40ed0b8bb6cd186dd3ad54d16a21f0fee0f7b31cdbd09e96b9f046cc2988d0b0a68c4424691f0899a6c17206cb7d2fd5ab172e4899b932626f589ca79e93e8f7d798bf7512f7e6b7ae1077ab0f6c51ecdb2d6ccd06338ea8f003dec3c6d03fb775d8f255c018589e268000be082f729d97eaeefe8277849e8fa763f225717cee2fb23e7d8a06dd655218f68de40b6ac7b2977842c68c73fd009d3664d661bca96ae9ac4394eb581e714a3fca0aa70c03214af6c8f708ad805d06c1286e9d9489cd3eeda8d43c97a1cadd39ab6e03c11052c20013503711e9ad2b58dadd6144436cb8a9d87c1a2296e3b25178123c994b2489c5d8f2da1c9a2bab65295ce79ce0551df2e788a399c5478025a779c2d79706d7eb21384221bf151b66e985ac1fea8b0f35ed8aac453a712f4038d7bf6448df380e8ba627d0a311fc919353684eec2757a98e06898f79b110f9c615e95c016cff848c8d9188004951ee82f6b458d15cc660cc15ce7d5b4fa89316a46e87bf83114907d64fb222b34f44a1f09822f1173d0b81e6df86996890dc44b5e901db2115930540d75e926ea959d45950d5b9752e0f8e53e0c07ca261079818c98620e7fa1732191ec0868f4c1fa3bd92f6608f8e4a538cb6c841a3bfe87ebe55d2e1da690ee9e67588581bcf99e0ef37cbcde7e82ce8404377c04cc5007bc66a51f1e81be8e43c439b1d765c97768637a9ae8dbd7b2256dba09f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had071580a20954e3c08af448152c21a006cbd2cacb1c6ce9d0f4bd8ccc44a33ef9ca1babd144d36b1622d23d9afbcb95a936b96412c17710a8e00afba3fe26d214979181f9da8c527625be03005a26ac755df99ac15af5a2f17b0a9dac553e9c78374d4b6986f693b683aa8aaf7dc5d90dd2a3b9b4fa1a737f435d8c5737825121737f315de5906fd3ce1e9abe50d4285d8b813e004515603dc1914687e790f03c7136f7fac207e4deb7baf782cd6047fe692783268e0d34052592725e36b3c2c08b308dbc32d54c8273dd9a75585549542a7799a82a0b2349bf6018b32dc974b7512761158b0f5af5e4aba480f4e0127147f1d45b73fb5df22550facbe84702c562190637fe79fbc8aa7b3a0e4d5ac70e5ec01db68a99214cb15dbe346bd71fc53d624e7bd35bcc427286fab650ac2fbcd035338f4176d1cd7f5f2334bf7259ea8de04af8266d643c3561526977b5e9598f405c2dd34f9d82e467e95fa72475bddd0047d57369f6a2186316ddef70c0172d0c4e98545388793d66466a807f41b2c4f416da8819530a46a6bbc74c36aa5384ff11fe0cf0886f3445706fd4d829989ed6b23fa8ab6b4c42f2249102ec6a5813aaa86540337f2091c5ce1a8a54d93667845a309b3cbc134c924ac53c4d1c6d6c0a87ab8043a89e2c620c99acdae2ead94f1e1316175c697fa0168faa7c190452024beb9b595df8e58a909191e8f3af2dd1a3088c7154752ac028719695df0e6980f2ac3df9e200a1ad06f3d07ef6eb9e7b05b4c597ce8257f5b80409ff5a3cbb3da8143db6598413381381e4f3f61e6c86b14873ed89ef618fc692bbe4405afeaf77a122b4790e8e51d04ae4a18cf9e24f340d48d158b77e8fc9183c7bef27fbac2a78638a6bf9f1e981553626b66206a0e3207041e7c61253c48fd0a42559ac2c9fcd09a78b8d955c280cc763d23dea9b38ecf8f7ad91f118880d765f9464dcb6bb5c63f7869c129484940d66ebf7f3b2d30127bf679b4c5fa8d335a08542ffcd26b7c60b2b8c16bf14aec8ce7f637cd0a8ad14412045e066b9c1440e9362b524533543b52db3bfb5253495c7bcfeb34b48de4f26d8c78220f77a6c9c0853b1064d3a8ba6cee157881ce7fe25f29fc6c908ca7dc82b49c11ea9cfbec67444aa669d3535f6abd2583129501dd06cf69543617de1eeea6ac03909197a5518266ce9a0b3a7bd25319bb43ddfc684a986e90714193c4473135e05a9bc5369502aadc504d2c5e7844bc9579129f5403727340db42f31bf56f9000a6be6a24cbef6ef3734ec270a544ff6b1895a90b47647de2eea239b912db38e99628d63e87cdeb8e0c37d0681b0c5bd5bdf358204ec45ae14d2255cfaef2684194da0190c92a8590b3fd6c1353f47ed0468cb831b2a7b8a14ee0e526c8598e6ffed3def7536a0310994c7cf70959a8bbd92a7c52a81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h444da63763e911ff186ad1da7140860bc4c8922dad93569c5591b7e2952852f2f5ddade7588a62f3a425e55409ad8e4ff7bc48c1deddcb0ee6e933714bff2c1aae122a970055e6c2e8b38d8e0f666ef0ad997622d8f31b6a830f85673c2815dc8fbb21a1b918b1dfe0813b83d62f81d1f9d0fe2e09fd5f21d1707e63e74d325a947e3f833851679feb6cd47fc1bdc7ce9281bd805950e705c44f0b5acc255ae2006a14441d46d50c7f7d81eb1bea90fe37f89b899b47e3beffcbf1aa45520b32d9ec99f6df75430a3c4cb68753ec8da5c81419262e59c54406af3961789f5cd5fdca9c5e9e266b387d990aab812cff0b792f9781478ffd8d3ffe8ddf3430e34547d9aec1ae406a968197cff3fdb55bd631a8042a8366a60f165c169ef185c3c8bdcfd31831c650502a27050c7bb475feb7d9c2f41c1252e7fa2426997e3efc757c2c1e7ba0714065d63fec058d6e44bafe24c4e77ee05416e1e4700b25e3f864b071143c00156094deb982abbfb583c3c4f1678291773032286a692f6a0bef367dbda1ae966ca527db585c536b381e7dd4614dde23554c0094c4a124fd788951ef8efbe2a1e3b830f3c506485e176646859916a17d4f80e78612110b233a44c22eadfa8206fd17d2fa74a77a94c6855e51605386f53cee19e00ef4c04e62499a21601fd8507639f1b2b6fce67927f6e197a12e2eaf9cc506a93f19c58e58be4f71eb7ea741173dea6d55f585c5eac7dd4d3e326aa7d45b9ed0067f695df347c44268dec1f55ecf0159847b13868e4a85ae92fafcbe21c0cec131b0f954a9d2c7c27e2329cd6b1554ff67c1c62de40f68af3f8861e7a504c970e4f75e5474070aea1469d44b894bca1b9c9aad80af6d34527eb2d7fe345e02df65ddcbd7fc68933a96668393b21bdc72522bb4811ee4b9159eb037cb332703db1e4d782aa1f80a6000f9cfdddb896e894ab1226ada95f84955faeb4ef67767216f796cdce484d1c640f647be5f9bfa60dc304da5c12235a3369ce31a0f8e22271963f0e2ac569d0fec37420cb1aa527dc8c5260a96b1fcf486ecb30496c01a4bcbfbd42aa6cddbbfa4ca74e786d838c242f5dea72008b8b2750681437e6366a011dbf94d171afb8624b7f6b9b9277e4fd88d640677c792048415d33788a6893663c5800de5359a03bd71459927310913e0ba38d661c006f9723f297327c444898c64c79c7950c1ba46fcf0eac375f3e72a815ddb5796f29ef3ebcc0a741df6ed211c93a28038e38e512818e1bf7f11c70c84a41ac15e013c913f7839ec2107b6c90020efb4836ad3901993fe0952efadae44769b3e1f4b66ba794cad61c7c9475007efa23e066fb5bb21dcbfaed9ac4e5165e0a561a6456aa1aa4ec28de0973c0ecbb046103a152042807651bbb4ababf21028ada22bef0bd3c90b2c687e68e87cb22d30a52133;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc9c778a7c106cc1c5a1388c3a1af99880de097d26a6dc6d4627eac3bb2fe74975745b7dd4b64cc64a9bbcc667a17b81d2b1ef620dcc3af3ff7250022b08726a9064fece5de428a8440baa92ef11a4844de4568289ee55fab84a9800677172e60196b2aa5bded4f022e478c4758c17eaeb60b87d74f68487749357c3a754a3240f4d9009689aa13413d427ebf43c2963ad586503f59064579913feae0606b6d8c01c2b3d9492661214fee350116b6f16c8e4ad9bab7caae83d42e8a746a586f8b9a9e16b92a2f2cbcc514af138909d52a3517b168eea246c1e4a774a8a1295c7839f1cd634614fff8b36ecb6fe6e46ee36498179866357c019ad1a86fd5ac5c0f79cc7d84093dbe798977b8c4eca5a33eab078da35624259ebeb538dcb07725d5fc395dedaa8cdf7e0d96b506c9628d2af99bd21bd779076e7a3546b0cc6121dd0829559a597caab76d9807db6196ff20e7609422228e8ea699b3fbb8b1e692facd841423d277d948f7e8fdaac13347f9fc14289f1f49c62e15da67266c8d08b561b8b41ea5093d33a9e610561c988f46890dbcc55b0c6dbaa2e8fffca475bab1ade489b81cd223a840bce457002e72640465c3fd9c225ea8a77f593e77ee91fadb8ba5a0daec189216851ea2084c49c7881d82ec2cc9a2dc88ae72eecf0ff756fb4985d83ff0da586da9ce8ec3d045f119f9b9621b396ac7fc8935545606f4cd375b081907221d9f93481b495c928e91d983a9b804084f1fa532bb7eeb80cf4b511f5e7fa35bee53cb4ccd5232c1cbe007be891aa9e154df1a38b54ec730b42649f89ba7ac8ee80388b906cf3dd40bbfb881ea7d43b7adc8a09d55722bf3900f715c7a7795178fd420532249604407a34d743b7f34b2dbf18bdb5d42a6747c7ade54871bb336fa9abc75fef4e4c3143b5b114d05a4e7882700cbd93dcc1121002c0cc5cb70ebc602bae28c7e717940d7de764691f8806582f3a7c411ee059265b862df7cc21d247c9547d52d7d2da360de8f7a4691bc323823b87ffffb3cad60a1101a687c0bcb9f484b81d7a78274b6f6e2b1e6c54f1d02f09113ff1a94a539a6f137cc04ad1d9256bb430cc4bb18cbccd48dc44a8a0cdd60e2a968c8e304f088cb398acd9f5f37fae057b39cfa2b2a3f501979b84f72198cd0a84998667d01c771c156a04630204f7fe69dd847a4f7051de4caf9fb1ff56f04cd2c3a53378b5fb4db1f25b58fd5bc21126f60e1ad92c6dd75fc18802fcda0856b20632b91d5e3448bf64afb8fe1d535418cd1b67e9d7c030a8951717bad4728e7a28b552d1408ef78dea988899efa5f214b8f90af44dcb8c314fd81f5dfddb01688b5fe1bac9d8c515acad96e54882a027f9a37bca0da45c641848c9c4371a4a05255159515ed3e9b0ff3a65259816e3411e434f79e4ab5ed1405d223ea15428a8c96103d17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h412564893d0ff22e77129043898bec98b803c152df615c96bfd30843d6ac817ab5ad96ee8a8130b961217a9be8da43d8c5b845093e74d2d3e8f77fa144f6595f05a790fc7746ee4f4a6aea45cc001d2989346fe1f5e0ec7e6b6fccaf07b9785cce2cdd8c60a4417e8cb8e94b256b9f889d7b92b2568b429395d4ed17a412a17efc1094fe647e3720dcef393e0b70de02b8d9764708e77f96654b61b9387d42c5bd1b07e196b2721552a223cfe5fb7b922a476629932a6de966257675b2dfdff75602bd851b1be96fb68f2d0fdde532e578e95cbb4d4e35015fc19dad06da0968eec2a093514885694a0e4a587ee13ab6e305956d383c921e3818d7024aef99da4c519d393d637cacd17b9504d66acf7fbfd29ad681e68621db871a407c898ad890ad12460d0e1b898d36d9d2b57c05f1fd17e84a0d2d9437687bdd1de0795e0cd5c06e45932c5acab362bbdda96661d3c5f8d501756bee4adb4b82077d9d10d1177a3c5f2769146a1c520aafae5c4678fe1721b44f715c4b6740faecc5fb3a8541fbf697c0a654316248478c9f5641b79bf26cdf9d53ebb21209956b8041b9b49abf2e6112c46561f6a1088a77b0f1bc11e4e90043d5216d5da7928f7e3a4167e884216ca39adf7b37cc3e1bcf11bb557741938df94b9fe54f8ae81b10e3575ef8e5e203b327ceaaff3b243fbc08d73fdafebc0d16496012553ece34b1018a653429d024d79b64d5bfb0f90241b97c694fcbfbcd9a1a298b2c7a68f5e2d971cc641aeda17e3248f9e7642768f5b3d124070bea2bb04a59192c1e9a48bc898e02255b782a76300619ba503432f33428ce701c07bca9745853cc98c19cc27e15a0f7b413825f8f6e9b1df62ca8d8766228ab0ff630f0af50b3d96709113873a5a997e98131ae5a62ec5ebabac69b46f381e079f95fd8ba81a513dec9dc10032f9c21bb65cfecbf5d81e4731591fb7167726fe698070843c8d1f30dfe35ed3b2fe5e9fa243fadb5b2dac49f7b5df6213ef18365924e8665789465cc06120f80187e0acdedb040edb66adebd318bc80a0aa87a8bc1364205c4d36824f715ac9462b9a6c081edb9da7563735e5aeeb08d502941537aa1ab0ed63a23eeebd7fbe27a74c8921a2a5b8719dc0356c473ff07c18be7cfdcde75ca9aec6aa70238c6c4752f11f4cdd0ca067fcea5c4334b7965ce7dfed7ea30b7770bad2da442c8426354421be474ff242f86efde7569d8594eab7a5aac6ab33680ec951c07c82ecc4985ba8801f20dcb7060428c66cb72e80c20004957dd902ef8c41852be0555a5251b666f5d1179a315e17e681c67e3094b4482c017e078c2407efe5c8d923a86d670c81ecc141c0bd313eb1b5024ac70caac42a2d70a3b0c729a2e81dc96c4d4056233bd720e68db6fb536ea250b04db85e80068b4ad1040c40e8e5a53853e076dd285;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5047679171d4467ab4f8398007ab785becd66b451a1ee3464fba414d71859296302203cf059fc94a0113809892bdf4de6f4d2a06cb97fe46f5f066888cabc7b4a500046a04536b9db6c65765489b0b4bd8deeb4e01b10b59ee4142f3a1574cd8f0690df6282aa28e757700880277b065d29f4a178a05a8fe2503bb534ce305511d18035ff54bc7c8976e64973db60e640218732e1df13131961a88d398af817b2d8b88c07eed6f52bc76547b2c8a66232b6dc7babb38abba29d07e0ebc906b8e67041fe73d3f09cb097db9c938ef260d35f927d4432f22d445d05545eb2a403e3248735c9bc48257232a0e53e8226ade05d823c1ade24de7cf00ec9e5c18ee07ddfa89d25b1e7761bb3f3d075e620c9bdb2050973bf13a56c7644c9e32187a34855d62d693e1cdafee283aaa566f95aedc27bf749af744a6133793b25762f90bc42b8badc00ac24348d6b339aaf320aca9c2bea5b2a60047c8f3ab7c37659071ccd3185be6b3f24900121725f65b5e58e971f09abb2a6eafef5a73ea48a0c6123bc7020adb8d50a879b479e42418742be7a0ca336e4ac734469e79faf0eebcf4b667cf3f68fde4e77fd0c0735399414c2b744772c6ee38db9793bb99b7b770165d769283a31c72ae68c163be34adb4396d7e41b314ceac4d6bfa1fcbe74f033bb65cecdd37958fdcca38e7d2ce1613c5b7b59ae66f11a6f93592f65fbe13c2d924f241c1e83b8e5f75fc3e94e535babbbd02c5bc082f82c9a7c8805ab915df0a049ef676d9f6ca6eb28249c97f53186c62d19b2241bfa0af743477d45e131b045fbe4c4c3070ec92ae1e66944d7a507fe3b95bd52f68e5b22f85085049cefbc2f25071803999548ea402e17adf0921fb62a1911bbf955bfc4ed7816003d9e0f8f5575f90030d7082f522dc7bfb4303fd8cd607b60867270db3c9c7ab143d93b2129f66a6236a66879a1ba0b75628cad00e3845df7b23dcd19a8eeca697466d8c365f9d2ec5bbb3ccca7b39e37a8245df7edba79374c2cf7ae37251f41aec738019448cb1fb967dcecafb3d6f02b9fd279092e88d1e5d7b73e477a9893a8e660e83c38603d33df82dfe9790f15b1a1df8c5c6ecd0a43bd5de46b049cad2d62a7f53fd2385de44e981e5120c97d8210aa81d3ba2c953a616a66aa897846ccf1f41ecdc5730fb9112ac76257b1d492e18d8346d3c32b6e05bae115fe181316033edb8583fd7dffe0c49b734bbd816dd0913f2308681d18880fec356eef50f0cf1c473229e7cfc93a875b2722ef4b07e42bdfa606e9406afdcda446b3d9e4e4aa01c4f3e5ff6b0865b0c04ba6a10809024436e5e58f63a35cae1a7851eb5de0f401874ffdb41283b9d91ca78fb83665271a791d9cf21e430651bc5be8a6df76e9d3302abf98ea9cf96ea0a1ebc0024a385cee43bed7e3a576500f74762919e2934f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha9e39d3fa962af5af1d22a957d00ab61cd2d84be0b463e3132f00939f6db48daeb71def07712f3cf333984b379543a003e55da177a2eeb1d33b9853b565022296cf91946df4d1fafd5f8872f93b485518af37624c8a3a183a1e00c5d070b51b876035fd062de5f30c1fc27cc7b71bcf509e119b46d631fb6c4b371c1e85c18e585156fbec7c2a46f9ebaef4e93b9f1d8ff1af0a693415bbdb077dc52f26860e36167754b0322502d74a753a3331eee9355367b4ce4f79d090ab628dd679d549e873fc95713aad223ed607ebbb392303d93b225b294379a7daee1f1b5363e35eb64ea1fea50ed7fdfe429b77449f5b3db252af4c7b671acf3aa543e922a65cc7c0addb6dbb1ea24c16365e9e4ce09efe68810db03dfa9fc4e4518ba5188855b0a26d86a5f1ae1c90018d2a31a2aa3cdd4d89aa53456cfdb0bddfb058d27f585b3310b497dcd5dfda680944b41f8efb803c42de8b9500961aa49cb0670aed2272849aca387abfb97f76d803a913ff7a9acc75404550a72b04e8f14a7850058fa66200f3d84c50077026a277b19c01029389ba40cc977bc6ac08641564a65848efd9e887cf39c101ee862fa062e66c39661fdb316e14cccb4cb29a153524cdd0e3395244cd6171b818100fe67be9f181727fc2eaa84482b161ebc8f298d3e8372e718b2ca175d67d5a3cd259c1173682521a5111c2c5e8d846b67c682621fbc619396c77c8f54fd1b974e46b5b4b9da678eb2a2a9bad2d56c0fa4395ad9f16f72448e0ffc1d60accf51f22a963c1a4d8720ec3ae88cfc84bb5cc231972b47eca8050bcc79e2785c0650be221c02726136de769c6f07b3baa2eb280f3e7cacf0e203eb5a21e08edb6ac1f5c3d45dbd474db0016b02655a9f26aee8bd5634f395a00c0276bfd7c119067412089d43876c81f1fedd6d5b3d6034f1fd1aa67ef7879e4f112dac074828ba1deec495b7cf191c90284481fba707ed990b02d82b1d5984add2d784c40ba3dc9f014087d0256d758de2e43b0ae0e7f90785a780069dc4fe1a5f28b8f90a512e0cacd2f07dbf25a13f92c1d6f7e66a2095b2335efe5603baeb6e8114b666d010a39a284f205f875493a6abeb9aa0ab6d1fa3f9acbbf0fd3d5463be8b1eb82db4befc01fec94b26ea94140ac5ddd1f0572715a50e07e0a75e98db534da8a3d87249e8ef4bcad43402dc3f36a203f0076d0eae2caa273ba9bc628aa46d0d572d09e14813962fa22c0a83c52d88d140739c668a802a0375c745aa5c51351b91c6b886246fdec86035538686f7ca85fae2ca24a251e053f375b5a6f29061b03ce11ffcadd3793f078ead9d8ed6394ba90e8744c658f75eceb9fa94c28ac1c5f59ae5edc36ebbf65df5c7c508343b0c79de833d0144d3b32b6d4f53e0a52c3cde7f8479109658c9599d32f13f8cf4181ec6e83f83adf151b6eab5c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbda1542dd1ffd7d7efd302ab88d8ac6a2d671494a90cac7bab17f71956360e0ee0c9b80d74da2502e6301891fa5dea9a24ec04a68f5bced16270cd6654013f15a1a3138485f18ff06cc01c5a53110851adf7f28e5cbed7e0bc896ea26d2f7a1b7e8fc6ea1d455388dffd77e2c43d1bb0d93d925923729f0737f65566ba5f0fdebe020448bebb6fea779e0c52bcfca387b78979a0151a32636d44b6ad4715f7da64bffe669fbace23a42cc411a419bf1a655f05f6263093c5bcf65f50a5cc5c5f68a1e37cc7c5992e3af97ee85d26f189cbf14bf03fe19692cda653a6d7c2b5bfc4dd24473824f88517fad82cc53b71a92b1e9d0d997a3ebd2ae0aa2722455f2f0e18db630c5d926381a92b2d767573a5f8edf2ec9755541ba2e115d5196b76a47fa9fd8c283594cd740c255f18d00a39ff2a89a6ef4ea50214e6866ce3e6556dcaf22564c03cc19cb9d1c775ef8d9e638b3d263391454bd6553f8ec9069c4cd3f5ba7978c969730639241968115c974cc1484f5d2c0883cefbf73cc145be8ad778f80aada5a12f521f24b53e59131f6a864dd9e9c62d0ba32c3ebc263ecf30df716052b497c965e5af05ea49dc547444a464bef843cd27be44c92e16be7e9d2849d2d31719fee757205d5c2f039acc5da5a957c916fcc55eb7e6568d6b4d5b95d679869768eede614da01eafba6b96149141278fc64566b7d081ef1ddfaf2859ed04a1e736d7da235e5fc2ba7da143b16199e1b3da00759b1ef8917f8f0c4f0d41a5053256695203829c615e48bdd50c32c08f86ef8ead2d18a690457dba6d11a362bfd34a21ddc99e7f662f1e939be0a1a271ef93a7de58ac6f356a136c1ddc1845df29388bd3fe6c8a251826d7d4553b8cdcbb657f0726a42bd59de8eca4adc444418e099b74b930744ec17a747a96d76fcb8672014ed039e5b8488cbecb019193c1043c5b72ef6ea7eb58563e41ab3f4cfeb78ff9c36b94bb024d6435fea3170695bd573f2d1872041290d3c2370166510496bf870948ed215375edb3fcbd1e36ab9104cf94c5a5348fc721507ff9154c21921f78fcabf5613528ae4585d5601aced2fb3bd2b52ce89328bb2069885fa0fb92e807f372204cdc4004ef4ee23a1fd4c802edfd0da304860c9602057eb70607324089b78406b95c3b330dd4facfd90ba0ff4d294df14cc72b07b5a86a4b2b88baf1d021e578eee06cf2f77417f54c214253ed0868db378fd3dfe54dc202eb05f78d7eb0d1df5295040b8ae36ba8d51c91713cc983b0766d6ca2540f60948134f6a16136734cb6aa1ea7e32341dd98b95021b098f081bdfad39949af5237b25a022cba5a0ef5940c04018d35eb1172d6f544f3c4e69f3c63d63814863725deb6a6016684dd19d723de21c9eaa0f8b7629ecdd11bc6732935e45fdfeb165c2caa4fcf892fd14f41e3ce07b72a7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9012a0227f14ff185cb80b5c83389a08fbf964ea40af924c05060e78a20395d420265b389cbd3c1a39d270d54d68d74885fe2a7b990b8a75a5ec0cfa099973bc6b350d6cffc65212ee250bb1c912bcce6a392bd63529e32b594073444f9611cf01c44285efc1add8158aad4804a693c1492de7a6f07d6aa2e9541840bdbd10cf23339ba4578901add559deadbc7b25a7b1fd1909cc48849dc8b236b07e2be3a7bc5e6848d01892bd2c6cda900b39afd23045d5d9bedc4d3dd62f721ed69937f5f7805787fa09b0da33a0d666ee6ff4715049c20b23bea0561fc653647c0adbada96f3fd2a489d648a6b8e0a656589222da9d1ff75556629fc6560d3f7f54b7adfaa1d9310b382e8a68f6060b2bcdd9ae337a73d9a3aded34def98e55f53b4cd34a3587c13aace489b848f38f62d2b9a44d770435a7909465af6c2874c8c4520d4380d8b856eb56c3460ac7fb55719b74730ec80e72b4c0b796cacdfb7dc504e50fbdc4ae0ef6b0382b386571912929111c66b2d5315deb4dbe2cbe004b85f63a8e156daf6d737c1a8502528f5c638668e372252e223f4980a09785eb027db938c05914448148d0c08571bb3d4837c20e86a5f1207e884daa15e403a59dfc6ea1810613fdc3384c962828b65b623cc7cf9713edf995e0026c5a4562cbe3a4c0295dd85f19192760f1ff1b2dfd5ac020bf6bbea1b1d8973478864fabf6d3aad766a158ade2613f4205edf8be50ef16d5d728b604c85054d2e6099e88d7b9c912a5aa08f52fe1b66a4d87fa74db8c1d6e498827bd5e7f9eba26c6fe925e19f91322a862bd2e589f8b88d8b4ec38937e1a45246dabaf2a7b92568d78b788fc1ade8d4ec0ff0654fc8f11b4640f57185f5ec38bec7aac88c3f0d4488fa8a25832c0abf04bf1dc602f7f0a1ad17ad2eb0f7b5e18ad1bb65197cdaf70f6d44518bfb4407dc2993cad7204a55a358483990bd6c3c3a3477272341bb0717e50fe0d86285c7b9ecc0f56e67102c1404157a84663d49d60ca2c099817e547f46c2a3c5f67463831b4ab3f3e78491536f4ff08849bf0fca1bfa7fb3dd524baac3a07205c2808f37f35ba89cd59c2fa4c333a55be98a3cd268febbb0fb1e6c5edb9193ee3ebda86b6b9c003e33d5ad9a0c9543bcbee1d876b9d97a68eb5ded737a2bdd55cc5224012d7c7a451c9230731f3a8eca90143f3d0f7d6d3427f1b8186a0d0e6bb1450e57e4c7335d8c80e2a22b463f08705c47a6822237e45e5f7b30eb28703b101cd4f4c72bfb89ffcaac251bfd81460aec2e305ed484eddc047d84a289244126dba85ff05d1d8aa39236cd5ad6684b6f516e89c5e8c1558b49451df9ab87789cb1be628c35878367bb1fa118dea06fc7ab3ace34fd273ee02fd25a666fc3fea44bf4db3875f0194e8c4f423392b015f17371fa07deb5665ea35206610bec107f291;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcf05ff57d4a9d1cef30963ef8fc257f4fb21d04c4048ce900e13c9bfebf41cd2dbd3dcbb74bd3f7f04fc3cc7ccc1e02d83a2667f978bf8acf41a10a283b264b26b4f450a6ffa641bae68ecb6a82afe4e430768e18138666a88c822321a0af7bf38ffb14b8a8dea6f9cb35a0f9ff431cedc08f80abba50445d233cf9a720a3ca1e16bab1115b93159862669ce686ea8bf7e3f29720f63bc0d0f23f2687a135b280b074b681ab0f2a12d30c2c40c2a55bd29d26cd1e2af499b1694eccd5cb3b8072f20078ea31c21c1c42ba6cc1590f0f087dc2ecf6d04092885940b8636a0fbee63ba9cf0693a03c752816d854aedb9f99b5fa72408bddd2265863025d58884cf6492d1d0953b99887901d8217b3473bd28bf1f3fd8df347e4cc66ccd22d17d4786ed0f67a4fdd03b97c76a645b580d5119811352760970b184d1d2bb107a781cfce0b5e39e21c7cef1e7bd2b9e4cba2ef62e7e55eb9adb169338152f28710694a37b00f6fc8891b08f32436f9943f19c0de7cfe3ed63f31a1e30eaf68ab68faa6726fdd02ee3f4772c6027782eefc49741dc378ab0795b227fbfcc5c5f07b1fe173ffa3a998a5a9ae2a09f8fb5625d60a1c5d498c3f8d9aae6f413133319dae5201a52f7a508db9f1a6005924ebb4a62623d287a2c6bc2a98dbcb83dfe4c8ffabab72e867c1bb21a34c6cb9db845976bd5096b88a72299c6bb11ffc04a6ff13629c61c82c5d60a597b3d4d397010201a42fed40c518ff30c24e2b8867aa67646395f010a1891df2f352bb91fe6dc99f89cd138b7d58a2ca6e7ba7ffe42b2ef12b1d5ce438fd48582a81b78cb60a87a20e0b9f1ab1d0f9db1f17c254f5d56ca148331a16e3e584ba9f1eed25e1ce20c5baf1d580e4981a1cb257a960968db93ca7674989e2a6c7b185a5c91101e9cebc8bc2dae876777250c0281e85edd9dd64bd1a3d93430d1008ed2363cd8a13b7e1c1de03793b0aefd3c0c4f5ddc1023ce54bad395cb93c35a6128479f5c5f3eabf3c4ed1479c47fc1b99c8474f565c125fd0dd20028976f87b83e5f9ed221efd5cc077ceae444448f40d08d9996d9ba9ef0d168c7cf984851bcd12837c28bc12c6730696cfdac53c5c925905bc2803ceb6cae4519b9faa9aa9db2485790e1c3b1ec10fe810d0c6dcc3a68dc93e3da7bb870126ed6f6cac361ad73331f065346143169184fa2d80fb37e28250dbbf6cbc99e324855e7f3f553c95b9221940e7de655385eb4eecb6080790ce09bd4e93c8a229509ad7d9f8e465116c1867d5c7d6f3985899e463791bb04301e9374b946d7e7851995db21396eb0e5d64dd772a3f4ee09e42de2fc773d9b9a251c5a515cf4aba0dc27b165afe018065b987bf9348a1016941756777871e12c816fba902f57fad7cbe068a5de0a380f72f2ff5ec4f594547172805369e42aeba13ff19e174801;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h276f813f2331d3133e2896875545f7c83023e2d90d715cfa794da79cdcc4d255bb392cd5e1019bcafbc7e5ed1d16e08226982e5624c7c1a840b9c2dc978cf3cee61d8f5d4ff3e3f369782797bfb507506f8961683eccad181faae3295f2dc8c75a497bf94b85625ac04305b6ccf246497ca6ea5df7e39944405d50fdf0e3de85d6961bf641734330f810beba5c81811b3086cdaadad25ede4e5ddcae19c0f15832458ede6e45b54ec7621bcb7edc46727068653f1a642332c28a0ee76bb0171681f534da2a81d9a5ce15f7827745ecb13e7ba2bac42711f171fdd3d51360a969e401abd9b55a3bddc0a066acccd6fc99ba15a3bfde49b5746c4a05cfc6e19e060d66b7506bfd762fd7490e943f6835ef7048ed466623ad82992a817e985c88c5264850962d698598c22051385020f9b44ef4307c93d1a7461f6a749dd7c9dde34b7d87fb3daa8fff0ad47f0d7233b27ce9a93adb71e0582194b99d3a0b92750736b6fff84295964e0899e3b0918273f6b6ce584de805f33735593ae07c088719a880db996e8089ac98db4de52936ca41d6d63bba59de7e1a92f25d269dcda4e99fc7a470fb6306d74aad28e95101049baf845b528844d4433d2c297e4e1ad7addc36ad358d5b494b6a55319ddbdc41049ecf9b006a46e2fd1928aba9f90792d578d00cfd77b69ff4ed7de3e67eedc2c8a2b044541171b32742843af2730baca51cff63175518c019a2c32dacc98a0fc95135d3c77d25b565b21ca6f4b026d48b831417a0c35af1c0a13cc654b962d90802ee8c90261be5026321231b3f606a950ed1892710029105e58eba0bf4248df85f08c19ac4d94deaad87132c948aa41bf0d22555de19f3efc2e7fbe819862eab3eb219baf0ddae26bd1817f5b6d7340d9d8669713c54e6c67ee27ca5e28eb0b66b4c0f77dc5c206ec28e2efd3147b9cc3a153729c2da777b440515b89f17e9afa24f5c4dae44136f25eeadb44489dd16d9eba63ccf4adfca26bbf9054dbac0f97d46374dc3ef2f7fd2faed8f37e4396c92b01d3a52c7770afc000fcc3d3b44e0942f9907be18f7a27d47258b8b37d9af3f206d4e9e24190830639ff39dc9cf5d7a82ed3200930117c1355f0ed64332c38e4dd7dba8fcf8b470e4a16cb5627d62dbbd060ec522085e70a762e4bdeea784a654b7bebf0585c9f7ac5afef1e70f5deb5ddcfdc69ce531ab49bb8005743772c87c26d1918054c84e64fb0822e5eb0b2359a0ba201ec5296aef858a94769553493f5393c8a0959773cc2ac2177e42a5ceee387a504a87de275982815ed9af1eb0367f9d4b2c7109953c0c792ceab4fad4454317bf6c22b8765cf131740c159d8c2c1b1c5b143c2ab4fd55a40261ffa5a42b352758878a6a1b7f26e5cc32f0e489730e5bba3ec23a6b89e03a6e1ccfd2822ff3f72c5c9ae35f306095cb6b418c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6b2fe100b8b70b46e6c04c30f31db5406658e0323d6717b853807a43ac539ce4226aafd06120c204e3beca2432fb6c7286b37615425e6c586765c4a89a1343059be623d12fa888db4c00969dbe0da9ab469eaddeed9beba9959da3a2fc66313a8b3cceeae0250f35dc17c6ba17fe3ae116bff33c5be756e14270f99fca3326522d5eefb8b204e9107fb5e36322797eeaafd2fcc0c1786d1cd0350793c8d1e1752996208017aeaaa4980eca5a6d98aee798d0fb19d94f6b65a92934a8fc4d26b834f8a1e2ac60ec87cfec25c634868dcb4d735ad76bdd12b1806c028719150271375eb25989fd9ef5ea597674931af69d22d437cb136fd70cdcdfa6cdf47cbb8f293d52f383550849d8bfd2c38fd33ea8de0243b1b752611aeaea3ea241eca9ccfe9cc467672cc9ad0cabe5099d978329dcc5e0858926965165d5aec93cce1022ca965883db9389570a79de75ec11f23f02b09d51b65334a8268e19f1c3885a934416a5afa0e0320ec261a0d3abf4ec466ff437b23297de1ae187f8efaef99c3e8fc2422f1d86d9f7af31f126a1b5cc1159c67d8b26a28356005b6162c9533a2dfe0534864fd1c45880b725b3196501588a8fab7e1c8ca88a3a0319c1e003f9a91dfbfe9f46c71f7ea1919ceaf91b93c00a053385936c16d792db637091ede14bbdd6f8daa57b4db16a35ab61b1843a59d8375a0d130b8e08bab5effe8514e044a711e2d40ed59f592c7d486ed554ee3214cbfcd130631a341df73edb6b45376745c1e5a476b24ef3422f8580146d7d0419124016654bcd28b875ec77d8468ac2d3e5db89338f4895b96f442a55088481c2628ef2c196dce91fb640418aabfa63cb0d7231515d61dca3f0d0f9dfef75152b3ac7d7e488e3c14bccac1ff1b26c16507b452a9a7085d6d81acc2e84c0530b026530dc814aef44c525dcb32b1af2c0cbc083a822c2803d1d64ed65c250dbd4f9aa392b6c4a61ddb01d755501bfd3c769c8d0b0c042c5e30aec8341da8013ccd9b95fd38a9fdd5159a0a289a5097d83362a890f56d2176509410501424ad26ac4a4b50e57490ec377661437e1bd604350fa6d9ab059023950ca36e31e7a725b2f8284c4e855c5b97b4bad4e68105fc0d121dec22c613283e8f1ee512fa224921eb6c44f4dfc947ba603810853629d1efafc4fb1c0bf13ecde6b0867e77a0bd92201a8f12a30917807c606c9d28689f775797547f01d7f4ee876c2e68b3b5fda6b880ac86ef16329d233475db03725cbf457aff49a6cf7f2df2154bb2becd09a3a21c27d53b377f4903149fab3c9b9783f80834d98769558c86000d287812eb3f30f2aef0aa09017d7e728a9ee862adfcab404340c295e4678f5e459039e5c4840113ab72f31e38e1b9d423f5df6ff9207ffd0021b4d4ed0f45a88e5ad8d9878dd893501dc203e494c510bad6c9d61f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf7c69a61ce9595a52751a64450309689845a53b4c46b4c3591c1953395c2ee6c3106e85a7e664bc93901def6902b5bdcc4957f73e170f2caff76aaf3daa94e23156223524de0ec785c95378ad9286a7bc47101b912e2395e6167293d3d0f58bf066d162765cdf68ec2211438d720468257dfafe0cbe29b07a99d1d2cf2340206fecd27bc175616961a18332d04782a696263e39846051c7bc53db8515daebf3abf2c71c8edaf2106073f2182421491509ff7892716c2d8c24f4a80ef5241b388314e8b605459af5dcea220ec7a665f81a2fa214d0fe6409bb11a63c782fff4068bd7578508314231fcf8578abd7a203138574a391520e3a17e5498f765a62a27fa37a8686586ed691f6fc36ea70d072fe31628c7babab7b3a723ce921bd7e788f4551142c1eaaf3c3562653426c56b93d985d7cd8a8858f01df332d598ccdb51a6f99cd3618696d1e4bbef9dc1dbea008424c7f824ec8db48f3e1b670d1c2864ebb8c525adee227b0485c96658c7593639e61867c897ab2d9cf7b171d2dc1815cb760c710060a5f401dba1ce7fe49063fe29f8453d1073bbccb9dc3fb077753c9a9f0133a490978cf51ad59223c6a870f21f58a176a6b0c4f9d1b6d1c7c8cd29ecc2bbc9cf1e13a34f230e7e5b4f52e2ac588cf247ac7d519510d08f6d5a201fe56c04c0879106251ed280c735f2ef10354d8cd95ae397f145e08abff5aad94fdd275e58d8e012c25f5b46bc00d6250d81e9f48e582c0c83ea9cb4d84f31b230fe5beb1d5a1cda5da38237f6801f2fe953d3b2037a6abf6f97376b7c4b4cc1c1a7ff5c0c60f881b9cbb2b44a6f0f827e7e5929732e652969b8faab55b599aeba91051f72b8f377180403d881077bc4f764e5f2cb3525d819ea1ee3db531d58022950fad02f1658fc52aaac90eb231d2370486a26334fa5ee3390b93b0ceb01b8022fd82e16c8444d1a19dd3533f37ff6bcb647d310db0ada967257bb9de457a0ba1401591ef797530f581f2e9a5cd4cb9fcc1563a52b86118964fd61edde8553334b890a931bb86e17bf8b87e5019bb4ff95b3a77dfdcdf2eda9ba105fa8db41fad5381ff7a29337b730c1a422ad39d2b657704463e06d0ec95dd08f20ed2fcfd77f3956634c750b6786032db2bd5f828f7ac7d38efb9edd4728567d389ef82d2ae886c66da1e28f2e79ef794305c58c0cd62c60b1b47e9596a597b145ed3c2c9e3257efbc4631e8315a95fdefbb533b54d62d477fe9b883db7eaa3d881cbf7a78474340285dd70d0a1d65f4fa1d53ca8793a94db0c02b34ad5f0d62eedadfb335655ef8529f12a7fbc92c6c9a260fdd4dea95496854b1728486a9a9f94e0efb1aecb89221b09a5e54b70eed4635c2625549ab7291a8d14cc7011930f09f2ebd6bd8fae81939f610c0b0c3e1354a4db1bd52e0b3a56b23f8e5cd85532fdc38c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf09ab022db1d98a23a3d5b6e0df03b2f5bd2f5f9c54557c27c8e0a6dc99064e53eb9ed961c80157ee6dfd577651e815f7a0cbbfc32f54616b176d3f6fba175cac9a81241eeb441eabec07b2a221a5cfa1fa3021de7ea71345b9431753fb6c30f5049c36e259de51a57c8fde82ec416927e51b5c32bbe41e7ffbd757637791e9e3c37fbcdf08914db293809d455b48b63a1de13aa92cb6b75c9e9a1e741f5ff42e3a1b9000637e135de867ec67baa5b49979036b343f732b959f65377d0da95bb9ddca095d95a0d83038a465b751b222ceb8e847a0976eedfea55f1b19cd113d6ad338528dd9d27d79fa2a2d2520de3104295f2f7c419da0eef5e91b2df127bc110960697c6ccdc058049b1b3f51c5d1bff78fbf763cd4fd16b99c2def00c338bc3c52f1e59a20306a0add240f79410adfe54454536ebbb9dcc0c8ac4df10955facbbc9ffef918246e63ac7855593a0c332a9de7f6a46ac390abfbd5bd9afd358048d44bc2f60c7fe32296a7fcc8144fd83c3a2561ac2fcadecc53fc19b4b63b846b7cd0dbd3305dd54c2a7197c2faf4bc6c90099d29c514b66ede55dc66c32e234b9a6242e2fe4980477ffe8c6365ed88b07c435d1f8800183521ab2f5ae8a58b75965829c92270e58ec216b07660eeb7d3e35472e8e4bdde74a475bcea2071399ea48aad72e2f4101e208a8f9d8ca01f0fb4d0b0aafc051f06e094b087471c11b9d6f0dffa57f81176c203ede8111c2e4d16d67f3b47c98155f753265d019391c38d61e7fbf3de0c15b7bd22873616ef4d20c1da1e2a2a8e7ab7a88c11a0d000e9aa2af562fe88216c19039f3097e39e3464d42344aef04fe98bc5076ccadd58afbeb9eb65c3f0483c8bae988b6870814b5cf3128a4d07214ff8a7e649c062bd9bfa1aa9ccef39b20d60e780788d8964acf8d5c2aa4879e4e449fe5e3e4a52c9734d791db5c646b8fba0c74320e8b3385a908cc06ba2d4335bb14f212f267119831a8d9cab2abe51f4778567059fa31fa4a3d1624fe400dfb0af6aeaebfcec4a45414e41d59085368c8d2213e07482cd83b41a9aa70d02bfff3244492c2f4677b1e0dab495d874ef7bd61e42c9bac18b2323844049ad9d70515cb6be5510ceb35d350739dca4e96d73bcadea46b1a5530e7a99b467f1adc55dd29f153a9a3cc62c6bda02fd3f102dc8b704fe821254d98f61975182476f81577fa37798238359c0de8238a07afba0002d75cb7509ea247c4f6d645d92cb28f3874ea87c2d4abbc640c38e1122f17b9f72f109d0d6bed331c6690447b6ea1ebcb8f0edc82ad32df85b60f6dd194888b808c173cb93530984437e840b1a66153bd17ff67c8c94a6f8a05606a4cb3be8fffac0f861a283286226aee236927727782231fdff9eee168cdb6fedc0b9a528754c2c4094448ec2f1a05e1146d566c1565a5032268142;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5c42b2d3c97ec0181c2817dad34cc1459b95993edd2a5dac38d05201801e82e9a4bc9b31f819ed337d4b42e0c769f3e268699797822930f46e3218b2baa40298a7e25e3a978e5b9efac039fffa18c9f0e41153d199f03e48849a4beae27cff34ff8aeca15b7677a81ef60377ccef87ee348e327accebe37d8c70af75c300522665aa74759c006bcc3fc28ff4a34aab4f3e9b7d01aad216090b7e52d24107baba0b15c5685a1f71b6982437837b259ec0944ebe477089b0ada0bf8573d40b39769104834b91ad234d7e7b36b30fb643192324a05de671544bb1f068786a8bd826c08e4b9d76172bc2c167a8be1349705a39f0d27ea2a0ee5562e78113402d656554673fb214ff36a12fc8f869cc0e5ea86cf40c0cc2b07f30afcc06a6a722f4ad6ed8944246ae71f8aa97fe88b60acc9504cb084bdc2357a8a48c7b41ac9bdf7c54fea43494b2a242be061bccc42c45957e81da481bcdbf2eab03c60af8f676d71adbd5a0ad37a4b6b5045e0c16a869834a397b970936afabb953e7b0e848cc73691f7e00190b17c1c3361d7ad0a739ed4c65b20354cbb92b90a7d0bc2836d6ef5312b614b20096d732e54e8bd74d45d5e604294ee76f91e8348c71d5e66654eb845c5e10ecd4d8e1d297014c21655a13fcf2532b5c821643935fce4f90c82b21db1c7ac3d3206fa81f39a6f074ac79b89e0f1432f2e9b4addf265e11abcf3f831c7aeb3a387cc66e92ca90f76ae218e24a64df8d87f27081d4cf78cbddca361cb27c06acab0086e89ae38278b4707104a65f3aab28f806298181301546d0507e898aa3faed726b71477fff27c1b9359eb81835e7a43e01c45963385173f3484de85a1fe56b6cdff54fdb0544a47554765a44386b234d2bf29856219232776e5b65a0a17af0b066cdeb4a0d44b42e9cceece7b6fe86385aa78c674a8ec74e664192a719f2ca0ddbb551510dced6b20ffa80371a1686d6cfab7e1714f9e2272ffae239b3c585dfc6b6ccfc68e4a8201c4ac26e1d4e3e5a346bc1caa60565dba55ee4f51602ed2f59b5eedfdfb71c4f0a0420af09c706fdcd32b49aa7d67f4363ebba3886e8d4f1bd42f3979919b24e8197463be02930bd177e23ee16556334326511da29fd39482ee150610d0a0134a7979edd318edf709d6dfce796a14200946baa8e0beddc8daf807bd6597b796067067207fbd1219ab2dad2579dd51b036c50b09446bec1d8cf701f78d7ee3f30329f5f0167c601485e1cd0da1e56778d133ac8385fa2a0e9a7e1331ea1262e5c12bd97419f0fd07b5516f44e20fd47929bcbe0cd99cbb65e12cc98cdeb8e458bbde83a5d569f7b3d1969962ccae1c9c222f78298ed7ab67cb6694d1cd30080b6a2bfca46a9f95c496a4502763ca786edb59cafaf880af7effa9c1103353c7c9045272f4df0a443d04c54fa8300858d829165;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3ae1c1dc717333ca3de1ccab8c678b921e9e2d75af06683a778e8586dd85f11a312bdee3195d12388e170058d290cd171ef9b68defa7a7a70ffdfcf16e79b0595494befa91c887f17aa5923c1814f4342e8d5d6ec0267a6708e5dcea1389d126592365b75037e0d557d317b110434a6ffa90ce004e195c1e01239c9acd4168109356e6f60c8ca7a5de19c4d971c555e1c145e921ef3b179cbfb8e111c6fa6f82c11e328dd0d1d823c7285f24357f437fb42909c148fd72548305065f7e66af40e48a4e68f38f3a1179abdda831f8da0973e621e78833ce3ae5b05799774b318823a7441aa558ce70adfba663e3eba4754c9f9d64fedf39fdcc122c69f3cee27a918b8895a86b9c0398b54dc08f55bdbbd72a55a3ae98011be58914214be5a7fdb626c4b9ceb8a5e2247a9da9e79deb19c60379148ad1cd90e8c6b3a7294b14e10cc1db52bb5bf8248b63e8ec7f1e2aed24ee10ccc633f278a146c6f95abfef83bcf9476813dd24b5a4fdc51eb3fcc3207a03fab2651a23071e7f8d584f1bad8b7de37a13ab5531928ed4cac7aa5f8cb7b164219d50e36f52ef32b9e0c91978241f03cf288ac823fb8b6ee2b7f5e695c9eca053d5eb9f13ad8c93683cc0760b772256e16025ae0fde3c7e56df1c14c9fe7031c82fcd9d0f7f296449ac36ee394d9421e2e380e4695ba8f37ac7fefdbcdc878dbdf66d4875b625f41a300094406e8768cf81ff53935c9d4600d90de28e48add82a4a7e2bf8c06218e125ee50c8050fe832d3c9efcdf6aca7b4314c46c448e79a378c9c4b8f32b6a2718320edb3aeddff5764fe220b9ecc665a6b36f25dba11ed69e8acb8517df8cd716ce645a355dbb04f342c225f5cc81c80bfcba4ddc237e8deb56c732a02b110c26e8ba653f5da09347f46da1b8e384ba97a5828c8c7c85cda826a8586b6ca53aaf618f98d6c7f55a27d8a84bdb2f3b9814e74d1a7b04506b4e11c1e23c89af0904703c0d7d84af0e89c11499ab67e018d4a4bc7ac586bb8c2d4913c2eccfc768aa1e51138c51b10f26b9a2f6897fec18f4a245f6236d6a48bf6340f126636090f2376081270a1fff4ab24fcc13297d503826b6f931ca8bec8a59ab8b16512fe813668dfe8ac83ada6c29b33313d39d00d66acb5bcf471d676232b0f1905ec769781d843e6a44827fe44fa85e501aa117321a4194c7fae0d87a2bae30173438d06d3ec80e1c851dd48f821b3ed6808f01f9e9aa01389ec146d4bf19e4a997f39ccab86d9b50f842782b87fe6c52b775173f4ed37d9b96b5236b9ee04926b189525a4dbf918c632e58df693fbd077d6a435500f2d7c5ab3e33c928dbab6b3d39a3f1e34ec1cf18b5e2386bcd7e6b258da68698200bfdd99fdc5106c5194709b92abc7860afa7eddf216709ccf39049084d26fb1570a54ff69c4b7ba60a0a369b4b8825ba56d10;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h36c23550c41a7c0c89c3e95154ac4f52faebad8d62c6d128d9b5ddc2346b1e213c4d436413bf2c3691e1cd4f6ebba443c15df916ac7b74da34425a930e377db60ce39bf094a9d3e3b5e34a735edd9b98c3e2f929e843ec090565f9b9a17d2e1dfae48a3eae814c62bd6515c5fa0932d1e081a5b9087f740d3623097fa18ce456c63f0335f314c72ab43f43283405cc62764a9905d883f99f5a80af04c28e8f4dd3e5112d18230c10e960642447dd4b5bffcd2843432d0c04fd401eb1c722491edb8eadcebd580d38f5a11d637376656a11a881c913b07cfbf36748b3a8a8ec43879d58153fb99150ef4b2ebb0c2bab5e05727e527655bf591a464095f1a9e47855935cc30f396618c898657e65eb816c72f036396451fe71d9c735e15d95f1a80b7dce26e0eb4c5ac91581d7105a18b387096e228b9cf4432cd2153d5417a0335d03908298976727972ccdea0e9f5d0ecd79508578a1edad67aee06190364a8912261ae2b099488494d813b41f2764fe4469d96f2bfe6eb18fdd5bd603d0d494fcb09b3e149e730876b03f49a791a07131adf944ed1023faff8a80d8cee66a1e61db0486242206880dcc98e164830e445fcfca01734233cf7ff9e102050d0b4b92d912505b6051e3e11084049b1798f941806202c277f1b845c0012375fee05b0a215364ff80411b22ca1f091e462697b61c00e310385c2c957422e0a8595f07702769b4c6da31b012b03af4601ce0a4827d8467a5ce670cdfc8981933be92879d74a0ee07a7a9050b8669ffd5e6934700fff683ece405715feb77aaa6baba28f103dc2b92beb18062893f73aa5745021322de268a6151d7fad0fd2026b4d197ec509526e95e3ceb353b16955be454b1ccf9329084e68acdece18a5cf1d2fe6247bee0ecda7505f4a00b94962e7175fe48d4e05b69c8ba2a98546adf9f92e217be2650d835a28c51f1352885acd2d882dbb7c9398e5e4a07bb80f5217a5377a6c7a057430a531f0fa3826935aea7ced2734ed29e3d93bbef814608bb8d775df3e13c83e727ce2fecd11650c77559940f292058f23a3b488454f8807712b261b81e6ee329e3fa63188a2d05114e7b3f07e29ec1239086e59171c165f094abc42cd0a790f59148858f35c7b81fbf4f209415eb639196a6574a1b2574419f44b2da1b7355884176ca90c71c96ef04f330f35b190aad832c98d9fecb4a29949356f039d1dc5e012cbfe218f7c98f89ca796017ebfa03a1fa112ed0afaf7b7a8f8d5dfb1db46e75ad74354c5cdbc69e500e188a5a5b59183a881af1184f853b9193c97acc5e83e47e7c4466841d026f1a18f440a79103cb63fc14cbfb3626af7d9eafd9610868f244d2638bceb78291fb678d384a803d1776a77aa798336dca46d84dce58964b723aeef6be03b11532011b22ce40b50a88cef06e46ed6d3c3ded2c64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'habede5ea074150bfaecb7bb3236ebcdc2be1612532c5da5b115cc86fc53e486233aa5e47311e2a89c5d77c3d7a5255ff823f5119d4b3c98341cedbee1864a1f51e1e368a5b62e2d6f5f238e9188853aef31fc93adfd606e2cf011b47d37959b70b108731627db2641165a49d255559c001815d78ac6b44bc32cecc42412e05154912aa81c52fb580353df9aa51f9662e680d17fa9f7268aed198baed8cb744fa0336f2b0a406b109e441a64c5f604a930d15f70e7b52c46c901f01e24c3be7ef4fd9dd58b2e5acf303da43404a01c057edc09b5ee8bd723c29ad14e583ca7b9846380a254e2b3ab7a005b4c3681ea5e8bb0c249c8131e87fae7b2f1ac87f747843b3bc3c075ed44b6ce5e09d4c3ead363c3cab192e73fea51515fe6cf1cabc62651abc22c830daa9b9cfbfcad032d45fc44996e02770e907d82843524d2b6b33d254bd511a027c8f7157be65c8983019025d3a3cf04cec8a43601918439e322a1a744314fa6cb194e3c77126a509d57bbb69d880e1f64413ba048ec4dc9408a1f2049f18b75e3381b526ad9c247e209f70d77a2eeb26145e4bd8929c61a2d05c691726b091b87b370f003bc927b37c59d3b6b29a23d651f4bae5fdb97e97ecae6ccb5df3d79fcba2b16fea476f071d25464f3ff66d1da5d7d0661a086e2d0586737322414eb7985014fa8b79f91920d6c83fad9c3147d7e1e751b932356be41a8d6afedf74fb819399c14ca59c2b834052fc0e0026e9d3993a52a8f9b96c2516b70df22cf70956884f9b7ee7ad3193a0d9111de3404f1fb99ea3a08990ac83b2c42632a9b0f687f1bee302d687979ac3f7839301182fdc2dd01205883471a7623d7b390c61394475076059ce1c0955940e79e537baa6e84fc5818073fe5bdac0a1b0a26de6b3cbe128f010c3f5b1f730fc524599eb8d60c3c8bea3dfaa160278d0f9e50614b14aec98d32b21b3b65c0e108f804c74b2958f06735195a8cff0aaad5f889da97586064e6d339cc7d3bf1bb093a661c1344efd4ea6e4bd1905157c7fa7b48a53200160a3e586a1a30ca129ec016ec8684ade86e041c7e48458bd6f2d7f356e0e47f5062dbc9a87e8e00305dbc9111d833e8f8cd2ac0fd2613bcf8cf50172878ba3ff8c56cf15142535e2709c3a933ffe19b9ee9f7d37f33b65dcc5cb3784f9b59f8ef0f9d486ced1eeeff4a4d31f2cc2feb15db0c2ae67bd07dfe9519cadd8c2ad74a5b8be9af41e7f0f5ec9ca4aeab8c7110332097ae266ee43eb6a8bbc72e020aa030eb50e2b85cd635a7ad3938551ca228d10a148ee000ff3cb4f5ff7828a4c6467a05dc4e1fad52c89c00ee320bb75ee3e3bb056a1e9d7c29762e9410bb3ec3054daedfe73a41a7f72e7f2861245fd4b819ecddda07334ad3d96e148a10561bf7fa3db9f1962bb4906d1ac734fc0f3d326c88414f7395fca18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8d1eebcdd3bd0baeb4a2fb2530b1f3e518e0c221f00ee2ece219c1eab5962406dfd5a02bf9741f449242c962e35ea7bcb8ac82343c83745aea3f375708c758faeec9648b516c98de3ddc99f577e9aa0d395f7a989162e752f48137bccdabd9d22be638793718061aec2bbef7ced163d123b742f659e6de17a053ffada224586fe3bf41a21afb66f2879085115a1156504a17a2dbeacb2fe402ca0941883bc8020eab30b38fb0c764f7f15e14c26cda4edbd31b9c1f45abed9c34fc7371d7e216de63c23d27f76a5c26672b4244d8c5dfa3366a1e9062ab37cae6aebf77fbf36f2311db36188ca29b4e9cfeb38fc1bf15041692229ed2960613987b72ccb9d8f621fe0770278a4af04794c2cf742902ea652d8e49c823f1f2ce84683960cda3f01630d296211b91fae3dceca31ba90013e75c5b2adebbe9dbc555f50647f11f26973c26ba82ce8b1f76ae73edac55db27bd1326c2aaa0d010bacabb843c98836141f9543e8bb6675fd5f64231b47f7406a743e7b59c6275e35f96fe5fa58a10ca0ad62c6110fa24869747581019fdc218791423075b315d76fc6c56c597d4cb47607597b9724a8715f3b12adbb8d9d90904db09ba151d1b34c88a46319d990250f8a13a95775aa82c64cdbfaf1b794d9120543d3e24ceda8fb5b3e16be30bf135983f4ea5c45b5ce1e75db119fae8e9c9025391145e32a25ef3beb7ad586b30367d93bccf361bcc3a308b9a953a2e75976488a7bfa30d77be42383acd478129c9553ceea8ffe8e77da9326c7850e035d4d43bf65929d284b97e46e094e9391e024c4228c96fff2099e030d64dde1a83f963bc0cd0a5fa781a8d3ea5428aada6cfcf1ac611e7e69c4adde9a80c5757c59d0dbba35cd303f7e62d8bc48a7776d1ce1cc173730d99b5424e65b30b452c7c5a57f5285568bd15cc46dc77211e00906785e202802ee54f137a63b99dffe79559f388c2f13a54813592bfd3dae0583398da3db360f617bd37ee9ee340e4ea7f4976911c7833df11201707b20ab185e9d7f2b7ec3b45a087cd110c4a40ea905fe98bde768f06e1d706b1c03af07be4728cc26ba879940ddf23bc19f381887d9ca1967f6fd3f2bf62c21640e29facd1850ed76fdff2f9e6d6a491988f30f5ec62e741756391269491389941fea3ff317064e407f204ded882f8d029a48ad6367936ae768095bb6a53d2a0454b609a2fdfdc81226ef502e1ac41091bc896bc4fb0e66e0d49e6808a6949753792bb973fc6d1640b7ca5b582187e809e649204e85039936867524f9689e4a6fbb01e6384129a9293c90c70b48a7a78b56c7573457047754eda4b24474aa5964020f5d8efd7d35792cd340585a7f1a0892ca9fe7b3436689d6f51c0db021484c7b94485a192b10ebd608fbd74e764e1b2d24b456f334339806fcaf1111816c09b033d50f66e4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc31a358ebcadda2da3117adf5d04b587cbacac5b86194baedfadb56a29ffc32ed05713ea5f5c5cee2713b9a246766cf9b36d9404e99fba3a99fa9af88804ffd03ae1b909e496a49dffb162a21c3031b50105997c740ff3e114c4e1f76006fd96ab6e9e1b1a12337c17aa539a781f287a96bffbbaf7f4e574fcf83a5ea1e03e23a8edafdf66311bd3c1c0eb1abef6431bd786833fd013429a73c2b37365d2094db9383f4741c9da9b4a73526c821bb6411a6a33f910896b95920520e9210c797b770a77f89ad72cb0dc25bd1281f16e81d688bc3afe854b4340b926c0dfa3f879cd3916eadf43deab5acf59b92f7deb84fce82a40f6fe073549e15e492dcf9910d8b8dbbba5bd9f8430bcb65622f033189ab70f3d5d91427cb1d238bb13dd29c1685e9632ff4e64db36bafb3fff5376a1c26c12922e3acf7658a187053de1d0c3741f517852760600359b705f1eb44f78086663b6764a8ce3b615a9c60e1007003d93ed885aaf9d9c8c5c8616e684c468ecfc2d986d81e35fb6a361417a1430818778c9f266ffc8876f5003cf895117a58cb3e8e273073c967dae75fabcafa22034125f072590aab9f56b145abff46fa1a7b2466f88fac4fa94c15f5ec01063b50f3ea03997203d0dd81642df67c494fe14031ca9105c10f0ac53529a1ffc2ad847ebdfb12b92577fdf0b6b7ba10d60c764c0a680347e499f91912e5d21290312141b8da5b2703fe2ce67e2a612d321bfe18e4c987e4fb30fcdc67e2f1d9311d11651a8f18ffcacae753fa36e17aab92f5556efdfe149db685dfb330fa7902bd414f5b888ed257606bcdf61af3ce26bcabd03487f9c3862f02f6ff05d2691c92bb5401eef7828e955397f29b9faeeece33e999db0d3e648f0ab6956c87017a4ea0d20e3cc4a7440a407b259de556a80a15df294642c14b1efc3ee5c42eac46535e3da861368cb5d5e6c0975fd5dec07fbd7d9b6e58cca81d49113ff70c39de9ed29ab52eeb72c4f66bd3e0b0fd89acf80964b4813d409bdca6e727c5c6bce53d1c344ff3c22abb70f5394d5948e196181b9490410b984f0a6d04b57782e378e4a593900779794b5f86426dc9b1899d4bffb78891d2f0d65020729add9dd8050c66591e3b67140de4ce93f3d19b080f3e57032ab7d6fba9a043ee7834fa97e71e571b2124593081069b923926b35714bbf1ef54b8b3576aba57d90e53ef1b4eb33f95dc6eedef3f1a9edabed9a671bab6bf67917b01d7fe9c2469a706d6944110d34822493ba958c9df9e3616947084aaf0f769e43a57afa24dd75b475c1663f097efc657094be48e09e425735778d1f3cd8ddff5f0127f1704e9f932e617a8e835f8754f05ca40e20ee0fce61ec42bbb0142fc47a5c77f25734f0c5f5792113eb4803f0f9b1135ccb38dc2a1f22c6836f4fb32fc3a878531f7a8a2b0dfe4706e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1ba4c01d0465515ecef3430cd64147e2004e65bf2080d51b5adb57db3719e3887002a9bcb2e9edb8cc1b0244ff03499f783240ec58b770c74f5ad7cfd0ce11f72d8a3077b8039c1f64eac7505de50a586b4d57e397f68fbae246505f88ad71b3fc1340990b7d7ca53d0fd41d9f077e64ee5af94aca4d225a6278b3ff0ff3d77f4a7a4871b7646d3182bb28f7e36109841707fca810e25a0062e07179f7edc62039ce3fce630285283caaf857ebd95b1b3ac55db59a40d5d7fcbdc02b3abb12d51cea7c2909f3aad3748700684ca4d862bbf0451e82af1066823fbe0545e61e2b3e137b1d5854d39dcc4821ecd335875ea6561dff3bfac1bd2c1afe9777adc72b99e068bf93a4eb8418cda69b9012136b39b9c63798d340eb6b62fb767690f1ce6cf745200e2806eaba3f58e07238df90ea0dad8c3f2c5da9526583bb5501914f7732efb7fb134b1ef9f693617b7441d166ccc5156a878905d3ee39f77d2cb64608de78efdef901b54576c6fa8d942931edc62edbca8da87f9a83b523a5949495cbf6cbd764b102ba25f1a9e4ad3149916ec8efa779ae1ba64eec3aedb8a63c986446eb6f732784fb388bbbfe16464dc5b5de81289781f4712fa9e964168cdc1f1f35ee747fcdc370592fe7dafbfcf31484ca03d7a6611473cbee3269f926354b6afc46e9d1af58714055f283bb02278b8b9df4445d10cac657de00765d8437b9c9be7a607c1c5b699df6e9aaee9657d796b7c312b9c235e0cff7bd2714ef75ea26fefd871b6293dbdd947e6f9a503edfcb0de0bc2067ab5dd50d2da98f09dceb877dd57432493a09283741dee8addc8fb53bfdd50d4d628522a44a682ba33654909bd515741a51adaecb908c279ecd708466213da9bc6768138c6959ec04343820ad96475d5060179ac889c509af91a50771fc9ee037995e36a49a1bb2d1b129ce831b12992bee44bf7232172528a960f3d2cdf54b6aea9b082b7fa2a8f3271dbc81b1345877edd5574d78d8971e346a8988dd529038781b44bfe15c6e6c70f503a33e52e1f1185309705565ab11b234fd1c4640e0914160198fb4fd883eddea94f0bf5251e729b3581536d1918401dffd45da4a79ee86ede03cb36997c546f93d175fd4a98c7710e1fae332cc3ca0321469f1bc63b9a33af60601eafc055381cc7c7a65f9ac7f1725725e1507cd881008955442674e9f28b2bd4f71936e599ffedb5f8ae52ab0d9e5d4ec06fc746ca7e04c842654e370cbb3866c163361762afabe7a62a646322d6f2806cf6d4a0d90c02fc35616ad8746ce404674e1462e3b4bd6c26176c152b5db586d9c08f914a59bbf1821b2bd094dcd38e72a844abb5e0a05704e9858be4b791bb9f6520618f9e772c01b55669429061de4639b9459c7e849ce1c2c4937bdcfc27c0f60fb1a87eb2c7d9b032ef0a9655d2f507cb226ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h63db01c5c0b55c58d4876e1f2107c8d55e255119faca8d48a1e844ce59018ddcd5b97fe6d01c250e8dec23b05b525727936f22a9a31c24f2d98383fc83e46ee12aabd51e6ccfe38037fce4393290b7d1a7c6c1435ef9a9b3ed0d0924f2cab93bf7e093ffa2f9a871aa5d92f3ea6e2dac112eb5eb4d7ab6e25e64fb1f39b816c01e00b7eb7fc419f1b4d0a523796d2ae5b59f23c404cadf20419d5ea5a6c756258119ba0670868f0bd76ed94ce01b3d52de47201cbfd1b6636f41eca2809904d28dbe065894b7c8fa995008a1a95336af850670b5bac7d86a346faac302e81f311f07a03fbb23d414f770cdf9ab47a9fdaee135afd767c4fb6c18811772559c0419d57d7e799800e67e20f3f1a1a4f0598abfa4fcf25c2958ebb2bd9e92918cc22e4daf8c00b6d7bcb72f0f32b22ec473a44c3681edd17d690900e21d72d1f6ae4761915bfbdbdf42593be842aa8ad5adb473c757213701966f160087a8e2198565f818c9fc63fc5189944765f0927cc67ac77a69a5a49037398a868e758242e7028895889cef789a958a6dde8fbd8301c0ab1f8ab9a53b5be6ca1e29d354e950e406e9de0682f8ec47c644831de00327130b156f37c12756684ebe4649800c512a74c1aad213b80801f09ed13bfbf61c9158da57681c6fa212033697560ba4aeb8dff3f4d4d386d66e160cbabed1980e8f488a180f20788b8450be37a39ebf26be4cfceef93a34235efcd1c9074372c7cab5c31b0024cdd827c1b28aed8e99e202ea8c421c2d21ab171eb1dfde174e33d2516557fef9ef0f9e6af4893e7e016d58004cf21c907b2ea32cfd566ee85063573bcecfdd9e266be8f1ba8815fb33fb16a47099c255e5e973ce84d10eb036a60a1f54a6e4031052b24731b08af8658373d2daf4ba40cbf31db534fba0d6a156caa9c43c6851c87d394ab950e6b3121e0cc8d1ecbf1247a3c5a0b6d9fcaf6b4794e88c8e35e8146e873d53b414291a4114eacaa02dbc5821a7f3fe2cba6f200732962bd6ef3ec3c54af389df9c33c31e2f06e9ea5cae1f2c0113fcf88905eeaee0f73cf3edcda8e18c605241846e4f71dc90fe940c8a73b19a9d5b5669e7f4ad0ba432e215994e1cb95072b0506a8fd4d8766647df132c4f346bcb0c0f7aa2f7104e5116482a20dfccb1eb2cd18e7471f84f581bd515b3747d18482fecb8df478f235de0184dfc682654070f3ae1d2ffc694971867f7bd2d4fd726fb6f04f37260790c6c82ecd914792b319869fb6636a41be216a6e77acd0cd43c42069083d6daf6cfc56c5c6ec211a0f726354e4d0372bb7982eaace8765aaaf3b5d088f815aae6bf285a1b5c926eba12adaaeca1f945af6680fa6615ae5c45974fe0577bef5dfb07f8f3635ea877c39a4b88061bd25899548f74576942c1c3d98905f2e4d0d38ccd0403c0104ade977cddfcbe6bbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he95d931851f21f764e462adf976ae171707d80c0dc63775611df2004498ad86c8387d55553b9095efb744e95151782d6886aac1bec6b320db955bc1965a6fb0d0ea27b4876388f76b82769b47b59bebe06f9507788d4e5e1c57e047f18446db088823fce6d892e4aec8fec73035a2637b24a893209fbf825ff154e19cb8790db9a10438ec51f0e2ae034fec0d8a73a549d9d381b15207b67acf9c66716a0ae1cab9e32cfb3c315e1d0405fdd8cd75b47970ba62d6f82f3570546fae1be441e2c6ed9e5585eaa1fdafcd309fcd834b5bed32a2aa73e94ccd10f3cf8f9d99de47ccbf659840e586a64217a6bc8511660f99d0b8451b077c802a5e88c4e21ea9b1a085ca6498a2556ba4d18f4e4e7698c775dc086b64c541c32854ce816afe7812adf5172ce97a6d171270c6d48339e0adeae1c9509c889ecb7d726e3acf7fa724582d6036ea05d6c164c8b7699da6de5765f65ade2e06f2d560c2e04d7f66c1a109c1eb05c0a6ac450b597cd036919ab04e583d4d3f40ffe80bf5f03b62fec953e8033b9848157b1bf7f3835358ace2959f567b57bf3a9269a2a65e623d49446924db2c1940aa029905187b7673d3bad6807c1a75a89539e7f2e5544ae4be746edc9abc4753af9a4b07eaaafd4df2da6767e6f7ac4aa8d0280936f782c67ebce9ff75d1f66d046885322537dc039316cc2d7bda372ed05cd1680ac4620a4addc0af9fb18d7ecd91d26b9334890a5c3bfa1e7009ffbf9534d008e8aae86a5630f387414d04e97979c270f24d23bc1d26958f8497540943f967ca8cfa4dc2d27cd5b9266fca9ae17f63a08542be4511e8b09297f7cc14c564a68707d4bf4306a7e74f55f1072fc94e92340ca5b15a715e840f6fc6e695d4d998d12d29c21a33dbe77df1bca90f0e599eba94308dc69254b59371f75c0dd5a7efd5a97cc155a3d7de43b7ad9cd838fb53a2cf83a49d12175b91c488c06475b8c6c962f9df5ad9247fd3af51514dcb969bad406cf3f7b1806b8e065b021e4679ac1d82ce72687a14967dd000ecedcab684ade9ce41719f59deb2f7ccd5bfeecafded47d351246805af854844a6ae37e59a8e4f6d7acce7fa913d6437b3e5d52b65cc84447b0f883d1ce30f232126afad0a04f7a4877ac11f4c1b1766cf690435746becf1c84a873138cdcf6006f6dea220fc77c1fb2f4383a9a719df7f7d46246d1475066ee85a98001a2a6757b2bb4c13e180aaacc74e4145b660eff284beff7120bc84035141c7cff514b2f899a679a59a1dbf0678be6bb19f13310349ab09c5bbfdd24feff3dd0c64471f92d84596bc56758f2ff11eb75b8794b7232584dbbecdb2b5766e9f47f4fa88d0dc7cbc0236c6c0979c51873448e2e783bf4822298f177a49701619116699f4f81f6f30701cef965cedce88f878468dbfd30d55a1378687e042cfce56b05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h79bbb4ed14ce1a5531fdc7dc3a36ef2f3447c5f209936142b479339fb2d89446053ffce5cfb020bc9ab19db880148305227ec38fd4bc3584e8d2bc4dfe761ab5e2b9bfbcf106ce4734c53685f8c136d451de2badafdc7a055ad025a752c3fe5a88f8499729f8c430a41425e8f3b6af92b0b5ec0f83fcde9ca779df3d2c888be03106216a5c9c7b8946421c5930cf5d5a406b9826ac0af06c922b52ba1ad26d62bc1a440205ab22f872ff5039285c7ff07b07b5a7dd012e6901cbc5a395efedc9ccd2d8e504ba98e228b84403abe67c683cfcc864809b73ee36d4c4766f554f20db9b7b14d0b0b2c5f928b406fcb2fcc6628c5572f6ef94ccd9913bdba06335a7c5dc23e815e4073e86fa0242e9cfbcd3c154e63effbad15124d99bb7811fdfae4ac208da0cd3b98d4e818e82b2a8d75aea2164f23aa9182d3de6f753b18a716bd99c448635b980f64c327c34560df05176c2fb664b5ab8d7a8294dc1dc5a2c37fc5c56e6bb46a19dac4f16d23e3c833ecd22d976ac4475876baaaf10bff6d18320e71ba5c95cfb763f11fc7348408b476745d4661f0bafcd7fd06b0387280f4eca0fb26d4f3b30e7bd02e139c145a9aca1de19b2644a00a6171a33a05574bd7bcbfa2d310ab1bf2e918ab702f0e19b45c7053abab423d55f547735811e9073e7048b08beff1398ba8511eb00b3afc4d54e2c980be32321bd2d4d63cb872f8c3fccf859d702a42c4f79ffe99b31b3a1c603f7c6a11a75ceb657c6dde834c027810e849475160340df8db23f6c2a22859ab53fd12f2a938a5d8b594e23e0e052e93a1b529c8d96637ff70fc0dffc1d5c326913d33d94424f48302d6eb61df29640216c9ccbd3d3f15c3db05a551a8c42f2775cccac89627f204ef25341e09d614bad8b894f2ea73af556b09f89c219dddb6d885950be58c1ac98f7b5eb5114ce79bcd7c9b785e2d4714f125fd80ccf937093e2c16d7a31c85dc5018bca3e27ccdd6cf1cf037a04fcb17417af330bef25bd5a952582e80d24d8711ab8eb51b0382a1d4eae9603a801c17db96d518226b4bd84ed8f41439fd73f776457f12b93067d1cd29c6656f985d0ef09c276bc21d04c72044f20863981fd0056d1f89106f482e9e4a7043cc3a5c26f93e4c7093830c1864ccfe880eec003de52eb0074a13ddae4559cdea63df2061c09a9834a81e94f44025edf6ffd83cdde477a760c7b9d117a6adc5ef985ab7a1f6d9285013642c7a4e20e64c905dc425420106a98dac06c5685dadf11e34a35e4d4cfde6d7ac3e5d666a527534a359417226a386d64d519482217061d954b0ea19e9aa740005cd55782e55d6b3ea9a2bf32b2eb08078a2a8ddb1b83c21579ace529e233f241993460fc238db432679bb405f394a3932dcdd06140e840777fa44befaeec20813473b1ad3017eecc80f78b9d4fb426723fc8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdb346fc26669a2cc5c45cc1adea253722d7fa50294f6e51c8b3154c735b93af7f5ab06e9c003e9e2f80437fee7e0f0bb6bcda3aee708b6fb508eca53d71520e002870b2018dc91a34eab0e758be97ee813a550e8426ac285d562172c76ab7e9c8c6b19d6c97349befef10367814d80d385d4d55730a8c2a4ba5886c8293450d694fa5fae2e21435ab7b8077b1f61b8345af75ee537a95f1e95c63e642eb65dc731243f7853d380dc7a3c164336daec193c3d5ccebfd40bdca3cd423cafcb32b1976181910f0b444672fb5a9701e01c9c667715872aeead548b95dc74f774a73b4cebdf35ef9597fe12b2afae1560fc1418d797fbfc8cc1c5a4791758437ac45be96c679bf8fdae5f66bb97fb020f0dd68144c96b84cb37cfd646dcdf351e3c41b19665a73a04cedea44a041b6759cd6521ef5cb1030013712aa5f6ceb8154fa528a5d66e91b8e346b5c4f8d9b364cf467facf4b0d0f41056c1777f9c2b87b59911cd8560257a5bdb1ad7681c590a540cf8080b7fb89a7dc158662949d32d4f54252440ba4ec610a5af4ab76fb14f4baa2e3965d36b9ea1cff4c4c78f12136d0e613b8ab07417cd9823bc4a51ef0c02122643c55efb7b67e0d98d5f0e707d4bd2de5f06b5145d9fdbaa3c12114ca5c104e91e889751aa003605f2163a16872a8558f6be52a8a67b24bf2630a0041093a1b88554cdc16c9bf14550a0e26bd979d9f3ae10562fa30abad99cf6b41bc6758534232ad52fb78ba31f456160e567d1d2331477ef44a4b658c945d4fec6574b6512ebc71097116ec32d130d65fd4494be4f8672051962dbb31e92f88b26152cef081a5b008fff42f4e7693448347a9712db2aa6b1703c950de7ec4a0ad248fddaefc5cc0dd90af05755ed90ed11aa5997ee182e5f958a9b4b023cb1dc8e831f7730b2d4e18b678ef050e900af72682e163fcfc3e6390a4285e5d0d9c13486bd19a0a8b458eab412f02d134da63556a01e71ddcbb7200e5540f5a577ee26472d2d320cf39594615e0d6da20316d5d2e4ff102409a996ac80d70a022f767d1e7fa2e57ef14c7c62d0fbee7688e8e4ab0e1dee4d78a694c89a5fa7c4a8a71d6106f08b98610bdd4431efac8be909ba1fe7b1fe40d65be4c3a30d9d72f7cd5dfb51e2c69e848eeda9b2d3d1e55fd9fc03dd0ff45db62cb00de48cb5a8d2b4e7a1769ff7c6f9b8a6957c67c6478f710cc5ba07da3e41fe5ab4596cdbbc4a25b6d627161b8be181b44c57d1c5da2d8ce311643905fd77d3bc43b8a1be8a57e77564d94cba516904135e54f69e0be9d82b8c868db5c59de4f13f0436092b0c39b28ff6963ea9b13edc9e51846450320d5aa5a6509fd803decc9246ec71a05f9b1dc7f90ebb611aa28a6d159a8250acbaaa11643695a2eae3c5531600374fe67fcd498d858d00d682ce739e87488ac98a5fe5c3a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h778e1058594e451e0a7d067507c32953cdede7fa308cd7ffd43323de3522de41b08be62e1216880f8657c1ce0a98dd72c8ae44c48c4b96ea6c956106fa2667ebd937b46e41e390b53796f3aea36ed33688f038556c10fb2722c6548e8fec6054a6d023294f4262c0f25995806093cee1e5a52ce517c0ca818f4c9d7b0eb56084819f91e6c6a3f8d6c47c92d5af76168742dce203f31ef60b5f4d225d5aa52675dcd0ad42ec8138f36d8f43eda8af1fa073a7c16aed4cf3cbcf4aa3e5e9aa1f30ace152521fe259dcccab9ca293c763100e8a0ded1c46f8b3be0e968787d13f1a934793863b1e3463c78390371b56b7051aa3e8314cdebc720b2ae5465b7688db2926c5770ceec75693eb8b65449fe1664e0560c0a609026d9ecd4553da564633226a18a629e5a1c966ec3ac7cea46639d52d730f8ec12c102638ef6672588dd5effb8fb084e8d66896ac500c34210455afde6a17b648a1dfb2470cad2280c7c17694ce81c1354c02340da236ad6d516babe0ae05bb0b60f74e726286976aa34e199cda7caa39a6604f7935fe2c0f1077149e4312bdbce0345726eea15b390e8b6d2fd8d8636c13670a3c008d5757383352b3d8164ba404f975dd16ea27ecf9e4b42d17ae514608144e9c03051a1a6926ea6c9b3f37faafdefe1aee022cbfd7de70ff2b515005ac4a53569301e9766249e67a1530df5e8388b19ee4c43f4cea3a08e8a78ee25fba3301dd7bacc886aba28fca66066ef475a271826a5e1f7edf81d02f0fe0c8a300234545266cfc43440bbc1a2ebae5ee174281837e2637a6a615cb5a486e354d5c3f798058f1eddf8dff1622312f8fc1f89d9f679f6fb2832ec18e9187e9f63e61498534f22dc922a33e6c9bacc68798d695f9b17898c8a06163952bc64f17821e699eb43593db847abba4d69c3cc39600c18e3f2fe57a2251fc4e34e7474ab9e71e28ca2508f52931a7444b69fddb1e2d28982c62b77643c825a97d0a450e18949ea998241246e76102b06c493d7c2316db9333b8ccb070cf397f0054ca57438d8896971f056f40d9f9893e13c7e628ada4623d8530c704f54a1d94372bc79fb7e5b66cdb308976274e28c9439c053ebfe1701fe0590e8a08913a99e4e339dae4b4f17ffb160020e02c657f5249c384ad13272a0a314f1ec05cd9de0c69b3b148b5bf5c0ff1c62810723446765822fcb32be2d183be6dcd21bd030701eef81fd2c85be8536e618519aae82b7bbe02b0258cb8ee7a0a425695c7c868e211d6c6629cc71db4d9d2318ea4031785180c39173f9a3c91933038186ee8608ea92cb0405e2161bab2a4119c679f5ad71702546088448ad34c8ae157d790c27807c7ef50995f263942fc4c070697926c6e46c9851bd6824db35f72ad4f4464eca63409719334806c9d9e725643a3473a9dc205a8bf3fa8af4154c58629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h68bf302a9f3ee329ecea66b156fd01b7bbc9f82bc94b5ac80572e74c84e78dd107402893bb778dd9f16659d8210be52b75455c5b2ddf395cf8f1ebeb02f8dcc27bbcd9a1f57f6f13d54a51d95d08ee08c79720502881bb891b02881105db8879468425ffac6fac77fc21c22008c6e05e37489aba98874e8800fdbd9b8e7af60df438be272e0f350d5c22cb09a2aa5bce8dc89bca0b72e38ffd3baa82f28a440c73b806d245f9d429cc616553603cc9b9b83008c3ad340ea2d3d8562d91de98d41ff6fe1a0bf089de070d02179e1718368fc4a0019b3960caf72e5f1cd382faa60862c66358f262d109472ae218d664327a028985684243b786ca2e8b3b1911d544f312c9e341ff6cfcb3ed7f6f8efdcd81c2d8ba40be2db7cf080b97150ac470a0868db5ebef5a9ffe85f6397170d19413273f7f0e2a3e3d8e180803f224b2accf31625cd87eaa656bb164160c840443983b8bddeb364330bebea3742476fa520cc966b0bf4dc5a8c91a766fde513f1103b7abcca5aae911bb8f83774dab93b2dc3207cb66f00ee7ea930a4c5d859890f0dea73c0e9ad8f0d748e45db4d90b25f9d69e9c6d13a4862f8ac1742285fcef4669cc57d6240132d72b561c0666d42a0c2b5ab886e8e70e415fbb200821b23de1c9b4dc886d2ae7119cf68d1075746c38b1673ba8c56aa5b9fdc583d2eee512293fffd0cfe5c93161b372dcdadd58c1b37e642bb51ba6e048cecde32ece2ac474623d59ea6b8cc815218e3843ef79fa9a0b87ecec3d1ef0ddf51469787dd930b918c9cc1877c20d3235dd2c272d3931e1f87ff7b87afe148d2134fbfdc43c7f706c1d538a368801165858221d2004a9a15eed2cb91fe1f549a471daf2b8b2e045c188ea140edabafc4df9a8781c819ce57bc1f4cdde91a53a07f25361ef62e9157d27d9178d4f1db26da00c3afe9d7fe132b5eeccb3faaded536981cfc7d077a83c4a0ef70de3aae81f456a60442074d69528b09b799fa36aa4d54590afa8bb846e70debf50d393644439556d70a49eac088a8b68404043f3514da3508af40769a55b3095fef4ae7c63cd050f59f47919b36c010daf53eda880c2cd115b76914f74562dc7d4a622403f12757a6a135d4803a70c6adebd913f2e264d10c9ad533dc2543467570963c3621c7052d13176ad5f15537c91184f218d7857f8397b4ccf03bcd50e70585f14342356655541735f947518092fca6fec7b655532045ae0650a44efea0dc1fed07768d9019a1783f0ab5c29e192a2c3b0721ecb4c69361744f71555f5713d18285f5f44f366002b87e2bcfaa5d590b5d8c0a30abe828abade644816553857be5522ef5f1a35ab622fe10f3988d5dee8c7a1070a02e6a818d7f5de6940638b6e3761cb487329e52d5f194f4273144b5c3c9bd9d30426f2d14f7ba22d7c619b9f29acf8782656f271;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9e0ec691af88809db5538bc6232e20bcd79ca49dd18cb8c49e7890c834be51b4d22fd71b11503a6ea1b1974cce93656a580902668cf40208be4ffc823083c588d3cd6d97de3508b89a4f8c4a531deccd5a45dab4595cfe9dfeb175d8fb169d76813fad09b4f441771bd5421c1e82233c32e1dd3755a3120f19e91248c75fa42f0fdda3aaf54ac05560c82724323fae9468ae24bd87bec8492c03959828e7d0bdd1ce93ae97edd78ff3bf0644e395d2a4bac850dc01095d155ae96afe1174d27c7bcbce888b0c7be3e82dc4bead218572610d8f534ee7f9541112c07a308ee6b91f745e4b2dd47640dab269b5cc18a72784c084b8c16ffb33aa2671f37e45f6a0f81aaafb3db6fbb81bfe1732d75ba6c1ae4cce6ad357d3f6ee4ac45cc0d8769d5028d10eed64ebfb1ebcb78b291b64fb2ee5e088288edec74069b5bdd351f65b35914a22acfb2f071a2384c59d4d06b6f94a74208f2df3f3049deb57e935c79164e909fdd7f05bf1038501fd012118efa3ed87a4864e294907d8dbdbafed990595a976f4f546cd3fc0ab4e354065d9134968b71306222bdb708d8779707b306fe74b8c3b6a2381ad78974dc2ac1d6fbdbfecca8ae7e47430d4eb835907ae76022232d3f6411fca564405b1da2e4241d2c5c804c04ca705e1b13a7e30a2e9daa7ef0ce4bf3f2e158fb0d87968533445c65769fb834066afb79ac2f15a72b0e72aca929ec7263735e2a9a9b468ee8df717d5abb87abcf1d2259f78f39c31c4e6c64bea4d2c6c05601b9692e5ca21a73c8eebdbbe6587dba96abbc42e48e4ae4318106bd558a88410bbdc37a471b210aa4abf0885c6088fc141706ca0e728427396c8368a224d7e5fcd1ba772634181b7522490fc00606a9e5fb54205f5614f02dd2b636b9d5bdeb2c7b816f833d588c96ba22a063937bbb7f2c43e7b0f4fb7fb696779f700d9dd87be622ef53b542917c8fcaacfa452979d9c38259453ef4770e25ab9661a0799a6b770816200e000121829adde1c716963af5fd8564cbdd1498e67e1d3ec86ba82fe570855aa2cdb19fcffbc7b75e4ad7da633be21e96aea216309d5f65a7a5503fb384246ee0b8ef44c851fadbb2c3fcd25e9a48951141bea7df01f8047847a216db363210870793e77aff7d2ae56a1813f25d6bd95a0cb17eed5474e9ba3090d61a94a7515dbf7f87c4bb7c95fa966a58bec4ed0061c33b7656fb2a307c2533f9b9f5de92b5a12744d53b3781d71df45530195beaa150641c23fa4873548843ff87a02ada9f8a6a417ead5136c242e8329c2551d7981f7d22389966cc9bea22b2e6127eeca3ad0d078924682a3d3ab70a12da55c480dac103cc2e416f5f8c394ab855c292bb7a603c308d8342d78b678036acf39652e84d64fc2c64e5d602a10c0606cd36d8d40300e5b46587b10f8e2ac0152356acfb68aef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbbab0fdaefa10d608d4b32f805e5f02d22038c67de2079717232b09117c0fa592a11c1cfd16087564a7f5b50a3304fd1cccd536e198c9dc18a966de92ca7baa289cedff0cc71e8b848d57955d074622308a88eb0a41470d462fac643f87dd7ad16ed8de91f0bac5e0c37f1e5066df60799fe1414bb59a86d3f479fe5c0c0789ae1cf894fc97de770b5686bc30007f740619d5a09f20a2266e972679f1e3156d555800f910b30e75519d02408b9c4771f12dd5d95c482fe8587d31494eab5c1ec7e597c510eb713d1ffff8c3bd028658ccb90144dbd8acd5e90e09ed2b3c36573c67044d813c0de3de3b2426e1fa97079160a47973b2ba55b0e606b313724bcbef2ffa4163fd9e558365ea2eb67c3f09efb754a60ffd2e902a813700ff8ef02291b8f837ebed1777653d6e33fd17bbcf8cd2b475b8a4a4d5980ae4edb72113b586ab9b8c3edaed7bae4511e4af8ea769b99887ad716cf1eb088d48dd5b4eccc6111b430fe9c6299a23336eeb7e62c23e05f12e4144d5eda532a4b11dbc77e99130a5b2617895e2f6bcb389e3ca83d0d1dda00fe9da45361f5a79375d019f86f219ca818cea882ed797df2af39da8e8c7b13aee8219db32faa2869724cc4bd60d78f955e51885632f483f400202c90a31580f1dbd69e86c372c4427901e57d6c062a79c1d0f98402c93d3b1fe5dd4efa314b52dce6caa51298d9fe3e013f71514d29371dff0e2475181893afa66013276abc7f439341bb95202fb2862c7cca30e913bcf3e7d048a9a382d55663ed2bbba96b560d6b5e4ccc306eebbf3d7b2f9613f1a19aca1b7ff2fda25e3cfb16e4160ebbdb7d2089b843d2878212a2d70fba394d655b02b984cb97d1fa9c317b9aaad5937bcb525c64e3e5ab5ba34b811e915e49f1d524949ba03757ac068cb292c0c63258013635a6a18aa9d77cacbd4b43ba61c3942337f4e4d6d7f038a098953d66a4fe0f7f11c5e9ca98aa09d4a618097a3774532facd8b3f61e2be43901d0501fadb5c837193d5dca53245baef0c7958a496ed4210870a19f4dab2dd875501b32a6456dfd8c97608e79f48703583cd81b4b7173a0f1ec33c1783893a62c910dc7e596ed8350ed0eec353c07ebcc3743143138161934ce278a6fb4de05a934a9e38a6d77e80db5d26864f9de4551a3e69aabc7fe4de04c2df651b76bd90c302ec97ac3663272e1f708f0903d981f4556963565694090c670a2ae5d9485215ba5584d15dca69359e8317442dbf7e7eb5e47c03fbc618ae07375d751844a75aabd14e379799a9864837699712f9bbe4a95eacd52b7b9ce836c5f507799ddc3b56c3da1c581b948aaca6b913bd8ca2ad6816344cffe7c2bde1bf377074c765b948b89a3c67c125b3e3d46c525e3e7a677308a9c0587e047a2ad3ddc9c8cb7b1e09f1f84b619b44a76be0f6fba0558e249e46c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcb8776220a752b50862d8e4fbe789562e298c909192f9ceedec7f5222d535c00bbd657366445138fdd77626bfb3d0b0f0655435d41db23b3ff5d0958706174c3dfbd809f36742da04343ddfdacac3209a1f901dba7916b4900fc2712993f7c020d7ff9691c666798b90fec1cb142718a3144449c35a2b3ae3317ab3c5476c4324d936c1b9a35c7fa83718d1092743b6416e078d355bf05b2b03b6844a03d839a313f1f8707a11ffde651bb362d1d4948b0be6f18315367f0e5ba4531c0a0aab1698cafaa0bcb5220b1c2d554e577fe9e131c419ae4dc0999689624b9eb92ef56e543e7a4c11a74e8513ef95eb0f677d2bc53faccb03f871fa4ce6eeb25371b5b4aa906d8c7c2822ea0c5b188b0617582ab5cc5af9cd33195fe2058cba4b90dc34dc3b3474095df290df52fcc82f0b467d4d3f4a3cb28b80200ab835841c7fc0ec8c5d0aacc90cf094279dd6a13e24fb91b75176f392cab674b456beb80c5ac86e3e8732a75725e601b92bae00fb3b436dc222095e6681000aac1cc9950a94b24d894e210491c4f539dba6e17f0577fe3939fbdc68b4ad16835aab9de5f9c67e045b4322ad9901a3c82bbf446e8964d328a19fe0281914753c7b75837f8cd3805a8353aca290fd5335531507efa7dba71f43c8e02256df940a9db349a3c624cca016a774aa246a969f41e94c16239cde5735714d499b7cffa748fd046cf42806cd0f336a466f3c26b9d90bcd2451fd2cf67d025a86faf11a66c7b9b404aa0af12908ca7ce7a2add25ba223c12302bf680e65a8b25a93ca21d7e98a1aeddeffd2bbcd8c502eb6652e54787a8532da7e110ab342afd7212346db5ff2f35459a0c5ed6c2fb6ff5b2cbb01f5462307b97fd5609dd6d8dd2910359900bc65f0910905b22bfe8f9ba99efe17e50422d892986cf9167c94d2e4cf0d556c739e0db7a2ea1a2b22b9dc18e7d59e32357dc17e9e28285b4137bc38c1e27bb85e368891bf43e28fc1579ec5b4f2390f5a122b700a235b9fce3c34f3599b5533e388185102265302d821d3dbd9594c6e8a0b47d6b828e4ba67f1f0dcb4bdb8c630862a561be3b8283c4c005df0619b825397a31c78bdf6413679089a9c02b225f41d3e475ef4260be22fb1bc30e342cb90d2a7bbb1637c53797cfd0f3807a9dd27459f864e0cc22426446ca987b2e8bb5aac6b9602226063f0fb93ba42015e20708b6b08eccfe8b6959ac338735221eb3f0e60dd687bfcef36017fd9b73e2cb264edc93c543a589671ca9dfcb5ed0a62e83598ae13f8758dadb569e16a99153f0ab2f2027a1c11dcd2fcc0349ce375157fe4340c1ef9995285b7f1a24bc7dd066c1414326a222be76218a47ba10486f81551a81399a9110789a74f2c21e22e515d50108b2a6c5c5c9fbc900fc8955dc3cb2974b5b6890fdc5696c4b5989c3ab3fd3b5eaa384b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f1491d2d66f5bed0aef8a8f9bddc94b538283b0b89ef2d78db3c585c27c2f4256bdd1488bac3ac179de370df2bd144ed311bba30bfa88038623fcc031d10f1c79e2e81381e35e8d27900b9fb0cac30475e3d3e1e3eb77258df72a33aaae73a046d2ddb536a42a3e37d64b0961f677cef5c3b2da9ecebf7e94eae7a8d5d40259a70de94f36dcfd528ab1d60fc04da827f148aad7b8d7c3383610e2b2540140132dd21f131f0d445f15ce51b5acc1209c1f7fea5dd1c9b29d3013b7509542567eac1386e4619a96d28c4e2d3303ae3f20d255420a6daf3f4dc90e225e65ef7e9729a1c318f55f7b0dfbd6d2c67ab660873ef51c03edc0c031298a7d16fa0ce7ec5cd21bcd7edd68352facfe0e51693e3489f91618193e9d145b6a91cdbcbdc0bdb3c40e8e8469982524240ce5cd2b0a0ebfc7326d1beffc0c2bace7cbe000db886898f94d67392d22ab22db11bf9908610c90b6b037552b415ddd4cda60fdb0ff237b6a4238efb64139f248eec2d48207f106dbef6b31fee69b5c33dd0891ee29f6af30709eb11391f240784731eb0008a437ad63e25c78b7b340d855d447a9e7677f75130b467e5fb250a1fc27e6d233cbcfe5ea575a9ba22fdbc44f11db879f93b6fbc60ebd1d57d44a46b825435afb56d61473e0d9af32203c9aefb0b95ff4ed3c35e71a6deda184946d5c01d026cb2c343fc85e27c5dc33f5df88f095699f372ce36a75adf83cb80306208391eac56cf0494774eef322d0590bd9f5a3787557d18f3c15c83f5fcd88292cd683e1b1871b6d801264443e34770c5c6f82f92c182cb191c5ff84add0d86e3f7bdb8041953fa4a9235d4053122e0ce9adf98e3850c17b122c823cc35b795f31c9a320dbb2ac41f4085e788bf93787c968d7649f155f395a7d2446458262a29889f67d088972467f340b112fa5fbf278bef15605079818426cb313043374af6b1d286187d79d323f016233ed42edaa7b5300b7c0a09af245a105862efbb066e69e503ff4a76c4baf834b713799e32a24d34b18c742c68ade59500885e7b611a09829d981e83a86be63d150e7975cab8b993c7d4f9ca253aeb9d902af209f034720ac29219842f1c64dd092056b2bcc23a5e9d391fc8ebdbd68638ba402eb92360b0f730ed7caa255a1380c96df2b6226ca0f18ebd14ae412fbf6c5838319d036209ac8b7029fba98f6674cd2ebac618ad6dcdb470a9b49a19b20a7b7504151000982ba7d6734c6632a0e522b4f64546d5f78cb412099ed82486c97dd918695fe33a06739d7f9b3d0f63fd456a40693e54262062230ca7db8d1de5dd7bddde2d37e20d15dd60e367d0df19c02d14e04b9ffe1ed33797ee02266347fc098d8d343bc6f378a68b8f0e21e417545647da44754d911b939ca2eb2681eb60b9d1d4ccbb7e495aeb639ee8613d8182f8278a3e93ba0f67e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hebd4533405261264a4c8dbde2dd22a37dff3095d4c691f1fa4f33c06caf66ce9ec80a8ecfdafee27e4a7ee3b6d38dae8ddaf3e1330bcfe90b459e0f2398c76775cb12c9c02ebf4a9c1390b511ae688c63c2367847fe542dd07aa7afb6865976a02ddddef53598af8ed03c2766e579410e2bfa9e399f04a4fd89adfe8ff87e9d7276bead98db922eec601780d7ede6ced484420ae0207bb47ad433b58763e99c2fc7ae265d7b0c01ac41e5a7b58c86d172eedd2f07a7366db6c5eeea219950b7aec4df1b8ac97e36564ad93397680431b07dfac5267bf95074f8f0fde136c8640087f12ef6e44bcaf3ef94bd458f4f32626289c75ec8a7795cfa675bb13cbaa4a1f61572ee0a3c67fedfbdac358375ccd5562946a086babe78b95e836ff47bf2f88d8ffa68b4b9025d7831d62a03aece8a819a775ba1d099baac23b0450e51d7248c4e55ee4cbf28b368d3a7e11e708f89c48890f5fb646c1bcc50206f21e5f0224432314d6f42b4eb48b731aaecefeefb1dc4420655040350c24bcf4e5c18b5957716f1734d47ea28c46483a4cc0cb25feefa8edc26a8e4ab6db325a2d4edf07a55b887e9169e76b3d5360cb72eaf4aff1423694661a9314106a932bc7921b1223d49730f7e42a80c0bc1920963ce10cbc6db33ebc87ad26a24bcf24dca8557afa8c1718fcb5d565807ee2678a49f902df7bdda5e35862b9aee065a47b169d70aac9761b2edc7057d9dbdc72ccbc5e114a3d2dd9730a191ec74fc58971dd4bc684055ff8e3851d01cb937ec3648fbc2bc7e486955119d162e1daecb5063fe226b793a50cecdb451a44b4ad643895c1340660df228ebc9bc43e8f1a4c107d8af9de50c3473a3f73182eb96a595e63117a8aba331461211470ed6d648d0d41095c480902d1b0cacac74dd3e2bb68cf0b0e732a7bc9f8ededf053ec21f3f05347123f6c623b49495d6195ec44bbb66a419e59a726090848cfabb45096847354d52a0dc2e480a7f12ddb32a09db080f6bde9017f1c3f5c311205e023ebebe87d96fb17fea537782df1f9f9302171e5ebeaad3b1afde5d85be11e44e9f437d6942c953fa615fde5274f954c1a3b993e68873d1af9518b8e883e4fa7e6ae45d297d6c23e73f9018b7b92e93c70ee21e44ee2eafbb6a817a0feb09ad9d80d813c11ab9a4e63a9f73dc76564517c02f019baf3223fe64c62f31ae6d7e7fa490070a7ea0007a0e00423e6c94f14ec74bf590001a0422b6dc77f8d763341d96aa9eefbb60df3dcbf872a109003ea99df0da44bd8566b3f28bb3166a0cc5824831cdc521fcdfffb67c6ba91f3ef31842ea603281af41f6fb164141854ba915a691a31794702f8d6ea48acef4ad95e142c50a567bd2c931d4ada133cfcd7da25943633a1bf7f02a8f6c34687180bd866b5d50e0adb1f21598c23328388714433d931506886be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6e5498fb01ad0245a824ffe1de67fda2c35921078ba1dd2f5aee3c446980413de3edd9ea45d6acbc998f5317dce62945bd5ea3a8a37b0add5a833541d76709ae05517744e92dc8fef87893e21ce8caee22df9f726d4710a2f4e213eb6a762c6cfbc8e69ee767d15fd20686dd2bc23ebaccb4388ffec593774d97aa62e7aa4c85073a95298f60732103421a9f8055199cae4d817b1f6dacb7c7bd497c99fa8cd5823d8c85a2bb3a52c76baaca9d53400f6a300b0098ebeffa443ab83bc113ac096972b7974d0f8f4da7ccca086d958b0a9d068e1666f2a34dceaf71bd2d359d05ad2ef8db178eb99deb7c1d94cdf776ab97db49269e3916a910ba3d1a232a595961169957cd1d39c7a525ab256e6292391103fec4c80a83f80fc66a4b8c4fbd7d723a74116f4fa74c5842a2fe2124ed0e70d42965f475e8bf9291bbdec51cc6e21c3753d05f13b329476747d6a6a0edd11a9f076b9d55676c6fea0809f028d9560001e32fda6911a596e38891775bdcfcb78e191dd3c10a0b9d33deae78b5f7ea9f1041e9442bbf064570cd252a7e46a080a3ac60e9cce12878f97a1f19265e06ca6bc49ade64eb9f57b4fd6d719be8a016aaa8163243ef4a42bb6985f597fe165a2cc30feb0bd00f43f604f5696b58c9cabdeb90c6bc32efe82e3e7212e396adb0ba0f6e8f3f247d348dee83a844ccf39d750068deb31e026d80dc2e1f714875dac67f69b4d75e07e532230e769edb16fb9e4f0ea649f659437e0742bf672c8103d1bef379c421b1112561c0c8a59e9e500b767636b0f0a45b259907cde98e5ba66e3a21ebdaec1f198f78656e56216c185a3371bb1685538745c316e420c7b1d67c65bdd01c675b63bfc5bfffaa8df6fbee18e023b203913bf0bfd5b17c8dc6262b0c434a9f637eac6b88349878f94d40d37ae1b4780873bcd2d17c006858b80ebfbca9f54d658e6e61dbc102aab2dfce9a83c8fff7df0bc0301d51e178bbbf0e5ebc65c3a47d76c00424886427907b909ad53edbc4c63331aebc0a450376fff8f9c8874f693c514fe3017c3494c2f5ac53a06e4129a47c3a36417e338818cdd81dc09c71bf3b08385b356d8e92a01fbc2fbb0f25a2dcb4c4649ed22ad76e6ce909ec1965059930b3b992d265f214bd1d8785431ab38e71ed770abfee20fb343cf8a733044b9dbe561e7b803a8ad35619be6da9d8f861da38a7f2ddb1a98c4f0c8ac481a7a88d8149fe3936b2dfab58c67eb2603f1b1856445267a3b47ff2a8382bf3c6ba225f6bd89624b34c8ff18479243bbf5e12ea97258eddfac2b7568044ac9bab12a04cd69f124e8202c8d4292e36281fe3cf68afe059ab3e6ca9a7b89367aeaf12367bed44ab31e9802197a67842ceab7076bd7b1bb66d2d7904193d0a11fd75577c955a13b02d7f01677a92bca3fc4aa14ba8df5069562534d9392d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he9532628c380f20cd9eee4490b5e43a6a7ac3a7793bf6ed4d2611ad46fe878a9e76fde4197d0036f34d2b7e78f46e86e115bb64379c26390964765074e5578df00337e658500238cfc7c0621aaa3dc9dcdb1cf74535e90e8487ee6e226425d71e64bd17fd4ab52d07a1eafcabb2c977648b50f982025d5312c36b4d3cad732edbd1edcfe24d1ab7c932fa66df3cab264a7c91638a23c68a558fe267bd398718f1905fd23655dc52929f4a89e8a13c8b6d8874fd2417b31196342cc0ba367510789df51e347530004d5d93c2badc70e8a9ee1a6fa76d26005e933a765417aef94e206d5a6d52f217bbe08cf2a8c769e3f63b253f13ac9e05377c57c67722996e71f6ac68713fc1e5f7053bae918756ec8382a7fa9d5df2d751eac7daa18371def29ca75e3338bafc421cc56edb1a4db8ad2f07a0920e87dd25e7d3557db013986465651bd555312bb5d0466554e33c579bc768eec3a2189a5d307fbfdcf80d7b091b818b0897eebeccd7f8650ad5fcb2a2ad26017eed97ae4e42d9f4a9c774a3c966bece6d77747db973b5a334cbb25ad356ff084080ee6d9594bb43e4265b201c1cf8ce9a1dc26561039f9ef0521d8fb0d92d6f5263ba8c1b96d64216a535cdc15e3410b441a31d04e1f178a501efabb88a537483e7f7da6159b479c543f22ffaafd5e522211248cdbb983839e30fb238864b263dc91e95fb29e698b7c9629e30c7ba3ca8ae24941e82c7f58e9fc46ce267c46fbaf74b03ef7699fe94f57dbc26d9de3a213ba449b2bf5bd2766ddc82bbe5e314f7b4cb9d8aa0c3ea1f83082325e39fcb2ec5111c8e98a1effb971b3d56dfe7ba68e7e041531df6f416d067c92d2d6400567fc8d16025734f4b7573e515e463d705d1fe1489961c089d89d990fdaf4210aa6959b8b662e22d9de0704091218e2c330f6d1ac8912640cd7d7a583079ff12853445ff4285031a8406382203575383f762e663d158f728bbc727f77c071d7bc557fe03612d434b5d32079c5ba105d022e5bc0a66fd07b193338e7f63767115f0c721d63c0584b40ec8b967093b452f0c6764236cd2c8b75736fec99ece8d1389c15a0fc71fe94799be5e0db9fa63434340e74c8c6109a4232e4a2b0450d4e88e8ef763aacca38028892521609bb9b4bd0a87c9da6edf9b501ba5bbc2e5508232f0a7c622c9dcd96a620f75f207b2d84e4bd947b0f0e9dadafd8911d6b29d11e522652e7d95099cef25f755e77c38d820c7706c0ee2e79d117fcac22c321b1ca3f995ad34ffbe2208e1dd777c46f9ca7aa2ce7ce406208ed6d541d241b351ff6beb843f985258d798805da5ea6dd8c57cb3ce1cac8b4ec75870e57887028a6afdfbf6ba2d63489bcf3289a7ac56d600aa821236f1bf44942be7817f6b3fb4cd5aee312760d37a30d5896abd655c02e1a9ee775d6d87539deb067d9f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4e724481f3d68ee8b899bb0d0797ef412d9822d45f6b90e488d1d03f999f943f423d02554be1341a36983dd8d86c92392973e07fcd09cd1fdf72b55d096fc3d5e95cab818e00e7d074cda57213e0aa071793345573c42b8d59df49ab1c5f6881e372948d9830103a09a7ce2de49baf05aed6463bf7c5f32ceabbc7836785831ef53abe71e1b73d435916d44c8b95bd4ea02ed5260f7864d9ca278cf020555a82f1905a6e3ab64d4c7664a5d88e907a5b7bce471ee8eacba2a89ae7218668adaf34a24c26300cb83dedb4b0c400df386146592bbeb3e8f89070dbf61effebcdb6bc3074fe489c07e3da7088d45d55e1e99eefac8ebd90e4250b112b6ecefad3d05305349f328c357815729d98df5ba49f9ff543af41d198d50a15cfdbaed458ea6359a50eb57d59181d69d7b7d874483c963ae05fe35865fca80e3ca3252304aea2c0b131ae85f9ecc95517ecce075fbf0d88ba138969a009e12edc2854819f17a41e5c46e3558ac43770a92103a0feb04e0302039c0b542ce7844225d6ab7d0054561af456c29f648ff7fc9657edb6cd7ad52e3e43fe1f15f7867801922a8dccff15eecaac77abf1fb3278a71ebc46d94a59485dd1f55a94bfb5058f392f8430e8e24f03fb4b8943e45b9aab96ee6e44c5d5c3dc9aa174f5435629eb3c31db9cf5c712eb0428f4751952718bb7894085ce2aa79ceefce7df8c774868bd400d045a88229dacf43d55095594e7307b80642f54f8d83c939a39ea8e9cde66c2f1c143c98f2ffaf00a5a7f70869ca6c60e8f867216e4a10d26faeab8a64b16d275a6912cb75646efce51c7551c28ecb192600dfa0a4dba91d5b21d1d6fbc294e98b69e880bffc6816ed8e12d7a43107581b8a61ecff70466ddbb2f8cfbc304d47155090d5eead63fb82f01b4d948712348c3723aad4b0d3548a205c8de5ea5bc739f9f64e31d24f707ba16dad82e2a721be5b57db1bff354adb80a025eec87d19c7b5db5d190402fa4523c75a5a58657f51398f5e39999d6258914e1099f592629dcd3612f60cb3ac2874bb46625ad7bf3d2295485bb174bbf394538f809b20020887601d5454b8e135de48b1aa983e5f564f19e1e48b857217160416c4919e391f0cc0059e8e1dfed825db004214be2388b0bed93b815eeb901d1069b54f9e5f725a74ec2022f35343730403427719c62e5157841a072a9ab0a23e5188e3fc432c0f34b4253da8d32a34b8e0ba3d6af5d9b3e9ec29692c522476ba5106663ba571d7f95151547c39dc77a0061b044093231e43e32affab7cdeb45aa6137a5f7f06d8462d0292b59a283ca42a771158682e734576343d7ac3724a5bcfb328aee8bd5f97bb6bceea60bf6adae6b1159725477e3de973167e85e1115404ec5665c419a0409b55ef11f5183e77a28fa5c82ae407df8d4915674cd5bacd9857e8719847b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1fb08cd7251952690e222d3b43eeb25a963a7512d3b8526ec97a265e1d1d0a5cd9381675548817f77b3b860b093c81b38b8bab1e893a0d7f5239dde5e5fb367bb8348c51272db55e1047bc69a9650c6229fdb1510302a1edaf5b237b0d918b69bb93e002dc049ec82992687dac4dd35e8f5b7511f1a8c185cc75b71658c9b23e308b6dc48105cf8ee000808183f5bf62f6a646532646071fbab5e3ce27382d587ed62297625687357416d36bb73c141f67565bd522b04ce9ecebdc1af858e38bd657ab18c142857788060b5e5ea0817386d937d1efd0fec743c4b96bc7b6beb3beaa6a53f6baec41d4e7efabe5df4db5632aa4b521c1f78ea6abf1b35860ec1c30d3c3564e508d17c42aad280d361e72b716e42e900a14edfbc27843db2f925869edfef6406ef45f3f6f320f417460ec4c1edbd9609380f97e693c47dea7dcbda7c67cdb5fc5e69c0c29abde75d821a0c736c349caedec3f2bbc1ae7e6d834992d13f59c69d7424747a9cfae2b254d0c2a0df632b52d97235b6684c3fed19daeb3816c30a28b7a4fdf825cb32f247ac14c7fb8d8ea2061fdeb027320d06b8298b383d56d75339208dcf779be6b6d5ce81adfd79a6521a376404b742a913a3bf01eeea4c883b757804db8d5b4e844900f8a14feadcb99d92f765626daf41ade9093a0ecb0a02777cb199cc13cec6867a57161fe30b9cacbf36db6d1621e68eda4b6916f0d574712e7960d6efd59f05589b550da444f37a0925a4e8f553aac4a1f9f6421712efeb7b497c413e1d70a4694bf288ebb8c27c5e49b8c8f186e342e056307933a9eff673c20c109191982e732ad70815cec6762b6a253b7de2e03a207822eeed3ed98dfdc37111ff43d4c965a070cfdfb475bf14685275cdf5e8029d75f4d7d2bc7a72e2af7924b22beeb5f82ba150f8c03e40da784b0efee0f9b34133f01b9c59d946f848c4fa61cd403dcc00d067292a5fc4359b60542339ce93c072fb730c3b502f3d9ea3e19d33fe1b58baf0e76a49499a3aef8512fd3042ce9f1282c722f9133897c657f2344aa357992e9e3ba207f059c1ee428f95b3457ac653196e0302347bd3960d0021517f652343e820c46eaa99cb2b308cca1a86f3fe85b558e25aaad494aa15e12635db45c2c01e24347acca10a5352646a97afebcf7bf2bc5bc8a21193e987a36f1acf1d4b6b6f934f7287dc593d05234db5137452efd513b8d135e50dafe08ad2ca7a266722a639857072c95d0cb172586b6040f0e5ccc1ea224b99e475890956fc2033c8efb6db7df2634917b5b9f0185885301db5c98dd9a4b5c473ba94ec4c7641ac3548ba5a6130b8ce3a639085ed47b3fec4b3ad30b12143b5aec5ac16467e8878618c6679850213158b726f640cba030b78de6ee8bd46cf3e0a8bd0dff0d79ebedc0ba030b8b59d1a39e6a0c638adc92ce43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h81a540735a51afee023793f9a5bb5e6b142698233cee735e67ee8318d49b4cd657c68472f76b7805f9f306aa9b802d0acbb2888fcfd85d7eafca69dc189f0994a300fb941ca04bbb8f53c29e8241d27d94a956d9b16bba84f7b5f85b5f1d36da5fb2ec66091e4c6d6f05baecd3253a56633c1f90383902225ca19762d6e4e2da53454e4b125dc3a0231bc176a759765ac24df76e2c9c43e588cb8a1abb509bc62d008d76438ab243a313ef6b530c4c973ab14d88175ea74dc443a9afc5666a2009e3ce5e00635b651a7bbb8230230792f9bb7f181f412e39d7d776224dfd0829b756659e478d28ad7b45a81c0e42f1788fcd01a8e63fb8ab0dec486633e6f1abb328f2f13332749038f9bc93ff7888da77f7816d25e8b0a749c30d28fd91f01097c8cc9d3d7e67d7566085c01e141f115113a4ffe4e3e38c80da435618fd1946b2d676cd950d7bb5bcf5792639c18983033778d2b9716af3cc3f9b42772ac72f69b1f8d3a2c508a3b8ee1a1f1fd917b5d8081bc1f8ff5882d1eaccf7d5befe84d2de35ebc7c7f9019236faeb2628ddf22f80598d2258c5de37add1f55f3f69eec0ca43b9e13c81fed5e85561a037261919675d4be6c3e29435c4df4ba65957c9381a37e1a44e88f34eb4dbcab0c089ab6294293bca21b1cd79140969d0bc647c44d4423f05516e2af1c79fd5e214580ab45e5f25639daa2c61724e13ff0a2ae4ac3a1e72b548a6c2c992c0686656a1e7ba7649dc65ba52e3276fa8db748190a2c77838d9a8beb918102a938c39b88ec6f8a26907dafa6e73fa11e4f4abe1cbcad2f40658ad06e42411f733aa479975956f1491ec0c4da05a860681c74bd6076aeab2266fe2e1c036374cc09b53eb822b0ebe2743bfcfcffc661e966cc13a173dcbc28598346459a6af4848372154f0bedf724bc10f92a08a94eb9f37323fccd8378f5e59bd1e3625a3a06751ce0a1037c37bf2f313caaa90468be7381fee28b6fac9aa08d26fca96b6723e10e0f6132b8112dc6e96f079fa95068e25d5a7c2d6a56c6561e6681024bacfb8329b7ced5f2a36150b00cedf45b494eed4f5a88b46d3e043b64adf816ca07a6febed3a54753c36f9330e50b433d77cc837797405f0a225be19e6dfcdcc39b0591cd3001285b6469a2f1c8b8ad1d0789e0253da8ae5c268eb1dbd81484ec34c639f4dbc7a4a7d590304260fe5d33d48deed7b1c449757f4be5180b9c8d303974b8fdc7d24c8e27440433ea3e14b43b5778a0ab796dfe6e3d35d16aa5c730020741956014199c8bd9546425f0c0144c8f0e07c4f6ec83324c5a0282d0b41946665a10d2fcba6b698afc79dd369348e970b6ffcb30c1b51cfcc39605f88837be3fd105da799c45a4adefe2f598db542cf0da98110e61557a4935c4bf05663acd93175220fd32cf01717ae1455fd4ff82fa1edf5c32cdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he9880c6959b33c4dabd918cec395efc07cff58ba72ccefcdfd65cac0954a63cefde32388276564d04a7eed2c5f98d35579baf6717fa4301c6cc35188618b1871de271a786efc5e576a0dec40ba91c2909d8d1e7ff3b8c578e86aeba82afc0c33dfa5a52ccb63a31c539c82078cbe85a20459bab3e8beba4ece4484dae77f3584651c9034d1b932965fbeaadb1224fe3cd4ce24dfa8a5f289c59e4d54b764c8473a21f1b4671f4973c3b15cfcb31f4f97344d20265ca5151493540d3a216df525aa64d042f9ca33a819fe95722f38cc0937041fb34f4fff24a6e15a775f626c18eee5b9d6c193d6b7aa7c6b278bdf8fe42c7f67961556e38a9ae37daf70d32e5ad3feed8d1a81592963e206c7d6aba0d0313d46a19ed4a4aad9981be3183317f4b51e7cca7bd4a0a322ab6f6ad8f6a49f9b0cf73cc8602cad75e4050e060bd7abfd4d23221dc1fecc617103466cd767bbcd3c7861783619a5427cff1df6838dcb62b5d96ad500387079d7ea3ae373b3449e318bc16e032befc2116a5c83731932b2320551e4e8d4b957e2459682c8bb781fc392957d8619c26d47de5f371a6d5585c5ef1b6540bc961febaea663b3e5878566da55f96fa274be4039a48360c71d6d28dbb98630bba96a195df32da6f0c9f15507e0195ab817640f4c3672c8e708c4be8f7fa3eb4b208f1b749fe30878147f4b5e6f338acfaaeeb7c18ad308d76047a679cb09bc960fd0e1ccd842b4e822ba4db3e8b164fbdc138775daf20d2c24b0ced8d8f78d6b3e5e743054d295b8925b5890973e4191cb559630e9899c0177a8088f575faa78243792f71e7814a1365add9518eb907da63aeccafd02e924bb1f153f36ebc890f8ae7b34a2149c6405b6208f51f3b1f262cd90e3507fe7123242f802fc7ea6678e5955d62ea8170760bfa99fe90aa3d6d60d5880f1d72a8b9de0d920faee91fdecf9923b67d291b506d2be58db5ed9282328c57407887ea42843bd9153a6ad570fb6c45ed008773c40aaa86423c0ff3068ab1c179a7b85e3a7bbad28c3817a22bb8fbc8dbcccfa443cd9712bd90ce0490dd076b17b34c53a34a49b74068640159bb97b0abf0745c8c7a923d67caa5f2880948680725366850c1213f9bbebcc71009235d20a9e7caeef48d48a48d2d3e8baafb7803f8a837790238aa567804452267ac0ef8d0988007380a1de2a34ca950fe7bd4c28c21cd0c76652709343dffdf22dca860302e0a6f9cb0cc479c4c3c200f30f69aea35ac3b137f6bcee89fe31e687616b41a6a229bd98a3da6b7b47dc2614bbe3fce071291a3236d6b8e4699fc2f1a7ca53146231a36332fae240602233f558057c5e6134e6c6529db6d7656eb9df22bfda9fe9826ff886bf2015045bc3d2d98675d7e2635e7e2f596a6f3f647a5fdc151751485b9f1497344721f51f94bae20fa441028cf7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1300daa07522e42af7573e9ad427e94aa217f52253fa0565c7ffc2168161b797f2306542be7d488f2bc4eddf8f5cc4da3edf92bd71e1a8f7a5e718123a2fb1dbca99ecfcf9abe25272ccd3e665d036aada86109674074479a0e6ac23beb82a7814739a9ff3a044a3d3dd79c2a602b92b9481f2ffab535c543e13ac1c22f469546fbd454ccfd0ed40c34130f82887ad02f277fdbc884ad1430d919129ae82664bd64b15b73c7c63ea755c66078eae97dc5999bffa32673aecdd9ec5dd8380edebfe20d2a38f0ea3f8d8d13ab3423982e0dd7452dcc3c900274f46853e93d01a0f5b156e34c9c754ef9cd2f741d2846ba7053fff01cdf7be241dcebc63a0f61c77b2944dfc31185b1255012bd5a6652627010a67533de923998acbe91c04b39a0c0c66225c3579e5214aab4c7b272a97bbafaa804984e4f6c49daea725ab2d993f817cbb0bfe05ce0473b1bac0db206172da7b8d070c4d7eddabcdde10bfa62a0a17e6ff113d806c45403d55806f532c4446193aaa7c0e70101309e57a7d0d9c64a60b8d5df3c1ffdbe6b2473e0de6431e5e35b20775bb16fa2048b90d59d842e38f24babd7ffe742edc1c56a8c8b89d0ef6f511072e6e69ddc45fedaef6fbd391c24cc28748e13ce859eeed008cacbf629bfb5186c748d395b03ccc673bab7b8b85cff0e651192822040b5fd8948398f8271a9f0623ffd5090ec2c3120fe77c7b095b0bf45248871c423db4f9a2729e63fa673f2115bacb8db546b0ecad5354209798f8e83e1bcd80c9586d95998abed56a090c22ec8eec77850efc7e32df0b6287a20a4f3598ff6f21d4791706f3e986231da3fbddf51067fd9c2f1b88b618d9c4df11881fece40fb938239ad56d3a48af87e656fbbac5e5f58b6fcf03558ec72f962c3c1ecbd6347ca53f4938fb780e67c5cb801aaacefa5d199ab3988936d3059dc3904ccd27d22146ae79da838512d74e2f090d50934f6643dcf3358da109ce10e5cf0432c7d831138c236d2524260ffd642a8580bb9aae698b0ec2af276c6d55e49d6d78aa88e1837181711f37873ef65b9c0b2195ff4030998ee21b8a25515e89c4bbbfa9c5f3cefb557a90156d0756a76d7c1afd2f2f7bf39ad35e9e57f79e57d49312e75efde6603c1689226031828c02dcbcb464e1fda18b3ae391a371b4062cc0146dbf8e8e5f329b1cb026702196b7ea441c544ccfaeedbb98fc8baee67da99a4e0bec781e9ec13bd50fe901d775fa78172d096dd6701d3ef5c1fbfecdd6d957871c68e14887987b431fcb2dfa15f81963b5a5cf5113ab5559f309700c60767257317d7364c3d7d657ece55c0b764adf4ece82bed8ddc56b3cf280ac0f239b18b4a71e8433ba5ac3f64acaab4458281c625370fd87e37462c5ab59270572e903f7517268e8487e50e9aa2a1733e6da2c3eef2cac15d00b17fa0afc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc15cfd43d72fc637e0855868e2039264b45f5897ab1c88728f7706f7ee5e47e4cca909b5b9fda543bd141514a96cd3253783a676339ebee700935e9535973c02be02d7c49ad8a0e2c13d0b4a18859d59334a07d4113a75bfe9c48b3396deaf3f2e5588b77f8c8835cb07ce73ac5ab37e93dd7c52388b2626ab45e062e947674320d3a0a8554616f75d88220fdb9b300039a5f451c35026a7466c3ede04063d9d01b11c064857b8a9cad054be487be0da12389f5d97c0958cb5a5f96478911c7cd4ce4f0caf02b31ddebeb29c545c86cc149eb4e1fc705a5ebbf0c177565d2a62d3829cfbbe663c070032d203259369b4a5ec4bb9b62a29d5a794641e620c8eeb9809c2e04495686caff2858e5a914e3a5247fd25e12a2ebe35957f1deb9048e03d2d51fc0db3175952dfaa7a62a23fcb696e917b145bb5fb456afd280bde4a6351e5977926eeb86a6cbb5b769017f7271bd4fd91d6bd6a3ff28406c631473efca1d9195f3b9dfd6acdc9c3c7e173f7649ae8d5052068a376c0a9dca0e093752ddf0c7c154368ffafc7f44be6662828f17e1c02d8e2eb49431a709b172affc8f066231d15109ec760d7678f27ec506fb7ca7dcfca5dd4fc667449dc416ff169a6ee857c64c9f05cc480377a84ef4ef6649e36efba92179e64165d95646c354ca1aa3d4dd588e491c0bd9f2ba10ebcce1c27824bbcaa1bf7e23b066f6b1af548ce45494d7a3230a75d27599344d14f1ae129903230c1a5bfbcab4d05878c8ca604a4a205d60afd9e02b90f4d722ce677a1dda9f3106fa28592b2a1315d93d5c1fb65caf44979a436a00b3e29e850c496c37fb6fb8ac17820ca6ca337004ab4b14f09ae02c61436db32d8185b17c42a43fed699359c9d869f50023b7cd004903b4f9ae5cb8afc12f5f2ffb02756c1b680b8b768e99c17c4c15d20a28de7a5e3b4e3d6b317028a52e2a9e511c677c36ac5c3e000649028425d13d3ea6f454c195d8e3f0d7afb307050c39256b8fe5a7c44287c2940262147e8080abbc048b8e49c75fea3a4241b037bb45f1c56d6d3289f846c96a04cca9be310db91c956c7696f715f2af01d607c45f303c77b77065e13ddd06db1a3ab0deb9a30a225e274498e9db2c75669b87a2ed97f18be3564c8691a78bc17841f749618eaa1f1c8b30f4a87d60bb8342f4bcd8112b3f0ed220b4597629e4a2651e3781e0d9c86b5a9227f451867a11179c36f7e7bdb08a4ab9c226a64eb81b6ca219d584a8abcb7e72768865ca2bb15775e08fce9ae1311eb250237e09629c5298461b632870f06e98e39c29c9251a540134b4afca071aea96c5027f5dbde7ee8de17df6689981fe693c0493b7d27323a4cface44158e4b69a5a41f8f71ed5986bb10a30345a2b13b3f2d8ef749839845af33df8f594582d3c51d2bc2a8a4e27e390186ed7a59781a29beac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2fdcf4605c687c10834850718105bf66e514027378d49c27a122d884424a0602e7fae49bdb7d67ffa5f00b4fd0a1fb8a5d1dccea5a8902f833f31620aff6be4c230dcf511ec8905249c2d81dfc949a955d293476504ac71cb8517db9f508c68629c2e8e5bb507358456192f5b47ed6518e72b8e0ef53b2b0a71dd9aa883b60764f1ccad603eb7668f780733eb83f530afe8ec3d8c2b8a672771ee34eeb9ae0072385945b3f9bfb86581c8fef3e077895f7cfe8c07e5b0f5ba19c9bc7c2c34a4ca45ca8feb1904d5fcb2ed0c3ee2b2d45f4ac2515b23d134e563b0c382e94bdcbeda6953e5fe0aa3601fe15ea23a968d7f1d1890fbc075799dbcd18a79c11de3423264ceaa65b23f15d9bb9690424a3572d2fc3e176543f36e03ef78c5830feaf4b230fcbac921a2edc96a8d898e8ae65471b3dda164b3eb47b4bafa31d4ee5d8e6539e8d161b1e3b5d969470ba18dcfc6cf6c1b0249af3d858c14f99944931ac494f5d8f2807b5d3feb77350012f5526129bee71ea15c0c7e71a6fe84b843ca6bfb22aef22bd1ab4204d3eda9a8b86a75bd5287f3f8809fb463225938f5fea56eddf9c5c340182bbdfae00362c2ac0f399a1a8350c89e7c329c5e1803032b07c74dab2ee821b90dcdae65e9afe4a1a39045c7464be970594f8f149b7f955264b18d69c58d7464fb85a7d5ab7fbdb0ed1b09669dfb04ab5ef7b0412deea4932283ac4f25bbbe9f37cc151d440a5cc03c8bdd351665fa899f88c25e1422669ee9a96a76dd608469dd21a48a33dd7b344f24c815b2350b1d095f7e1cfa2c84d8dffa4d8f6ef68eca5cdac5095fb6744ce618eb8292cf91605b332efc99689f31ade487701e12ccdc86e206f6ce2643583b9af676afa892a975237c283cd1aaad81baf66d2e88e97a2927e8fa09a4995f295adc26d001ba5715a32739577dfadd94560789830180f0f56b15c66fe782860388a6971d7195bd9850dbdc3a3e44a1be1d9ea823cf5e1705d433974b1964ef437c8ebc5bd4e7f86e8da63d5319d7d7fd96aca2c85aafe49cb6d4c967af53a64fc7912c0a9981598507b09abeed92c568b62c2018add9a39bc8c44c8513e562757b347b1b5b98cf64b42b9e6ba32c7cb1a8ed47b2b936fca3a9c74adb1c630d804496c695fc312628bb343affebc2e16fdfe90dad26cb4cf97e3569be0176ee2d8ae017a3a75736d9ae058fe49c10a99578d13639173561ff3afcc567e646e3474852a5063268583f857028830a23888e5685d209b2bacf02513fdb01b0f97681f3bfc2e1c0dd9787b19c8280d7ba152bda37a1ae0d082ec22ffd4c022b3fa7b458405d747f0a3cec2bc4a0efd0c9ca3ab53dff64c5271ad7889ccec97a7a3ec9e66e6076e76fb89728dffe521d4c860cffe30eeee491fd1bf9e86c6a27eafc9cdaad245fc72c769c402306b01cbeb683a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf43cd66b08d7872a0a4774107ec9607d403199461847d05b2a9f4b647eff1335a215d140aed6582d06479b005050ae7380c5f3b3ad2aa82c832efb7a540bfa71c23235536ac8a4b6ec738dc0b3146bc1851ad6da41378a1e38271b5c4f24d940aff4097dd4efe6fd47bbc06d3b4367a19b8c2326c43630d9cbf10aab2067232bdd7f76664bc78e3623ff694dfca301bfde2e411e7c39a6d7a74fbab78ec1dd297f738d8481bf4cfe7f97ea0ec156721fd05b9a7b9174c3a5520b17bf77b68e7c52f0554ae1f4d721bbe2ed89740ad5e84442cf36ba12c70f4ffcfca01792d055713fb8bcfb6807e4102d926e915f1e794e7fa71d014708a661c01195a5790c559cf7f45369f1b00b70f04bea8e537644bc1a6286c099518a5c7b35209ec45bd062e516b4d276a311baccef3245de23aca2447df612d58240dfc864f13520a14f7d67cf2ec30ff4e206e2fbed7f5c1a23c41ea669c9ae9469727949ecc7b398a0b9c94afdf0e0599d9454284ae8525bb0d150bbb86534c054cbd364be691dce647a3d305a8b4bce0060efa66232fd8eee0a6346f122baa33db416d0771b4747503eff50b7e47115047653ee5a883f2f332a74c364d5c59e9d43846e688dfc7ad9a505acb6c434605fb581b283b8a07a8e4171dcbdf7f7392f95f1fa28f4ac327b6cf99af5aa5d54503d8895fe64855ec8e30fbc4d0ab386726a0fb6aa22d7e781e780d9c0c1b33626d7ae4aa6ca9eff2f8fdb952eb008672a267644023254143f41dcca3bbdddd313e812cba66bb6e958a44a1ef8eca2d39edd8cc5c5ce2bc3f7ff1e4f5f211e05e2642acf4f32ebeadc80fa8de2781fd3a1bb09e74d16d281084c0feed7e109cf66036ff2f1bb0070aa3e3eebb931f7e29e207670db438faa3037271330d1a77cec61dc52892da30437e0b732bb63d894c303d5bc70f1d0a1871ff17b91cd12bcac839f0d17966b1a52829421054f14bf03b6d3eb53b46195c55f8e13d63ee8f0cab9688a5a5505aa0839843f3fe9c18ae985a64fe6e431fee8738cc8effa3578d0d4be8ec5b245c7f6f351d3520f5b5bf7f2baffefbf30447cf5cfa28764125b3baf49b889def946f94e1a229c9018e87f69e0f06dd37f730048906a9a54cbd4a5ac94b76a7c30cb15c1fe1f8d26e2035430f456942db80f91493abeaa475517cfcfd048bfe671c15364960a70c712321fb9d9582d80e6318a84a7b41d52909d62c7e4b3ad148797bf9edc25b003e06b92a30575c6543447571beec7321aaff9985d296adf76601ccc282b26adef6fda2bdea5bec306d84451c5692e8846c5df2ed99d7c94b5c86def93497906afa238f6bb17359d147306a385060c3364127366da3b52c9f29828c7d41da8cce1b6f32545abc5d2973a8858913d9c5f65af15a31c1b76063bd9bab67002cb6ac0208742edd7cbfbf16526bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7f5d003a6480c4d6b3a23e29f08531f807e454ed9d07a12d053dba799e5de9613f4935516a7a1d96d3a41172fea378d2f8f90b601571f254e4d27917aceab6c918d015bf3d5861b78f2ddca8cc4ab63a26dafdb6f31e52ce406bc089e7d72068dfe5f858a27843c058b9206b61dde9583dbf9701acb6273d275c553a839b816c4064609524f2f5985ce369c01cc3e80451258188a4553b6eb4c84728d78b46be84b201a2abf0edff1867cf7fca2f15f88c132591da4a564d21d80a4b3586c5062185c37b229905afdf10020b9bbe75d5f33cc502a007368f25a5e46f487dcbdfcbea8082389d91fef4b4f6904e389fcc06dfd8f0cb22694857a39fadc040b49d2ae578f3e537f5c779d28b20d6075e64008412f46b4efede775b5ca433f8ddbc9178da2321b9b30db1ced2352f272752f0e370d1a4fbab54d3d2ade369f0d24c6adb10fcd05b8a909dd29d945a025d5d8cb2879ef37363619b927f83255aa41085406f12170f64b95ab2e06801a34c6153848b2838552879aa2b67549394704e3fd90fe01aaa788adc153112eb370a2817aa919f91650a2d83b444bb36ea19ac78033cd34b420cbd979ff506abf48d2ec0cbb2e8016338a98b27a38a749e6c4cfd600aeb45680b71768bb9b34770128465a6f844f4fb2111d6134bdc85469a97cd18f384fa77dfb422aec6154616e20f1cdee36150c0ef5cd0288cea9bd2fb6dfd0bca440efc2982096cc9108c583b373da8661108a8e44e8db6768dbf079695a4e1eb71478a1ae23146a5f5db0fb6e25a04e72603bc8b88f1f0ef5027028444c1544fad32cf5fda91ca4558713d3baae08c562d057a491588c7c72c0ddb8970e70f99c898ddfdc62643635d1891c18671cf9a087ca6225d5a3be72e8426d2114e1ef593c83bbd9b104d44747f519e78f23da58f0a3e2d8ec78882e0a7d3da74f5dd108977247232800be50b7f5a6063e7ecc793cfcc44e3307cb981d3632d5d0bcfbd40721cf29a5f30dd6e0cd06619e89fc4ee9919d9645c5b0d3b4271d1d0cdaff090ed30b9c745b930b1a94f29b35d732253860e49cd62c742518a0bad06aabfdd1527c046403038c0dbe15175ba589898786c5b0216b326ecf236dd6557ceaafb21c873f9b50935832945a7878387e43f1a1d7884234fb61e3615f52ff71736e56f789478aedcba73073a5f246128a165d4f6d89c09935f997d149a1ce45dde2b5419b946c1679160086f03ad8e1fe2236578de85323a5c318530c8baf0d2e0effcfbf4eb3dcc54e0fc483b745cf4e70a82f9a0bcb3db4aa43018a22f158412e510e39b554a61f728bb8b4eaeb90dbdbecdfb6b9da05900145679a485949daab82c7ca8a4bd712bb737bcc31e1dc5e5a1ccf2f9794725baf4560fc36455ed4a1bbd82aef6fc27aeff1a0d64742582b428fc7e7ed846cc08be0b656a6606;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hff919ade1d2334e0e488aee88e19a14cc61f56cc46f4adc09e2adb7fb4ed34e00ec2f29615b0b04ce598800ebd1b95e5c47c36a4109b9ed61320d52438cd4b4c2f06dd25757c7b0de8c7c23fa5404883150874f87117f40fd83f692693046ff2b7fe19afca5c19d54270cf86dcc5bc84324844dac77d79f49360853f52696f881642ab9a108f9255551ceacf81f4164071d255eb7a52861ee98536bd713f1c2814d9fd8e3c258bf3ddac4b7f88f47e1bb2e7ba0784176daf779e3e27bd4687303fc184a5cd515189c7f065b1713e518fbf326ac4439eec0c0e939c399c11531c0df4a15c8d86d27e2498c7f2cc6731dee04cff43cb64bf09eacfad15d163ed07139af3e7598c9e3436b0e82c22d7657306047638a9ac5d06470ef8c93a528dbdf98ad2b70a953e8b5eaebccd11f7fc405a961f7e539ac77c5ef45f6adf8d866ec59b30188730c6b09f4ef190cf37c2d0216d88c543f24ab2d747fee107ac2fc713a389afb95e09a869f1b85c0bc6392b8b5fd24282381df7345cb425447adbdb5b9beb4246665dcefcb9dac12a2dd2f80689e75b1a70862d77ef0c6b43f996d6af859708371620fba73e58dfaac37e85f6fffab71e8230f7030c2e357129744ca2a746d3c102775c4565c2e7f2bf99d58d30fd810094ca5be10b4f1abe83b4768a9c282ed0b704b3143d40531cc369385d34fc29b9ae93ba42f6aaf251c885556c6b7a0f65541970cdf67b535ab997ceb101d48c927f58e8c2c2ccffdc81bd24507ac8ed834596eef3b13990c28f1d7750a474aee5d4695765df66f86319654425be2af9ea4d07b8a991e66336da0aa4e6a1be0b33d8107fad1485ce75681254d443bac2fa5ae3f062610cef16d28d541daec760f415bd50baa612a7093099cb3a4e4c99b2242c9ba236b5271543684d9342261f5740f286574d39f4ab19434462d97a95776a6412551dce431fa33cc22f32e9a034b418cac259e76ff47773c5672d2b43920ca3c52eb41901ed8faa3140fc39fe26f35c19c91c4e1585fcb54c46e1457fae1cb1c02756ca5527d0cf8cc2b1c96976d889ef91056060dadf5dce524c6fcbc7efbfab8632811b40613291d69ddbdeb416fc2b8080102681e3137623d1ab6ef016a2fc9be20fb62699582e1f2f7cec92986c3cb677b515257873d4b1d71c164094ecb33354afae30fd0158c44e4e405d61eba689babffe16b559ce3c1e68189eb528d2961c595e33f1b78b783937e1c5a99428ba5e2ce47d5c8803c853adb29ba96077d334f3d27fb0712fc270255c786569e0b6eb781258e8a26985dbb2252e90cecf6c1b26952495dab7f6bc56baed2bbf1b9cd461b1761c22de609eb7b179e33c423c070e11afa99dcd84f1cbf57a6e10f9c4883324d9f383bbad20c8d0b9075c4f8988f18fba5a805ac0b9e0b8d8fe12f11a0055a3e6fbf2a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6946f30e4df7de385c10a4ab0f8bfba27607c150e9624480efe3948fd658261403fb9a8cf766fde01c3139228b54e8ca3cc3df51abec177451518623700193d475dc6bf1f0f4e84e5c4691aad25f544f38c8cb36857a84ac623eb0407c02a3daf0ec1aacb113b1eb47227a2af9a61db0a2d302e39dc1890a2d39936d5d7815e5cd2d98f2a94f5d46a40d698a6fe73131a9cd0772eb4f8e54077d3a4bc43267e293705c1817dd289a957ae666d37b8ba267507980fb57df8c3b99861a136f9d748e8c4d5e5c4a3358efa777df0fa59da9f73a3524126bd65aeb4fa755edf749f6a9fd82a51769976e5f21c640647b6f0337131257db531a4b5058c8866443e852e7716c95f3973597bfc8abef937b2f4d49a44cfb9ded6acd39b0ad02b767934ed0cd2a7f0edd2e8e4071e24d0c14f292104666542ef766f3c2de42125c398e94e9bb9ecda2682563cdacd0a1449aafd992ca25be7785cf9abda88775573a6337a73f2b9b7f8784b2d597ab0c107438017c6c25293ed04f59d706e47c161c9a618331f9b20475ebbfbf1b38f31760ff2df734e742ff1863f298c5b7567ee2e968b4184e364d1d8866ed214ef2d930064ed759d496c86e4660f1f3f7a53dfb2a452d052489a8578001f951d52b45b97782d1bde5bfa709e313636a3234575e307c4a6de51628b34007ef99b2ad52844ed26d327da873707ffac7d692e4faeac4bc0877bf86c4e8edc23bcb2dfc47d95a2d486bcec819db28a0cc7d7e202c7636701fe15d1d3e3fbc6f7538f59dd359df7fa3218d9ca76226e63c9fd2aa4e4664e578512f4f72819f1e5912a22781dece8dc84d4cb0a3ea1adab82d90a0459550e44b2c71308ae4f3e923a275c8fd3f9836d5bb5dd1e564630ae7d75a4e69aae5e02d1b9c741cfb811b63344e8be9e591866a9806c9a02e84f17dc8d914e56d783c332574e220cb8bc8df05274ccc64c6a7459c991c22a87c2487b33c8ff11ce088599bd7a338c08e150e002ef324ca444e414a8be461aa1ba70af5cffb036af0041ac9a0781866bb82b6548c680635b433408b2baecdab8ad2e8fbcfa86307e88c360440dc5f81c93a93970504b70efcdab0f19c04fb2a8b1c7fb971ed9db9ca71100037d1959691f86ed10e4aa77a2c18cfa32d138fc53005a1c2c82e7d87565b07cf910e302ac6332d6440d4453728edbd882c9d603828f9758d5570027efa425ebeb0fb3120f57244dbd2a2c8433c2cace8f7a33212212ed29e09802b06ac5186c96dbdbc63f8bcaf6a0776aa5143f39b0b8eaf2a082c1161c06360bc760350e40c64dacdc01ce220bdd73211c2ec9cb66e93c7c6d6f6b11d0748f62f504361b974590da60577fa01043d77bd8f7d538ffa93fda1398479102bdfd1de3e1f9c103161d2cd976ab35090e083a489658724ff1329069936a7e2f6ca001c03bd9e;
        #1
        $finish();
    end
endmodule
