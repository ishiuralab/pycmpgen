module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b655646e5c675a11d74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b04fa66f911acadcf1a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147ed92e164576db6285e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fd803589fc0e3f28bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145d86a836cded110e3c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b0441ca13e6c6807d3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135a2e88f37178806e69e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2790709304d5ad4225de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a487252d56bbc6f45ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34590c19a9765ddc0ee8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha77b6633b0e2baab0a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f73e4bb6f4614f307d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ffdb57aca5eb4482564;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habb68e1295ab66052455;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9f304d71328dce76f82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64352a6e5b2100d234f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c62e7b188d04b76e077;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4d467d14f8661f09e53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e436426bad227f85da2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142851a92da788789878c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f68efac26e8c9d03b9a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c14b3eefe6303f23128c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8664035547eac01882c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b6f4b8f1cd75dbfc103;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea1174171881a010478;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a35816cfcaf1c226a237;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d083d80cee0defe8b953;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c7eb60cc239e99481db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db48578ad648cb5e2591;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1719adda9fe103cb4be12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139c9f142736770bbeb63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1554ab04654c1855458e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc8ece767c57d8713cd4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b578248b49d96cffe46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2bacd5833a294bafc13e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1843eb52eede400f6bc41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1a9627ebb1742949c44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf72c8d61059012bab23b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43f21ca71f9a6b00bf3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144b4578693b2c4ff6d4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h273f28ca600b7a3b5504;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bda0b0dc090a6f27010a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffd3096eb0b13c6d2060;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4860bb3c87615f7a6c46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28d63bd3d39e572e9c44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ad8388bb5e39d41cf73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h637b8b1e0ac712010755;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8788dc63ef3db8b87603;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h708b35d9b05642aa503d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h216406ff92d06d135ed0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ac31377ddf3e194f1a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bddb2896f12fafefa9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ba470ef867e94dc481f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1094d43945a8fc21731e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15328d3f3a2cfd6b474f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d99960f474d47415965;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170a5fa0e603c1494e702;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34653e124f586d52d058;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d21137a4626a9f93beec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd8d80278a32b12a4a02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e24ecd0639533cc8a2b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a30014e94ba1df2f8edb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ba7e4abe02920a80578;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f9477862f2dc5d26a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37ce50b2ad9a3c43ca21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc206deb487bda470202e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4ceb12d686e166c424c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha66c06b5e6997f13e219;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h220c9ccb48aca1bd2c47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d8f75961ff8e137cc67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a466d2c584297934baf6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b91590a30ef5a270e04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a384baed5cef07e53ef5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16152e6a90d5757036f79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b695a6dc3d3c4ef868;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c3f99d3cad8e2bf2958c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1192776c90d2300686b65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e447c911bf12c7dfbc27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3cbf1b1131625132c9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62fbe464c095ae97f6c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d18252d1c24cefa379d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170a5b502cb4502d03363;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f89e6d160b45c0b2d2d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185345e2a581f7d8386f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6012af9d1d603c175954;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h616300866ed5083cba04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1699f5685085adb312d3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf2150ab4d7f781e09f59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7118dbb830252889591;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111ddf631779550a84d9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7b9823d09b51ddb838d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145e4c4d22a00710940f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddb1773bd07ae9e2c4fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b1460d6e90864fe4e62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbf12c4a427bd3c664b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10df76ec1093e8b51d81d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83b8edfe266512241e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ea95d6be00f1cdc1c47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a88d669c268f101b3583;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a692d670eba0989380a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1183558a9d0e8fee39576;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h845f7e45edd578caa8ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd0f17fc0c7feee0fb71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf3a524257ff09baad98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73c91358844e5d31b371;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1408eb886ae83447d6724;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ebfbf783392eed5a000;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b38d58a5c14e207859f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac353c954e028cc169be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h569c1123d82ebedced3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfd886bc5f64b95dbea2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d94b726142f1f82028a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dada00d4a0a06e58247;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18313b91c58cbf4944c68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147c50be510cde528782c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d40856f44238fb5d604;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d96ee63e9f6b3470494;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2a53494ea2b7b1b55ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h814af2db18fd9a68e4dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1449247d50157d728398a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103a9c1569b4fe2f33305;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113fe25e8b1abe747bae5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e326332e5c3eaa21bef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192bb5b4741bc2e2589c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he99155b82c2c35ddee5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6e13e38c2ebef81f7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119c24f38636cf37519a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he554077cce2eebe2fa8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105ff5928434e214f08af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52965be1de99d0f622ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf57340ee7746c424b00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd5f47fa79c233c054e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6ea887ef5568b52607c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19fd820d157e7ed09a1ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1438bc6ee9c49a60b48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f74d5a60d81b214fa446;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc17507e2ad00988e40d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1222378f0fc0070d1694e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7d7ddc795842e2c0c31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea84531b44c2ba97f429;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ea727ab36e3b69c8611;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d358ce1eefc0b14fcbab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82fd8cd9bd77eb5ae38d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6cac51531e16477f418f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7d900f47441214a55eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164941d31a20291960e84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd78d0ac159e6b256d42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5773c3e7d5e530291eb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de1d6e1dfcd96951afba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2ecc25822c23dbb984c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e22ed0f8eeff7c072cf0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d2bfc0a80664292be06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd88af413f63fded1b76e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h136f41b3647b5a43ce4df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6469715fea39ce1ce82b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8de89940d98a80798e02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6725575acde19f6f2e89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h630e80aa68050308044f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6742ffab516a8ea6cc90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84f7c71974e4858f7058;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c9209ecd420f6f8ea42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f34c8d3831ffa284c8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h585eda9759376141513a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca98237bfbf619d9bb0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1508c2b0bd342ef7a8180;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76117d35780e504735c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8fadd06d7ecc9b89393;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf10a333c781ac8486f71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1283cbd8d49cf3c45f09e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3b559e40a5ffb908385;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161d3d74007fac7728f5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76543cff91a0e2452fff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbd7d8d9970a869f3ac8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fcd63e75f24aedeec6e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb91a1e7c0ab6bd50871;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cb741253ea541642f98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e6f25aba793b4c62da8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c67e211343cd19e537a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h362f376660d901449cd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h791b083ab2bc5df5e0a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18650c248701f9e09abb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1decc787a599c3d21ad1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138d9074a5c1c0804f5e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19416f8a7e381ff401da0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5078aa4684f133a89d8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1589a4109663650f42830;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18857c2b5800bc04b1232;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1838e0da85ff7ce9550c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9efd89fe5ebe747b1249;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b343c354f7a9a038790;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10154cf8dd3fdd6fb85a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f8c807f43db433b31dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff094f873cb0d3c9ffc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bc9da40bb806ad08f07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heafd1ca4ab904aa07428;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75364df4785065f20ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8accabb811a7d564e60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bc61be1463562b8e767;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cfc1953dea7037cd64ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h439a5348dc72168ba816;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb17b727b66e33d8eaf7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h770aa08bb2987aed87a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9947b78fcc29599d907b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7feab988425e48a13766;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e89ff25ac604325ccdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22bc2f8f260a7de11835;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd36fd4881c763f04f9c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hecafc5a15b5b98e726ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147d52004fbceef339501;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70fac2a4e1785b108ab3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe5db1c2d81486b48d8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe79481a9c4972dae96d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d379cc87ce6392829d44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58d55bbc4865a61c9858;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h205a2ff135af507713ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13338770b8210a50c3edb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d62e05c0149866afd82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ca2d2dd67751f3a3020;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1671c66c585f1793b1f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd18f7a22b5485700bdf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf68a9af692900ff6f895;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8d78047dae6360a7b59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2639ccccf95f0bf1f94c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a3bbbb6f68bb8b057eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1252c1ffb641c3c2d6d77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18205d9ec6144c9cd93cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47976cd35e37419468d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b187fd54288688ca50e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6d8cd3204eac5558067;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1995ef76c91999862bdda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa6826ad6882d6fe8f32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd914e4c1cb657091df4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143fbc40b432235b3870f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97113f6eff009158b89c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2a3bf1caa10b78c488b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1318a438b17f786acd1e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8169077eaff669faf079;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae00abe84fb2de8eda72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf194890fd33a9f432bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfcaef547b04416dbb79a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a370b99119fa36dd323;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc58a03cdd6c4d3a155d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152cf6c89896188cf2123;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d3bd0fc8f509b1edcf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2afe560ca1d73014ad7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43f913d9f8d026de269;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6175823f9c5bb5e4ad40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185337d7b0bbd3901d4f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6a77422528beff1f36d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8468b6a05e00bc0b579;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc67184239b4fc636155e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6cea85c93365678bc1d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8555930539903050302;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7954e07c88bab84de43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ce7bf4b38277ebd6cc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1943cd62cfcce70c3ebf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b78c88460ab2d021d58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ef26753697fbd665e61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbf3623238ce13760c0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb7c032131ae1346b53b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h216f71c69aa7f542c806;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dcd7163928a9379b785b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1d52863d9064b83302d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187661925a5164bd2c349;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h727aeb9d265737bcaee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8dbe864aefa24405afc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he01be85894035fec80dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fec7022f23009487913;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fec642f1cf678aaf1ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb108b8cdc8fcc7485e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc005e609da0118c93a84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdb646895bfc09127519;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd253851afb6fe041e2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38a60f6e624cdf61ed5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61541842566466cc3d51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40a7feb3cc149ada3d1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d83ad11400123650d42d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a83794ef608108e8b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf36d8ca9f1c9b89ebff2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b9a5a0381eb730b0e1db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52a81d1aca608116033e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b643f11c900c2b8a470;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1327834fcb23d25cbb43c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114f4461886f952290109;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121410d026b7c1a543fb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb16526bb27dbf194cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hebbb81d71fece8fbdf50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fcecea50fdf639b3fcfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1272b77db2025af00f6b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ce49ff3c542cff685aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h166717b66b5d1bf776498;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha45493ab31bfbc4b7df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189eeeeba8c0db8fcc9e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e7a382820fa8f52d7f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1ac479c4804b1afca5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3a7fff5a7e67c44dae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b8a972f176d235d49b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7b6c04eaf48e3e7c5bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196dd52538b4a1225d668;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd07c9252db99135ddfb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9821daa2c5e63e34d7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1602a1d3d288599be64ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcff9538a35d84b0bf204;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1856679f226fef5cecad4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13aa6eafe447323ca2773;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4cb3476d20368d0eff1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b79a8e69cf534fb537a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4ee539957e955fb8460;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168de225f2ac5b04c9193;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc318e3eaf873541f5ba5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4d858ce20ef52bbe182;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e3c649788a7dadffb39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1212b39864dee34fe528e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9d82af3d63c48ef0ae5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dece5571213f6e94d2aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a8c21decef0292540be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4778105adeefd156c77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36920354587c0fc8983e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfb3e7e259348fe91dcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc77dcbac6e08ac7bc568;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1951f93176541aa842637;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59215acad218c32f5553;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f82cfa9b42ead4dc01a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fe8f5ea1a4872bdd469;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31d4ed27c63b5a3b7d91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188c60f9c47192a04a423;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2e66e11c5cbc88f486e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105142cc1474502a590c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb370d6dc90d97408131;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf64a21a37cf32d17bbc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129721a41abc9e1a61107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e96710f109c6348bf30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1305bb421aaf5ca4d222a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1999a590ed2f78d723fba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e3fd2015e32ad9af29c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b131620e055745d52ef9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af678dd2967da1af0e51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4828d953e34e6be61222;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3078a23b67f01b420901;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7781e92bf5a3f0c4e86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc317325ca14bba9b6013;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147b6b7ad36e4bae245c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h576779d96019fd3bac4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebe2151c2451acc26508;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11963a6da0420ed31cf96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cd694d216f200a3835d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b50d442ba12c4e8026b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc77315b3912db5cc373;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h762b822510fd6224b08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e7580db6c2ccc1342ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5d075311a66412ff1af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd503494af0a54e0a1d54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79df374af43ba77b3ab0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2baf9a23793801eeef05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe291e01eae94ca07cc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1231f14987f7a32e9070a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1920b19636d741c840f9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9dca690dc06d23ea625;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd9eac4effa6b147e234;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf536b5116d093f230960;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19697490e2ad33a605410;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0106558ef2a3f8d9c91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69ccf6da85fa8f42f567;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1469c77237c978e734bfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10cf77247e5b38d0cd32d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fc409aa2fd2c603768d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2f8178a09636f37d81e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12054ff04146c2d1c6140;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa6901bb00c6fc0716a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h258aefc9ea7838b4c4da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf25dc0bda6d55bca6c08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h375125c7b96393aaac6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1919a25be7b1afc066d0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac5a1af701029357b2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8450595431ccef5d356;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eadbb928a5d9704a9b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1286571656d8cd1d111d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e0f739cd30e9b23e610;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bfdd283382ab1ee0017;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef2e960d4f6cbb6ad246;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11919dd114d986091648a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159a66e1f021a560bd0c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97c97d77066c18436e24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3e976413cc24a6cbc30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff6525f0393320549f57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba858b786c486e076318;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197016e5d9cc3441c200a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9e9e8390a1a0d0e4c05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146982b6da5cd0673ee3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb21462651ebca1135c87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc997513b2ac2dc97562;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d86563a4bee7a00d117;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24b8336b198b7108300a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5a29c702ef9b026a2bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15dfb73e176e4d32d2ce0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc99f33f17ea1d7cb204c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbf6a2bf61e3a95fedd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1998909ec1f8df76eb9e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba2909564a5331ed9a3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71c7fa2c5ca681c986;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5739e06b512c32a6529d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cf74f8a871c1ca4bbc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4123e6c93325e10b815;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cc32ffb2fccdfef3124;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89c8a180f8e27b47b58c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12191b5a437b074754b7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa05012056a9df0cf8d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1258d5976a1bb86187769;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ea3a74c7e3f6c4df14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81e642804e350a0aa84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbffc9715a82d33c6dea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d10225b88f66a8bb0a44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1528d53424c1c58da6645;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f9d17c6609c3a6adb32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165cd43dce778c4e05872;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h437e007fc2bbee5ab9e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5d21fb8ca4b75958e91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb445856161b9face06a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b65a6fb4b5a159cce8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9d4d74bc8280846b3d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5743fad729e18a575d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9292b8dd57a9a720635d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d62d6ca1a8f750c0335;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef7004968a135e10658;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154c6a05217b12e462f0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbe681c9cf78a5010dbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27df6acaf1b72268c274;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cea4247b579bcfcf8f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135c81e316420252b6aa1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13efe8277259d4b7ef03c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de04258cd67144b218e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfa149af17ca314d378b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dc904fd8e5a66117ee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd4d54dee9d84ec2b12b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h851970ef03f4d4cc26cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51c07d06627648e83fcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1951fb5cdc313ad555a02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1459633a9fe01119d1def;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f234f7de1494c95fca5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd79c0e4f6bd13865d44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1a07b22bd19aca62d1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d0fbfa106e459a4a7fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1389bf7105be32f84d1e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h836b8e65d4cf300c6ed7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dbfabb73088c6957f99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf61dd1af2f417fa1d6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h333f48bbade95bdcd49a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a23271e6b5e19e1a7721;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h153666d9f453f4c24be66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13aec910487292eb3e38f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5435445eab518c13b6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1fdc546fe32a87c292a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7bc3cca6cbd8c69b7bbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h541a4c3e762eda4aa0e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1662e1b2e9db8ae2fdff5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e5c5ada461f48331c23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bc804877a96e296d873;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a99d23a72af1b5cdcf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8fad87c9eefad8e8f155;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4cfe78a80b5da3a0210c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bda5cf779fbd77c53371;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6dca8ffd278d143eaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e4a4fbf1e235b0f311e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heea7860297a83cd295d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14973789c56a4c414365d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf01166b5872caa02eb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148284a107fec330e4bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3342971a1cc72e5f2d11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d640d0e6a0efd3aaf696;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14318298c54492f6bf31c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8976b3dc98b7856a6927;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha556c72aab962df345c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f211eb40ab88d3887b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5a14e03a542d2d1c5a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4eeceea8cc112d8d3de0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d04d74d6a83eef9cb0cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf470ffae57c510e10ffe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccd889328f6f10d8dafa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he27acbe2d31dd5774c75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c3641dc2e4a550776c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb2d7f7992cc7388fb21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14789cc40a5eff361e47c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39de1518a54620a16b5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab67465e48e81007ad1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc50c618557209b490724;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13668ffc46a5df8fc875f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1e435909c61b256d00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h122b35ea080e3e6ff8bb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102ee3f86cef724340911;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13be21b64784acb682ea0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h349529931f56ad56c2e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12836726b24551b6187a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haded9a647aa096a60fab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e897b57b99f0c583e48e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf738c1cb0ff32b0fba2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f60d9c88ba27db83113;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c05bf9977c8d4f67990;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1675a7394f85857f4c721;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf47a3874f97a963faee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedf82dcbb1720787bd10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140ab4eadf48c349558e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9d930df0f0e84af7c76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d43966283f8561ed3bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7c97e0d155cb768577d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a7a8c41642934e28cff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8fd25e9532415593348;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca47f0e6616eddd57b25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f79474685267d123763;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1251b8111a54960332c8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c7704e5f97ca9ee22eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce0de496ae5139c56f81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af5cda1f980f67dbc236;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e5e2af79bfb2d08d879;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119437daad476479c89d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bb8cf562263d3396598;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cdaa4afdcdb98184a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd021aa982964107aad3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c43f113ccbd668cabb8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e0a105d0ffde880e0ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114a2ad597d7c8204b705;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2228c00eb35dee8c12e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ad7c8e255ba7f35a0d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78cc0a6c40e05f696233;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcebf7a0b0a78bf0239ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87b9e5e530e85effeba9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190ee41087a3eb5c7039;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfa0b101bcdda2692c1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7d8ade431b33d3028e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f6b58eb17e6fa900c09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe0ae0da3d193131d3ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b44814237bcd80ecd945;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1f0b688905acab17412;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ebafbe95e68095b722e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa7489caf2bfb535757;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81950cd3f40f270878b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4153ab8c8f82c6d4a2ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eacd6b9ad01a1e2d033;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a89d19b461964153cfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2968ec0e4a9608935d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1036e08ec6879e28ccaee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23d1c9eb95811b62a960;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdf4fc614d2846f8b727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119b77e3bde3e10917f58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1550a00d4383113b7bc74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e234eab5901f453df206;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc279c2d22ff4877fb617;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12145badcb14c4ae0138c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cba497b4a03f40fe1ece;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1ec2445e7ec25d11a79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b223a698a36d9080deb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de52da54ceab524849de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2967441eb5dda368d777;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3208b225df6b67fe8802;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e2062c26fb6d8aa72af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7cf1d67feba3222c028;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb40b129fb51bcab52277;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1700b4d04c3b64ce93846;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a3deb86e30e0136ff1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac6de79154350bce0bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h973e338cd6d0ed7d215f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e0368cb801aa544ec8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfef5a10712ea6bf40a3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1291ce0e21fa6f3f9968e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124bb7789065abf8fb9aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c864b3d36d68844bab8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133236b49fdf435c2be97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffa35da33638019df477;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8d2684571bf404080aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168b96571fa964564509f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74f0b6cd6408be47d52a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12450b9c795a4fdd811af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42546ec3800a5bf70e94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ec5f82bc2dcb63d4f32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199e2d08c8b1be66374a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c3703c7516a799d447f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h207be7720fd4930e2260;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7710b4a3349bb0a77213;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2dce5c467aa31bd4c4c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3859e9182f8ea51f8041;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bb8270013e9d564e4e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121f1555bea18f8531d31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f150caace68498785cec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he587418515f821a9216c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2aeb83706a6818a835c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79334e4f7497a041c6cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafbf7fa88607f6a5a6df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcbf4779fc989f9c38d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be148c5b5e175b7c44ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbce02365e80303a4e4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1020f5a7059eec55ded68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cddf88b29382934f0836;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131034255c735a828abdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha252fb00243d725dc2a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f436f95c314d50a0715;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha29d5f2b1ae008abc040;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c1b75bbb96b33901642;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab0f5e2ea6bf649a6e83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1297acb7a6acff9a7398b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d7040dd25c108672421;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73fab3ab59bf7010746;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h533ad91d461b6c6d89f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1450bf3d7e58a42ecf4a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hceffade1fad2075e468b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f07ac3a5eb7259f36d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb72425cfdec82cc07a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aaefa63c60379acc30d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa5cffb0e37cfd74c6ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3a91d2fd8114bac5b9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123ca3d90eb904d54f567;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb4f4990cbaed610e4ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cfc80c617f875e73adc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19548b9d4da31f3821da1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103139324e9e7285d5642;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157bd37d2f6383c40b0ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16184516d550946c68b59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6414a4232a0d536dd76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1971de390ff1a4acc5bc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d4755ba63fd36f50190;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16683d0bc42adfff1dc6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0624b8b833e374584d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb483af03072f93e4bfba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4fb7e583ee515db847d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb68a85141afd058ba5a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5d899a172a5458c2e62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7cd1b88ce0f9f4cac17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130c005e9f17e14af30d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7de6c0206b799fd504e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10749c135cdfbbd6ea1c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162882bc8d59022fd7a42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141105dd8d9dd2936ab31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81cdca9cb6295fb8aeb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45785c5c8bcbda21d124;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea1172914095863fa194;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53a5ae3d43a229b2160e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h471f3f21e461dbaeae72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87b5f3f847a5ff64af31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d93ec575ae4e87dc4db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e522fcc809f6978a9048;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177f0b5f34b47082876f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18733dcc5cfb5d4598ca4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fbdb60f90225bc0a986;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e6a9b890de8370dd49c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be4d9736f04e2fd171d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d965ef1a53e4884c48b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb57568466ac47bbcdfba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d470195c36b2994b3188;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee44165e19b6c95738de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44b81d5d9e7fd60c0402;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3c407bc8eefa5ff5f41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h281ee26c26bb88338416;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51a7fee376c24c324569;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11154ef2bc7ce8b863c13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc34b46a6585ee84ab08f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h781eacb85207b326c3b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef16f67e42c285cd9712;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0b6b4b7747f623e0096;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135df177f1479eea4053f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1390a4b755e156a8d84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ef23c9d35ed7d952458;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1800bd08c8c4d577700b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e337c78c40d21b0c449e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd86ef18a86798b0ebb49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d44d9c15f402884993cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f589e66aa0ce8acdfa10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c2d909a6787f6c380da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h807e78df709c06526a85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b7d1cbff3281843acd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h946bb557a91148ab7b5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115e3032570e3424fcdbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b71caa4cbbe3f8f62cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b7364fb1bd46c6af61f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76f772f20246d3313778;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c3ad6de7fffc0c46384;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14adf3e38fed3e257ef6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2f38fd9ae1fd433dc57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b83c51f731183ff1710;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6626106564d25e1bccf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b5315d32cfb7a7341e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h850f8cfd5ca3e9d4f128;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143c71b72a026cbeddf2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19619ca6eeca537d3a9ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef6c4cb6244d3c804256;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c9294c03a1c1025fec8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa3b353be82ea5b76da2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6654e754468e54fcb344;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fbe08971385fd455f84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3439dd536484aad89d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150335b84b330a60c65b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2623de637cda48a06e91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h809186a608e24feb6656;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c566d35a11e31433235;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9e3e1c95c028bf0e3c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9d900f7099da8de2827;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bccac1ef37f54653816e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90d655444ea633a0b1a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf18ffb4d31cff784fb14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h444ab5fbfbed7f8b7372;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cecd261c2f5202011a97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cc6a00840156df3e14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4bbb881b1dd720b6caa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30b31eac7171e23fd162;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h593d7087194118f93244;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac00f58a94df4a46590f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18abce9615b9d2ee0fe7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96a022832d6f32732abf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f87338d277ba93a5d27f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6954354695ad4cb7f04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c503e734868561b26ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f2a62add78919202264;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d64fd12b70b62368b0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7de924a0a61b2fe57db1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193c5cf1f61abfe2f58af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f807153200d01d4ba6c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad4e6345eaa3a2993cf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5282540b73955f0c4b67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fd2f5958501eaade22c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfdaee67c0ff2518c614;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf2e599e214cc43f5e1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d5e202c9ab493004d9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c91ed82f734f285d7aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb25afecd19a80c32ac0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ee906fd9e732487cd4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1944ef2de95a508da7c61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6b32102f281f36d9458;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ee75f44ab48484ec2d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1742bae42b461eb14cdee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13de24bbdbf39bf711f63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fdc5b0d40b1bf620fe3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12dea2cbe6f6515505344;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa83389c5901d9ac35b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e277c3d2a5fd7c532c6c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a6ac69f9ec2a9c201a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a54c7067533de8ae6f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1358230e497ee56634fd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1754b388a0785b819eaff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1852a8a772af0c29be4b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3bcf201959bdd3c8292;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41c76422aa3e0a7296ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3221857faebeb20ff8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e1e9bddbf138ec02c7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff46590ed33d461b3f46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca8149b8b66bb849983;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h293cead13cd36e3ae40e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb004b9d38ac6078a5dc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffa3ff967b5dd5352c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c296490880b9c47cc84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192867c60feabcd2f2e2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16095f9aab304b1b3a29e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2208238b5bce8e641aed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f26312cda05646393ce3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db286898554e8ffea996;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3a8a9997b0e4bd64b3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68fcc195093176fcfef3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa5ab58cdf3c54a8ed7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106215124b5926c68a57a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17fce00b6e10c81afa039;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc888ef8652db0b82ffad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157e2876d313d4fc39aa5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h825d22bc976e1673d89d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fbfdf0d1d4f42bfe6ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18dd80b09d8a14367bdb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba206c6c3f2f5e1e324d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h259f70c3a5c1e68f762b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h740c4f20d57843cc794d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59dcf62cb218058e8228;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c010df44fc957b9ba13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e768bdcebc0ba74359a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86e748a0cc41a0ba18cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178daa11f72b7716964a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148549dbe502c4bbe3d93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h470c67b9a19384e9901b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafebaaec2ff5d3491ed1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19453d7b5999471c7baed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d3da2040c28e84fe6d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccec275a5704e2bc4a98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a655b50c8943bf09626;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17af1754faa3f6ef05b13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0dc37909833c8a39e1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e57b222d6e66fbf29c59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cf59f7bb2d2219405fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15789c8b5d004a2551733;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d4fdc07f434534ca0e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42917a1f3a0267ac7184;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2aaea2ae30420f73c24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h680495d67ddb10446ad0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc29472c9eccb0393dbf7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a31c5be385118a3ca3f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21cc7e6be764a79ab2fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7a219032e44e8cb2de7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1740f934427ff9903da9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af43925db2555728414d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4b1eae65c62a2cbc2f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c68eb4fb2846c883403c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d03ad862345e6dd0126f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1daae39fd101fcbbadf9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c752f7ad0752dd08aaa4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbcf0c3dd3e786801d09f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182569282cc9b54b357ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af04012f2d0cefba0291;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf35fe6178ecb62e6c807;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1458ce785817e7d58eaa9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6e6a07fb6ebdb830055;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f536a892d5a01f6997d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h440403dccd68ad245218;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1188250c5ae417f0d450a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12784304a03836a933f1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec4924a1ed180bc67cdc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be53044f68d537e9f816;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94fe61c954049897a501;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a7c17301b04eb71c750;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cd96803217d5e36de1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5127b4eb293fe8dbbfc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178b0ae7993a9ffcbb76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1524889d0b44440fc821d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10bd97f51a3079aab1ede;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3caf1291573a01338a12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169bbbf7baefadaf3503d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130328364257aac55bf38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d78c27ca9c544cb96b0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebcea9732786c8c75bd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118ce52a03ad471b31fbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f59621aa209bfaad600;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddbf2bf48cdebf89b4e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h678af14c30afbf71155e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159f845c53da67f27b72e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93d00b8a152ff4ec9bfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8bed42f4977486459bd5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bd754a59688d817b9b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193cd7e572fa3407bc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17bfdbd48bc5da5cdd681;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb936dbf020eb0977c3c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c18cd1847a4e93cb0579;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd02c6f6795ade74e6d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ba5a5227775b63761fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4a9b87630efcb314f4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119e492b9bef7540d4f79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150fa3205d98cd32df1f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2ab68d41c05ad772e98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1000b04eb8c9d61e809a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6317cc78f94eda52d83f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9f7116c13306d6942c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1784908ffa2b571611b5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec2bb3940468bb79825a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd6d2f8828d2d1c447d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h857984bf59cf791de008;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b305f89f6635075c3014;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10faaf76d1fac69f013d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c8f94a7b8b5b0947bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86c3e93d98a848680e8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he312ec2852100125794b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42db635a442dd4c84a7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64a90f373e06fb800483;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5cf9df7e71c2e4cd5895;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18978dae10d99458ccea8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1236b0f0ab28097ca705b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c61c867fe23dbc160e05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1e5908a1eda3b3fa94f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92a490f4854061a8d56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3171978652a1df9f69aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0fd827e759f5845351c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h883ef0826d3f422395b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha36bf2ee23f46c7e69ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6af2f77ef9aac0892698;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5381337ece504f41fb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bb7fb1c31cde71fc304;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1383842a2424e46be9e09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e204b583e17ce4365c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc98acbc9fe196b83a47a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba841045029f2abc9c5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17bd352277388f89c23af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1044c42b8bbd2390bc107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb9a2a67845d81be253b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h616aafc64f6178da7920;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15aaa40418bfa9c191b18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1687fa4c8a4e60310954c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a491313f08cefcbe0db6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8ee011e2546e72e7a75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2a8caf584ee51940e7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95b70969ddfe03c2032f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf98f7ba2714c1b1dcbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d469c231a7cdef7800f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h898162a539cd8bafff2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h845beab8e5ecbe6a1864;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c8f43e483857cf3460a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11af04c3990f4ce8f0c50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6241e7c41c236af170fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha52cf254aaa0ea4e2977;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h847658866b43f1581a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f5a419e8995dfaef0bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac10d758a1efc765a40b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de9e54c2e8bac9ae67d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152aa0445a62eeded4d9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ecbd836aefd13a05caf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfb9b3240f67fcab57ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c88a506990f37ad6256;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137de03a8f56d17c5920c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf3bde34a05e7b6b47d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177ad99f7c8fcb57abb95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb77ebee707b2bbf7987;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143b66203c13d1684b0a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4a2b7394a693611d26f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h971a7708ad98c859d1cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129da34e0bba341efe333;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdf4dae691c1d412e428;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h693bf0e44d888b4d7dea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2701bd3b6055fd3d7d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1277caddb19ddff88251c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57be7f4d8ef879755cc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3eb977297d0acc5f36d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3c4155d450f9ade8b7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1011bf0db96bc79c2c612;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc355e1556eafe3295fab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba0aa2a24fe6403a97d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha39ccb442803b0eda19d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4de20e37395463d9fa9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6c659b4c101dfd3f156;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2aed5ccc79f7545cdb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6bf9891004c65856b43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177c7e2dc6c39f0180a1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9ae3924a5458ea12a2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32cb4c3a2ed53a21adc9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdaf5cb09559909813d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h780d188c9b99b1b80a1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b871e494850dce30ff1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188d2a9cc0d1d966d9ca0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10529812778580380eea2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4210adbcc6a98556a37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f37852ef09cd48d4823;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1596da9fe79c18a92c485;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d4186964bfc810ff309;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e8a2b270638d46f714c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f48135551bf634a4923;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c735e9e17b229c502985;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154ea203360b1db52603e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8be36cf2aec3d27eccf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h584273791d1df1f0b309;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144449357c55fc51f4c6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfafe9236c6beb555605;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19493cc2f6b784ff42921;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13189496df0332f43e73b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198045f7bfdbddd76c2cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff7e0880ec6accaff00e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a062e9913f97b2d1d60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd135b56bb12e188dd7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ded67afd03a9c862fece;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4c562b2bf38a688b8e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b799de0371e885765c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3b453f2c71ca82138fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76ec6e1f2ff69a33b9bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18957425f4c6782a1b909;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f0437fb622596ee9113;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d18d203cd018c4e376f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1111c3563bd512ca2d627;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12836daa82ba41361a163;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb50d5d96f9912020a68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce5d752b76b53eded6fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175773c58553669916b28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ea8833861c5560c722e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hccd9f94ef07fd395f27e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39f5d343b6cc960931ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18251eea594b6ccfbcd22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba773ddbe548b338aaaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a3e512402ffe05d6953;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179d840dd173f0cff5384;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e65c1d0f7e022eaaa5bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1467b5bab02e71e6799e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144b1b7e1660e0226e38c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186203781d210a431035;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h396289718c9e209c3c28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h297194f1d2434029ac5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cedfc5bacc3c4c7dc7b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1055935363b72a62fc2b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa42622baea7601879c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha69d39869599d182c053;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11bb71a706035a341742;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3021a0dfc4d87850c58a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc470252fccfbb9cbc711;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d03bb03bc05a45148e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ec964b31969e0deecf9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf654be84b9b2c56dfefb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1584806716368f63f8bf4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d830e1327e3c29c09642;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185208e05e03499a0e58c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c114f026200818c6e2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42f8364562283148c45b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d7a02666a16148f570e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c440242b054f26d79505;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12935701c718b2be79d62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8ee6204312f30569da5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf6abcf8ac969e8df175;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1937574e252b19ceeac31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106474b7de99b13608c02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c09919d765b764c1243f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5ff59be9d5d036acddd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha31a473c0c167b666297;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8d657a40c7b4b9adeef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fc0405b0c49c50a21e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5b168d26a4180b836a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc84b2903ac7cd2fc694;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8e57be179779f25b1a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7ca8047f73816c84fce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9890ad856d946ad3ebf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h205c2cb6b5aacf59c5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c8ca2aab97bfe756d75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8fa0cecbf7c02bc81a07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdfc212ed6d86bef9f6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2f75c1ae190b6c69732;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3c1e4f6f8bdc40bdcdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21d87fdb3a1517e9a45e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4c4edbd8863e99f7138;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c25ece52378dc3411b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6df54a6e19a189107266;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d170dea97671ed0d6b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h335e6ba3d24143ee3a42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a20b006ae452f7ee72e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb38c471fa120f14e81d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8935ed1987baf1bb37b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1851aa0f6e331ca3d62fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca3c8ad71b0d39b5d659;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he45473c21c490e36eac8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d72c65c8460849ffefdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104af67b57dfbae6f651f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdc431593e31139387d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e390d6e18b2d9411399;
        #1
        $finish();
    end
endmodule
