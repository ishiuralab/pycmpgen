module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    compressor_CLA128_16 compressor_CLA128_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA128_16(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [45:0] stage1_0;
   wire [63:0] stage1_1;
   wire [38:0] stage1_2;
   wire [48:0] stage1_3;
   wire [59:0] stage1_4;
   wire [56:0] stage1_5;
   wire [47:0] stage1_6;
   wire [64:0] stage1_7;
   wire [55:0] stage1_8;
   wire [57:0] stage1_9;
   wire [53:0] stage1_10;
   wire [51:0] stage1_11;
   wire [56:0] stage1_12;
   wire [71:0] stage1_13;
   wire [70:0] stage1_14;
   wire [37:0] stage1_15;
   wire [35:0] stage1_16;
   wire [20:0] stage1_17;
   wire [14:0] stage2_0;
   wire [13:0] stage2_1;
   wire [19:0] stage2_2;
   wire [19:0] stage2_3;
   wire [27:0] stage2_4;
   wire [27:0] stage2_5;
   wire [16:0] stage2_6;
   wire [30:0] stage2_7;
   wire [28:0] stage2_8;
   wire [20:0] stage2_9;
   wire [17:0] stage2_10;
   wire [37:0] stage2_11;
   wire [28:0] stage2_12;
   wire [18:0] stage2_13;
   wire [34:0] stage2_14;
   wire [26:0] stage2_15;
   wire [19:0] stage2_16;
   wire [19:0] stage2_17;
   wire [6:0] stage2_18;
   wire [1:0] stage2_19;
   wire [14:0] stage3_0;
   wire [8:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [8:0] stage3_4;
   wire [9:0] stage3_5;
   wire [10:0] stage3_6;
   wire [8:0] stage3_7;
   wire [13:0] stage3_8;
   wire [12:0] stage3_9;
   wire [7:0] stage3_10;
   wire [16:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [15:0] stage3_14;
   wire [10:0] stage3_15;
   wire [19:0] stage3_16;
   wire [6:0] stage3_17;
   wire [5:0] stage3_18;
   wire [5:0] stage3_19;
   wire [0:0] stage3_20;
   wire [5:0] stage4_0;
   wire [9:0] stage4_1;
   wire [2:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [4:0] stage4_5;
   wire [3:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [5:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [5:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [2:0] stage5_2;
   wire [6:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [0:0] stage5_6;
   wire [4:0] stage5_7;
   wire [1:0] stage5_8;
   wire [6:0] stage5_9;
   wire [0:0] stage5_10;
   wire [4:0] stage5_11;
   wire [1:0] stage5_12;
   wire [6:0] stage5_13;
   wire [0:0] stage5_14;
   wire [4:0] stage5_15;
   wire [5:0] stage5_16;
   wire [5:0] stage5_17;
   wire [2:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [0:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc606_5 gpc18 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc606_5 gpc19 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc606_5 gpc20 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20]}
   );
   gpc606_5 gpc21 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage1_5[4],stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21]}
   );
   gpc606_5 gpc22 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[5],stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[6],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[7],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[8],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[9],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[10],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[11],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[12],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[13],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[14],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[15],stage1_4[32],stage1_3[32],stage1_2[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[16],stage1_4[33],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[17],stage1_4[34],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[18],stage1_4[35],stage1_3[35],stage1_2[35]}
   );
   gpc615_5 gpc36 (
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage0_3[91]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[19],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc615_5 gpc37 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[30]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[5],stage1_5[20],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[31]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[6],stage1_5[21],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[32]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[7],stage1_5[22],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[33]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[8],stage1_5[23],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[34]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[9],stage1_5[24],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage0_4[35]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[10],stage1_5[25],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[6],stage1_6[11],stage1_5[26],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[7],stage1_6[12],stage1_5[27],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[8],stage1_6[13],stage1_5[28],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[9],stage1_6[14],stage1_5[29],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[10],stage1_6[15],stage1_5[30],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[11],stage1_6[16],stage1_5[31],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[12],stage1_6[17],stage1_5[32],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[13],stage1_6[18],stage1_5[33],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[14],stage1_6[19],stage1_5[34],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[15],stage1_6[20],stage1_5[35],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[16],stage1_6[21],stage1_5[36],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[17],stage1_6[22],stage1_5[37],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[18],stage1_6[23],stage1_5[38],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[19],stage1_6[24],stage1_5[39],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[20],stage1_6[25],stage1_5[40],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[21],stage1_6[26],stage1_5[41]}
   );
   gpc606_5 gpc59 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[22],stage1_6[27],stage1_5[42]}
   );
   gpc606_5 gpc60 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[23],stage1_6[28],stage1_5[43]}
   );
   gpc606_5 gpc61 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[24],stage1_6[29],stage1_5[44]}
   );
   gpc606_5 gpc62 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[25],stage1_6[30],stage1_5[45]}
   );
   gpc606_5 gpc63 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[26],stage1_6[31],stage1_5[46]}
   );
   gpc606_5 gpc64 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[27],stage1_6[32],stage1_5[47]}
   );
   gpc606_5 gpc65 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[28],stage1_6[33],stage1_5[48]}
   );
   gpc606_5 gpc66 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[29],stage1_6[34],stage1_5[49]}
   );
   gpc606_5 gpc67 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[30],stage1_6[35],stage1_5[50]}
   );
   gpc606_5 gpc68 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[31],stage1_6[36],stage1_5[51]}
   );
   gpc606_5 gpc69 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[32],stage1_6[37],stage1_5[52]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[90]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[33],stage1_6[38],stage1_5[53]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[91]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[34],stage1_6[39],stage1_5[54]}
   );
   gpc615_5 gpc72 (
      {stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_6[92]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[35],stage1_6[40],stage1_5[55]}
   );
   gpc615_5 gpc73 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_6[93]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[36],stage1_6[41],stage1_5[56]}
   );
   gpc606_5 gpc74 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[16],stage1_8[31],stage1_7[37],stage1_6[42]}
   );
   gpc606_5 gpc75 (
      {stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[17],stage1_8[32],stage1_7[38],stage1_6[43]}
   );
   gpc606_5 gpc76 (
      {stage0_6[106], stage0_6[107], stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[18],stage1_8[33],stage1_7[39],stage1_6[44]}
   );
   gpc606_5 gpc77 (
      {stage0_6[112], stage0_6[113], stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[19],stage1_8[34],stage1_7[40],stage1_6[45]}
   );
   gpc615_5 gpc78 (
      {stage0_6[118], stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122]},
      {stage0_7[96]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[20],stage1_8[35],stage1_7[41],stage1_6[46]}
   );
   gpc615_5 gpc79 (
      {stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127]},
      {stage0_7[97]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[21],stage1_8[36],stage1_7[42],stage1_6[47]}
   );
   gpc615_5 gpc80 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[36]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[6],stage1_9[22],stage1_8[37],stage1_7[43]}
   );
   gpc615_5 gpc81 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[7],stage1_9[23],stage1_8[38],stage1_7[44]}
   );
   gpc606_5 gpc82 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[8],stage1_9[24],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[9],stage1_9[25],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[10],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[11],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[12],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[13],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[14],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[15],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[16],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[17],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[18],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[19],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[20],stage1_9[36],stage1_8[51]}
   );
   gpc615_5 gpc95 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_9[12]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[21],stage1_9[37],stage1_8[52]}
   );
   gpc615_5 gpc96 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_9[13]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[22],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc97 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[15],stage1_11[17],stage1_10[23],stage1_9[39]}
   );
   gpc606_5 gpc98 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[16],stage1_11[18],stage1_10[24],stage1_9[40]}
   );
   gpc606_5 gpc99 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[17],stage1_11[19],stage1_10[25],stage1_9[41]}
   );
   gpc606_5 gpc100 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[18],stage1_11[20],stage1_10[26],stage1_9[42]}
   );
   gpc606_5 gpc101 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[19],stage1_11[21],stage1_10[27],stage1_9[43]}
   );
   gpc606_5 gpc102 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[20],stage1_11[22],stage1_10[28],stage1_9[44]}
   );
   gpc606_5 gpc103 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[21],stage1_11[23],stage1_10[29],stage1_9[45]}
   );
   gpc606_5 gpc104 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[22],stage1_11[24],stage1_10[30],stage1_9[46]}
   );
   gpc606_5 gpc105 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[23],stage1_11[25],stage1_10[31],stage1_9[47]}
   );
   gpc606_5 gpc106 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[24],stage1_11[26],stage1_10[32],stage1_9[48]}
   );
   gpc606_5 gpc107 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[25],stage1_11[27],stage1_10[33],stage1_9[49]}
   );
   gpc606_5 gpc108 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[26],stage1_11[28],stage1_10[34],stage1_9[50]}
   );
   gpc606_5 gpc109 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[27],stage1_11[29],stage1_10[35],stage1_9[51]}
   );
   gpc606_5 gpc110 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[28],stage1_11[30],stage1_10[36],stage1_9[52]}
   );
   gpc606_5 gpc111 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[29],stage1_11[31],stage1_10[37],stage1_9[53]}
   );
   gpc606_5 gpc112 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[30],stage1_11[32],stage1_10[38],stage1_9[54]}
   );
   gpc606_5 gpc113 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[31],stage1_11[33],stage1_10[39],stage1_9[55]}
   );
   gpc606_5 gpc114 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[32],stage1_11[34],stage1_10[40],stage1_9[56]}
   );
   gpc606_5 gpc115 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[33],stage1_11[35],stage1_10[41],stage1_9[57]}
   );
   gpc606_5 gpc116 (
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[19],stage1_12[34],stage1_11[36],stage1_10[42]}
   );
   gpc606_5 gpc117 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[20],stage1_12[35],stage1_11[37],stage1_10[43]}
   );
   gpc615_5 gpc118 (
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106]},
      {stage0_11[114]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[21],stage1_12[36],stage1_11[38],stage1_10[44]}
   );
   gpc615_5 gpc119 (
      {stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111]},
      {stage0_11[115]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[22],stage1_12[37],stage1_11[39],stage1_10[45]}
   );
   gpc615_5 gpc120 (
      {stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116]},
      {stage0_11[116]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[23],stage1_12[38],stage1_11[40],stage1_10[46]}
   );
   gpc615_5 gpc121 (
      {stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121]},
      {stage0_11[117]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[24],stage1_12[39],stage1_11[41],stage1_10[47]}
   );
   gpc606_5 gpc122 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[6],stage1_13[25],stage1_12[40]}
   );
   gpc606_5 gpc123 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[7],stage1_13[26],stage1_12[41]}
   );
   gpc606_5 gpc124 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[8],stage1_13[27],stage1_12[42]}
   );
   gpc606_5 gpc125 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[9],stage1_13[28],stage1_12[43]}
   );
   gpc606_5 gpc126 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[4],stage1_14[10],stage1_13[29],stage1_12[44]}
   );
   gpc606_5 gpc127 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[5],stage1_14[11],stage1_13[30],stage1_12[45]}
   );
   gpc606_5 gpc128 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[6],stage1_14[12],stage1_13[31],stage1_12[46]}
   );
   gpc606_5 gpc129 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[7],stage1_14[13],stage1_13[32],stage1_12[47]}
   );
   gpc606_5 gpc130 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[8],stage1_14[14],stage1_13[33],stage1_12[48]}
   );
   gpc606_5 gpc131 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[9],stage1_14[15],stage1_13[34],stage1_12[49]}
   );
   gpc606_5 gpc132 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[10],stage1_14[16],stage1_13[35],stage1_12[50]}
   );
   gpc606_5 gpc133 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[11],stage1_14[17],stage1_13[36],stage1_12[51]}
   );
   gpc606_5 gpc134 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[12],stage1_14[18],stage1_13[37],stage1_12[52]}
   );
   gpc606_5 gpc135 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[13],stage1_14[19],stage1_13[38],stage1_12[53]}
   );
   gpc606_5 gpc136 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[14],stage1_14[20],stage1_13[39],stage1_12[54]}
   );
   gpc606_5 gpc137 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[15],stage1_15[15],stage1_14[21],stage1_13[40]}
   );
   gpc606_5 gpc138 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[16],stage1_15[16],stage1_14[22],stage1_13[41]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[17],stage1_15[17],stage1_14[23],stage1_13[42]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[18],stage1_15[18],stage1_14[24],stage1_13[43]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[19],stage1_15[19],stage1_14[25],stage1_13[44]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[20],stage1_15[20],stage1_14[26],stage1_13[45]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[21],stage1_15[21],stage1_14[27],stage1_13[46]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[22],stage1_15[22],stage1_14[28],stage1_13[47]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[23],stage1_15[23],stage1_14[29],stage1_13[48]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[24],stage1_15[24],stage1_14[30],stage1_13[49]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[25],stage1_15[25],stage1_14[31],stage1_13[50]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[26],stage1_15[26],stage1_14[32],stage1_13[51]}
   );
   gpc615_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76]},
      {stage0_14[90]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[27],stage1_15[27],stage1_14[33],stage1_13[52]}
   );
   gpc615_5 gpc150 (
      {stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_14[91]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[28],stage1_15[28],stage1_14[34],stage1_13[53]}
   );
   gpc615_5 gpc151 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86]},
      {stage0_14[92]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[29],stage1_15[29],stage1_14[35],stage1_13[54]}
   );
   gpc615_5 gpc152 (
      {stage0_13[87], stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91]},
      {stage0_14[93]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[30],stage1_15[30],stage1_14[36],stage1_13[55]}
   );
   gpc615_5 gpc153 (
      {stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95], stage0_13[96]},
      {stage0_14[94]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[31],stage1_15[31],stage1_14[37],stage1_13[56]}
   );
   gpc615_5 gpc154 (
      {stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_14[95]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[32],stage1_15[32],stage1_14[38],stage1_13[57]}
   );
   gpc615_5 gpc155 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106]},
      {stage0_14[96]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[33],stage1_15[33],stage1_14[39],stage1_13[58]}
   );
   gpc615_5 gpc156 (
      {stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_14[97]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[34],stage1_15[34],stage1_14[40],stage1_13[59]}
   );
   gpc615_5 gpc157 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116]},
      {stage0_14[98]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[35],stage1_15[35],stage1_14[41],stage1_13[60]}
   );
   gpc1_1 gpc158 (
      {stage0_0[99]},
      {stage1_0[17]}
   );
   gpc1_1 gpc159 (
      {stage0_0[100]},
      {stage1_0[18]}
   );
   gpc1_1 gpc160 (
      {stage0_0[101]},
      {stage1_0[19]}
   );
   gpc1_1 gpc161 (
      {stage0_0[102]},
      {stage1_0[20]}
   );
   gpc1_1 gpc162 (
      {stage0_0[103]},
      {stage1_0[21]}
   );
   gpc1_1 gpc163 (
      {stage0_0[104]},
      {stage1_0[22]}
   );
   gpc1_1 gpc164 (
      {stage0_0[105]},
      {stage1_0[23]}
   );
   gpc1_1 gpc165 (
      {stage0_0[106]},
      {stage1_0[24]}
   );
   gpc1_1 gpc166 (
      {stage0_0[107]},
      {stage1_0[25]}
   );
   gpc1_1 gpc167 (
      {stage0_0[108]},
      {stage1_0[26]}
   );
   gpc1_1 gpc168 (
      {stage0_0[109]},
      {stage1_0[27]}
   );
   gpc1_1 gpc169 (
      {stage0_0[110]},
      {stage1_0[28]}
   );
   gpc1_1 gpc170 (
      {stage0_0[111]},
      {stage1_0[29]}
   );
   gpc1_1 gpc171 (
      {stage0_0[112]},
      {stage1_0[30]}
   );
   gpc1_1 gpc172 (
      {stage0_0[113]},
      {stage1_0[31]}
   );
   gpc1_1 gpc173 (
      {stage0_0[114]},
      {stage1_0[32]}
   );
   gpc1_1 gpc174 (
      {stage0_0[115]},
      {stage1_0[33]}
   );
   gpc1_1 gpc175 (
      {stage0_0[116]},
      {stage1_0[34]}
   );
   gpc1_1 gpc176 (
      {stage0_0[117]},
      {stage1_0[35]}
   );
   gpc1_1 gpc177 (
      {stage0_0[118]},
      {stage1_0[36]}
   );
   gpc1_1 gpc178 (
      {stage0_0[119]},
      {stage1_0[37]}
   );
   gpc1_1 gpc179 (
      {stage0_0[120]},
      {stage1_0[38]}
   );
   gpc1_1 gpc180 (
      {stage0_0[121]},
      {stage1_0[39]}
   );
   gpc1_1 gpc181 (
      {stage0_0[122]},
      {stage1_0[40]}
   );
   gpc1_1 gpc182 (
      {stage0_0[123]},
      {stage1_0[41]}
   );
   gpc1_1 gpc183 (
      {stage0_0[124]},
      {stage1_0[42]}
   );
   gpc1_1 gpc184 (
      {stage0_0[125]},
      {stage1_0[43]}
   );
   gpc1_1 gpc185 (
      {stage0_0[126]},
      {stage1_0[44]}
   );
   gpc1_1 gpc186 (
      {stage0_0[127]},
      {stage1_0[45]}
   );
   gpc1_1 gpc187 (
      {stage0_1[96]},
      {stage1_1[32]}
   );
   gpc1_1 gpc188 (
      {stage0_1[97]},
      {stage1_1[33]}
   );
   gpc1_1 gpc189 (
      {stage0_1[98]},
      {stage1_1[34]}
   );
   gpc1_1 gpc190 (
      {stage0_1[99]},
      {stage1_1[35]}
   );
   gpc1_1 gpc191 (
      {stage0_1[100]},
      {stage1_1[36]}
   );
   gpc1_1 gpc192 (
      {stage0_1[101]},
      {stage1_1[37]}
   );
   gpc1_1 gpc193 (
      {stage0_1[102]},
      {stage1_1[38]}
   );
   gpc1_1 gpc194 (
      {stage0_1[103]},
      {stage1_1[39]}
   );
   gpc1_1 gpc195 (
      {stage0_1[104]},
      {stage1_1[40]}
   );
   gpc1_1 gpc196 (
      {stage0_1[105]},
      {stage1_1[41]}
   );
   gpc1_1 gpc197 (
      {stage0_1[106]},
      {stage1_1[42]}
   );
   gpc1_1 gpc198 (
      {stage0_1[107]},
      {stage1_1[43]}
   );
   gpc1_1 gpc199 (
      {stage0_1[108]},
      {stage1_1[44]}
   );
   gpc1_1 gpc200 (
      {stage0_1[109]},
      {stage1_1[45]}
   );
   gpc1_1 gpc201 (
      {stage0_1[110]},
      {stage1_1[46]}
   );
   gpc1_1 gpc202 (
      {stage0_1[111]},
      {stage1_1[47]}
   );
   gpc1_1 gpc203 (
      {stage0_1[112]},
      {stage1_1[48]}
   );
   gpc1_1 gpc204 (
      {stage0_1[113]},
      {stage1_1[49]}
   );
   gpc1_1 gpc205 (
      {stage0_1[114]},
      {stage1_1[50]}
   );
   gpc1_1 gpc206 (
      {stage0_1[115]},
      {stage1_1[51]}
   );
   gpc1_1 gpc207 (
      {stage0_1[116]},
      {stage1_1[52]}
   );
   gpc1_1 gpc208 (
      {stage0_1[117]},
      {stage1_1[53]}
   );
   gpc1_1 gpc209 (
      {stage0_1[118]},
      {stage1_1[54]}
   );
   gpc1_1 gpc210 (
      {stage0_1[119]},
      {stage1_1[55]}
   );
   gpc1_1 gpc211 (
      {stage0_1[120]},
      {stage1_1[56]}
   );
   gpc1_1 gpc212 (
      {stage0_1[121]},
      {stage1_1[57]}
   );
   gpc1_1 gpc213 (
      {stage0_1[122]},
      {stage1_1[58]}
   );
   gpc1_1 gpc214 (
      {stage0_1[123]},
      {stage1_1[59]}
   );
   gpc1_1 gpc215 (
      {stage0_1[124]},
      {stage1_1[60]}
   );
   gpc1_1 gpc216 (
      {stage0_1[125]},
      {stage1_1[61]}
   );
   gpc1_1 gpc217 (
      {stage0_1[126]},
      {stage1_1[62]}
   );
   gpc1_1 gpc218 (
      {stage0_1[127]},
      {stage1_1[63]}
   );
   gpc1_1 gpc219 (
      {stage0_2[126]},
      {stage1_2[37]}
   );
   gpc1_1 gpc220 (
      {stage0_2[127]},
      {stage1_2[38]}
   );
   gpc1_1 gpc221 (
      {stage0_3[122]},
      {stage1_3[43]}
   );
   gpc1_1 gpc222 (
      {stage0_3[123]},
      {stage1_3[44]}
   );
   gpc1_1 gpc223 (
      {stage0_3[124]},
      {stage1_3[45]}
   );
   gpc1_1 gpc224 (
      {stage0_3[125]},
      {stage1_3[46]}
   );
   gpc1_1 gpc225 (
      {stage0_3[126]},
      {stage1_3[47]}
   );
   gpc1_1 gpc226 (
      {stage0_3[127]},
      {stage1_3[48]}
   );
   gpc1_1 gpc227 (
      {stage0_4[126]},
      {stage1_4[58]}
   );
   gpc1_1 gpc228 (
      {stage0_4[127]},
      {stage1_4[59]}
   );
   gpc1_1 gpc229 (
      {stage0_7[108]},
      {stage1_7[45]}
   );
   gpc1_1 gpc230 (
      {stage0_7[109]},
      {stage1_7[46]}
   );
   gpc1_1 gpc231 (
      {stage0_7[110]},
      {stage1_7[47]}
   );
   gpc1_1 gpc232 (
      {stage0_7[111]},
      {stage1_7[48]}
   );
   gpc1_1 gpc233 (
      {stage0_7[112]},
      {stage1_7[49]}
   );
   gpc1_1 gpc234 (
      {stage0_7[113]},
      {stage1_7[50]}
   );
   gpc1_1 gpc235 (
      {stage0_7[114]},
      {stage1_7[51]}
   );
   gpc1_1 gpc236 (
      {stage0_7[115]},
      {stage1_7[52]}
   );
   gpc1_1 gpc237 (
      {stage0_7[116]},
      {stage1_7[53]}
   );
   gpc1_1 gpc238 (
      {stage0_7[117]},
      {stage1_7[54]}
   );
   gpc1_1 gpc239 (
      {stage0_7[118]},
      {stage1_7[55]}
   );
   gpc1_1 gpc240 (
      {stage0_7[119]},
      {stage1_7[56]}
   );
   gpc1_1 gpc241 (
      {stage0_7[120]},
      {stage1_7[57]}
   );
   gpc1_1 gpc242 (
      {stage0_7[121]},
      {stage1_7[58]}
   );
   gpc1_1 gpc243 (
      {stage0_7[122]},
      {stage1_7[59]}
   );
   gpc1_1 gpc244 (
      {stage0_7[123]},
      {stage1_7[60]}
   );
   gpc1_1 gpc245 (
      {stage0_7[124]},
      {stage1_7[61]}
   );
   gpc1_1 gpc246 (
      {stage0_7[125]},
      {stage1_7[62]}
   );
   gpc1_1 gpc247 (
      {stage0_7[126]},
      {stage1_7[63]}
   );
   gpc1_1 gpc248 (
      {stage0_7[127]},
      {stage1_7[64]}
   );
   gpc1_1 gpc249 (
      {stage0_8[126]},
      {stage1_8[54]}
   );
   gpc1_1 gpc250 (
      {stage0_8[127]},
      {stage1_8[55]}
   );
   gpc1_1 gpc251 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc252 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc253 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc254 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc255 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc256 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc257 (
      {stage0_11[118]},
      {stage1_11[42]}
   );
   gpc1_1 gpc258 (
      {stage0_11[119]},
      {stage1_11[43]}
   );
   gpc1_1 gpc259 (
      {stage0_11[120]},
      {stage1_11[44]}
   );
   gpc1_1 gpc260 (
      {stage0_11[121]},
      {stage1_11[45]}
   );
   gpc1_1 gpc261 (
      {stage0_11[122]},
      {stage1_11[46]}
   );
   gpc1_1 gpc262 (
      {stage0_11[123]},
      {stage1_11[47]}
   );
   gpc1_1 gpc263 (
      {stage0_11[124]},
      {stage1_11[48]}
   );
   gpc1_1 gpc264 (
      {stage0_11[125]},
      {stage1_11[49]}
   );
   gpc1_1 gpc265 (
      {stage0_11[126]},
      {stage1_11[50]}
   );
   gpc1_1 gpc266 (
      {stage0_11[127]},
      {stage1_11[51]}
   );
   gpc1_1 gpc267 (
      {stage0_12[126]},
      {stage1_12[55]}
   );
   gpc1_1 gpc268 (
      {stage0_12[127]},
      {stage1_12[56]}
   );
   gpc1_1 gpc269 (
      {stage0_13[117]},
      {stage1_13[61]}
   );
   gpc1_1 gpc270 (
      {stage0_13[118]},
      {stage1_13[62]}
   );
   gpc1_1 gpc271 (
      {stage0_13[119]},
      {stage1_13[63]}
   );
   gpc1_1 gpc272 (
      {stage0_13[120]},
      {stage1_13[64]}
   );
   gpc1_1 gpc273 (
      {stage0_13[121]},
      {stage1_13[65]}
   );
   gpc1_1 gpc274 (
      {stage0_13[122]},
      {stage1_13[66]}
   );
   gpc1_1 gpc275 (
      {stage0_13[123]},
      {stage1_13[67]}
   );
   gpc1_1 gpc276 (
      {stage0_13[124]},
      {stage1_13[68]}
   );
   gpc1_1 gpc277 (
      {stage0_13[125]},
      {stage1_13[69]}
   );
   gpc1_1 gpc278 (
      {stage0_13[126]},
      {stage1_13[70]}
   );
   gpc1_1 gpc279 (
      {stage0_13[127]},
      {stage1_13[71]}
   );
   gpc1_1 gpc280 (
      {stage0_14[99]},
      {stage1_14[42]}
   );
   gpc1_1 gpc281 (
      {stage0_14[100]},
      {stage1_14[43]}
   );
   gpc1_1 gpc282 (
      {stage0_14[101]},
      {stage1_14[44]}
   );
   gpc1_1 gpc283 (
      {stage0_14[102]},
      {stage1_14[45]}
   );
   gpc1_1 gpc284 (
      {stage0_14[103]},
      {stage1_14[46]}
   );
   gpc1_1 gpc285 (
      {stage0_14[104]},
      {stage1_14[47]}
   );
   gpc1_1 gpc286 (
      {stage0_14[105]},
      {stage1_14[48]}
   );
   gpc1_1 gpc287 (
      {stage0_14[106]},
      {stage1_14[49]}
   );
   gpc1_1 gpc288 (
      {stage0_14[107]},
      {stage1_14[50]}
   );
   gpc1_1 gpc289 (
      {stage0_14[108]},
      {stage1_14[51]}
   );
   gpc1_1 gpc290 (
      {stage0_14[109]},
      {stage1_14[52]}
   );
   gpc1_1 gpc291 (
      {stage0_14[110]},
      {stage1_14[53]}
   );
   gpc1_1 gpc292 (
      {stage0_14[111]},
      {stage1_14[54]}
   );
   gpc1_1 gpc293 (
      {stage0_14[112]},
      {stage1_14[55]}
   );
   gpc1_1 gpc294 (
      {stage0_14[113]},
      {stage1_14[56]}
   );
   gpc1_1 gpc295 (
      {stage0_14[114]},
      {stage1_14[57]}
   );
   gpc1_1 gpc296 (
      {stage0_14[115]},
      {stage1_14[58]}
   );
   gpc1_1 gpc297 (
      {stage0_14[116]},
      {stage1_14[59]}
   );
   gpc1_1 gpc298 (
      {stage0_14[117]},
      {stage1_14[60]}
   );
   gpc1_1 gpc299 (
      {stage0_14[118]},
      {stage1_14[61]}
   );
   gpc1_1 gpc300 (
      {stage0_14[119]},
      {stage1_14[62]}
   );
   gpc1_1 gpc301 (
      {stage0_14[120]},
      {stage1_14[63]}
   );
   gpc1_1 gpc302 (
      {stage0_14[121]},
      {stage1_14[64]}
   );
   gpc1_1 gpc303 (
      {stage0_14[122]},
      {stage1_14[65]}
   );
   gpc1_1 gpc304 (
      {stage0_14[123]},
      {stage1_14[66]}
   );
   gpc1_1 gpc305 (
      {stage0_14[124]},
      {stage1_14[67]}
   );
   gpc1_1 gpc306 (
      {stage0_14[125]},
      {stage1_14[68]}
   );
   gpc1_1 gpc307 (
      {stage0_14[126]},
      {stage1_14[69]}
   );
   gpc1_1 gpc308 (
      {stage0_14[127]},
      {stage1_14[70]}
   );
   gpc1_1 gpc309 (
      {stage0_15[126]},
      {stage1_15[36]}
   );
   gpc1_1 gpc310 (
      {stage0_15[127]},
      {stage1_15[37]}
   );
   gpc1163_5 gpc311 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc312 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc313 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc314 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc315 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc316 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc317 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc319 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc320 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc321 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1406_5 gpc322 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[0]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc615_5 gpc323 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[26]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc615_5 gpc324 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[27]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc325 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage2_6[0],stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc326 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[7]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[4],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc327 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[8]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[5],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc328 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[9]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc329 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[10]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc330 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[11]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc606_5 gpc331 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[5],stage2_6[6],stage2_5[9],stage2_4[20]}
   );
   gpc606_5 gpc332 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[6],stage2_6[7],stage2_5[10],stage2_4[21]}
   );
   gpc606_5 gpc333 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[7],stage2_6[8],stage2_5[11],stage2_4[22]}
   );
   gpc606_5 gpc334 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[8],stage2_6[9],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc335 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[9],stage2_6[10],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc336 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[10],stage2_6[11],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc337 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[11],stage2_6[12],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc338 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[12],stage2_6[13],stage2_5[16],stage2_4[27]}
   );
   gpc207_4 gpc339 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[8],stage2_7[13],stage2_6[14],stage2_5[17]}
   );
   gpc606_5 gpc340 (
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[9],stage2_7[14],stage2_6[15],stage2_5[18]}
   );
   gpc606_5 gpc341 (
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[10],stage2_7[15],stage2_6[16],stage2_5[19]}
   );
   gpc615_5 gpc342 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[2],stage2_8[11],stage2_7[16]}
   );
   gpc615_5 gpc343 (
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[3],stage2_8[12],stage2_7[17]}
   );
   gpc615_5 gpc344 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[4],stage2_8[13],stage2_7[18]}
   );
   gpc615_5 gpc345 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[5],stage2_8[14],stage2_7[19]}
   );
   gpc615_5 gpc346 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[6],stage2_8[15],stage2_7[20]}
   );
   gpc615_5 gpc347 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[7],stage2_8[16],stage2_7[21]}
   );
   gpc615_5 gpc348 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[8],stage2_8[17],stage2_7[22]}
   );
   gpc615_5 gpc349 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[9],stage2_8[18],stage2_7[23]}
   );
   gpc615_5 gpc350 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[10],stage2_8[19],stage2_7[24]}
   );
   gpc606_5 gpc351 (
      {stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[9],stage2_10[9],stage2_9[11],stage2_8[20]}
   );
   gpc606_5 gpc352 (
      {stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[10],stage2_10[10],stage2_9[12],stage2_8[21]}
   );
   gpc606_5 gpc353 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[11],stage2_10[11],stage2_9[13],stage2_8[22]}
   );
   gpc606_5 gpc354 (
      {stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[12],stage2_10[12],stage2_9[14],stage2_8[23]}
   );
   gpc606_5 gpc355 (
      {stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[13],stage2_10[13],stage2_9[15],stage2_8[24]}
   );
   gpc606_5 gpc356 (
      {stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[14],stage2_10[14],stage2_9[16],stage2_8[25]}
   );
   gpc615_5 gpc357 (
      {stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_9[54]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[15],stage2_10[15],stage2_9[17],stage2_8[26]}
   );
   gpc615_5 gpc358 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_9[55]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[16],stage2_10[16],stage2_9[18],stage2_8[27]}
   );
   gpc606_5 gpc359 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[8],stage2_11[17],stage2_10[17]}
   );
   gpc615_5 gpc360 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[9],stage2_11[18]}
   );
   gpc615_5 gpc361 (
      {stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[10],stage2_11[19]}
   );
   gpc615_5 gpc362 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[11],stage2_11[20]}
   );
   gpc615_5 gpc363 (
      {stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[12],stage2_11[21]}
   );
   gpc615_5 gpc364 (
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_12[10]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[13],stage2_11[22]}
   );
   gpc615_5 gpc365 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_12[11]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[14],stage2_11[23]}
   );
   gpc615_5 gpc366 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[12]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[7],stage2_12[15],stage2_11[24]}
   );
   gpc615_5 gpc367 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[13]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[8],stage2_12[16],stage2_11[25]}
   );
   gpc207_4 gpc368 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19], stage1_12[20]},
      {stage1_14[0], stage1_14[1]},
      {stage2_15[8],stage2_14[9],stage2_13[9],stage2_12[17]}
   );
   gpc606_5 gpc369 (
      {stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25], stage1_12[26]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[0],stage2_15[9],stage2_14[10],stage2_13[10],stage2_12[18]}
   );
   gpc606_5 gpc370 (
      {stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[1],stage2_15[10],stage2_14[11],stage2_13[11],stage2_12[19]}
   );
   gpc606_5 gpc371 (
      {stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[2],stage2_15[11],stage2_14[12],stage2_13[12],stage2_12[20]}
   );
   gpc606_5 gpc372 (
      {stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[3],stage2_15[12],stage2_14[13],stage2_13[13],stage2_12[21]}
   );
   gpc606_5 gpc373 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[4],stage2_15[13],stage2_14[14],stage2_13[14],stage2_12[22]}
   );
   gpc606_5 gpc374 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[15],stage2_13[15]}
   );
   gpc606_5 gpc375 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[16],stage2_13[16]}
   );
   gpc606_5 gpc376 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[17],stage2_13[17]}
   );
   gpc606_5 gpc377 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[18],stage2_13[18]}
   );
   gpc606_5 gpc378 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[19]}
   );
   gpc606_5 gpc379 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[20]}
   );
   gpc606_5 gpc380 (
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[21]}
   );
   gpc615_5 gpc381 (
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_15[24]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[22]}
   );
   gpc615_5 gpc382 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[25]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[23]}
   );
   gpc615_5 gpc383 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30]},
      {stage1_16[30]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23]}
   );
   gpc615_5 gpc384 (
      {stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[31]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24]}
   );
   gpc1_1 gpc385 (
      {stage1_0[42]},
      {stage2_0[11]}
   );
   gpc1_1 gpc386 (
      {stage1_0[43]},
      {stage2_0[12]}
   );
   gpc1_1 gpc387 (
      {stage1_0[44]},
      {stage2_0[13]}
   );
   gpc1_1 gpc388 (
      {stage1_0[45]},
      {stage2_0[14]}
   );
   gpc1_1 gpc389 (
      {stage1_2[34]},
      {stage2_2[15]}
   );
   gpc1_1 gpc390 (
      {stage1_2[35]},
      {stage2_2[16]}
   );
   gpc1_1 gpc391 (
      {stage1_2[36]},
      {stage2_2[17]}
   );
   gpc1_1 gpc392 (
      {stage1_2[37]},
      {stage2_2[18]}
   );
   gpc1_1 gpc393 (
      {stage1_2[38]},
      {stage2_2[19]}
   );
   gpc1_1 gpc394 (
      {stage1_5[49]},
      {stage2_5[20]}
   );
   gpc1_1 gpc395 (
      {stage1_5[50]},
      {stage2_5[21]}
   );
   gpc1_1 gpc396 (
      {stage1_5[51]},
      {stage2_5[22]}
   );
   gpc1_1 gpc397 (
      {stage1_5[52]},
      {stage2_5[23]}
   );
   gpc1_1 gpc398 (
      {stage1_5[53]},
      {stage2_5[24]}
   );
   gpc1_1 gpc399 (
      {stage1_5[54]},
      {stage2_5[25]}
   );
   gpc1_1 gpc400 (
      {stage1_5[55]},
      {stage2_5[26]}
   );
   gpc1_1 gpc401 (
      {stage1_5[56]},
      {stage2_5[27]}
   );
   gpc1_1 gpc402 (
      {stage1_7[59]},
      {stage2_7[25]}
   );
   gpc1_1 gpc403 (
      {stage1_7[60]},
      {stage2_7[26]}
   );
   gpc1_1 gpc404 (
      {stage1_7[61]},
      {stage2_7[27]}
   );
   gpc1_1 gpc405 (
      {stage1_7[62]},
      {stage2_7[28]}
   );
   gpc1_1 gpc406 (
      {stage1_7[63]},
      {stage2_7[29]}
   );
   gpc1_1 gpc407 (
      {stage1_7[64]},
      {stage2_7[30]}
   );
   gpc1_1 gpc408 (
      {stage1_8[55]},
      {stage2_8[28]}
   );
   gpc1_1 gpc409 (
      {stage1_9[56]},
      {stage2_9[19]}
   );
   gpc1_1 gpc410 (
      {stage1_9[57]},
      {stage2_9[20]}
   );
   gpc1_1 gpc411 (
      {stage1_11[40]},
      {stage2_11[26]}
   );
   gpc1_1 gpc412 (
      {stage1_11[41]},
      {stage2_11[27]}
   );
   gpc1_1 gpc413 (
      {stage1_11[42]},
      {stage2_11[28]}
   );
   gpc1_1 gpc414 (
      {stage1_11[43]},
      {stage2_11[29]}
   );
   gpc1_1 gpc415 (
      {stage1_11[44]},
      {stage2_11[30]}
   );
   gpc1_1 gpc416 (
      {stage1_11[45]},
      {stage2_11[31]}
   );
   gpc1_1 gpc417 (
      {stage1_11[46]},
      {stage2_11[32]}
   );
   gpc1_1 gpc418 (
      {stage1_11[47]},
      {stage2_11[33]}
   );
   gpc1_1 gpc419 (
      {stage1_11[48]},
      {stage2_11[34]}
   );
   gpc1_1 gpc420 (
      {stage1_11[49]},
      {stage2_11[35]}
   );
   gpc1_1 gpc421 (
      {stage1_11[50]},
      {stage2_11[36]}
   );
   gpc1_1 gpc422 (
      {stage1_11[51]},
      {stage2_11[37]}
   );
   gpc1_1 gpc423 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc424 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc425 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc426 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc427 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc428 (
      {stage1_12[56]},
      {stage2_12[28]}
   );
   gpc1_1 gpc429 (
      {stage1_14[60]},
      {stage2_14[24]}
   );
   gpc1_1 gpc430 (
      {stage1_14[61]},
      {stage2_14[25]}
   );
   gpc1_1 gpc431 (
      {stage1_14[62]},
      {stage2_14[26]}
   );
   gpc1_1 gpc432 (
      {stage1_14[63]},
      {stage2_14[27]}
   );
   gpc1_1 gpc433 (
      {stage1_14[64]},
      {stage2_14[28]}
   );
   gpc1_1 gpc434 (
      {stage1_14[65]},
      {stage2_14[29]}
   );
   gpc1_1 gpc435 (
      {stage1_14[66]},
      {stage2_14[30]}
   );
   gpc1_1 gpc436 (
      {stage1_14[67]},
      {stage2_14[31]}
   );
   gpc1_1 gpc437 (
      {stage1_14[68]},
      {stage2_14[32]}
   );
   gpc1_1 gpc438 (
      {stage1_14[69]},
      {stage2_14[33]}
   );
   gpc1_1 gpc439 (
      {stage1_14[70]},
      {stage2_14[34]}
   );
   gpc1_1 gpc440 (
      {stage1_15[36]},
      {stage2_15[25]}
   );
   gpc1_1 gpc441 (
      {stage1_15[37]},
      {stage2_15[26]}
   );
   gpc1_1 gpc442 (
      {stage1_16[32]},
      {stage2_16[16]}
   );
   gpc1_1 gpc443 (
      {stage1_16[33]},
      {stage2_16[17]}
   );
   gpc1_1 gpc444 (
      {stage1_16[34]},
      {stage2_16[18]}
   );
   gpc1_1 gpc445 (
      {stage1_16[35]},
      {stage2_16[19]}
   );
   gpc1_1 gpc446 (
      {stage1_17[12]},
      {stage2_17[11]}
   );
   gpc1_1 gpc447 (
      {stage1_17[13]},
      {stage2_17[12]}
   );
   gpc1_1 gpc448 (
      {stage1_17[14]},
      {stage2_17[13]}
   );
   gpc1_1 gpc449 (
      {stage1_17[15]},
      {stage2_17[14]}
   );
   gpc1_1 gpc450 (
      {stage1_17[16]},
      {stage2_17[15]}
   );
   gpc1_1 gpc451 (
      {stage1_17[17]},
      {stage2_17[16]}
   );
   gpc1_1 gpc452 (
      {stage1_17[18]},
      {stage2_17[17]}
   );
   gpc1_1 gpc453 (
      {stage1_17[19]},
      {stage2_17[18]}
   );
   gpc1_1 gpc454 (
      {stage1_17[20]},
      {stage2_17[19]}
   );
   gpc606_5 gpc455 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc456 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc615_5 gpc457 (
      {stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc458 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc1163_5 gpc459 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[4]}
   );
   gpc606_5 gpc460 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[4],stage3_5[5]}
   );
   gpc615_5 gpc461 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_6[2]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc615_5 gpc462 (
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_6[3]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc615_5 gpc463 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_6[4]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc615_5 gpc464 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27]},
      {stage2_6[5]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[4],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc465 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[5],stage3_7[7],stage3_6[9]}
   );
   gpc615_5 gpc466 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_7[30]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[6],stage3_7[8],stage3_6[10]}
   );
   gpc606_5 gpc467 (
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[2],stage3_9[7],stage3_8[7]}
   );
   gpc606_5 gpc468 (
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[3],stage3_9[8],stage3_8[8]}
   );
   gpc1163_5 gpc469 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[2],stage3_10[4],stage3_9[9]}
   );
   gpc606_5 gpc470 (
      {stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage3_13[1],stage3_12[3],stage3_11[3],stage3_10[5],stage3_9[10]}
   );
   gpc606_5 gpc471 (
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage3_13[2],stage3_12[4],stage3_11[4],stage3_10[6],stage3_9[11]}
   );
   gpc606_5 gpc472 (
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage3_13[3],stage3_12[5],stage3_11[5],stage3_10[7],stage3_9[12]}
   );
   gpc615_5 gpc473 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_12[1]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[6],stage3_11[6]}
   );
   gpc615_5 gpc474 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[7],stage3_11[7]}
   );
   gpc606_5 gpc475 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[8]}
   );
   gpc606_5 gpc476 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[9]}
   );
   gpc606_5 gpc477 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[10]}
   );
   gpc606_5 gpc478 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[11]}
   );
   gpc606_5 gpc479 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[6],stage3_14[6],stage3_13[10]}
   );
   gpc1163_5 gpc480 (
      {stage2_14[24], stage2_14[25], stage2_14[26]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc481 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[1]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[0],stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[8]}
   );
   gpc615_5 gpc482 (
      {stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_16[2]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[1],stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[9]}
   );
   gpc615_5 gpc483 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26]},
      {stage2_16[3]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[2],stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[10]}
   );
   gpc606_5 gpc484 (
      {stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[3],stage3_18[4],stage3_17[5],stage3_16[9]}
   );
   gpc1_1 gpc485 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc486 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc487 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc488 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc489 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc490 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc491 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc492 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc493 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc494 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc495 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc496 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc497 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc498 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc499 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc500 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc501 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc502 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc503 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc504 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc505 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc506 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc507 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc508 (
      {stage2_2[10]},
      {stage3_2[3]}
   );
   gpc1_1 gpc509 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc510 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc511 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc512 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc513 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc514 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc515 (
      {stage2_2[17]},
      {stage3_2[10]}
   );
   gpc1_1 gpc516 (
      {stage2_2[18]},
      {stage3_2[11]}
   );
   gpc1_1 gpc517 (
      {stage2_2[19]},
      {stage3_2[12]}
   );
   gpc1_1 gpc518 (
      {stage2_3[14]},
      {stage3_3[5]}
   );
   gpc1_1 gpc519 (
      {stage2_3[15]},
      {stage3_3[6]}
   );
   gpc1_1 gpc520 (
      {stage2_3[16]},
      {stage3_3[7]}
   );
   gpc1_1 gpc521 (
      {stage2_3[17]},
      {stage3_3[8]}
   );
   gpc1_1 gpc522 (
      {stage2_3[18]},
      {stage3_3[9]}
   );
   gpc1_1 gpc523 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc524 (
      {stage2_4[24]},
      {stage3_4[5]}
   );
   gpc1_1 gpc525 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc526 (
      {stage2_4[26]},
      {stage3_4[7]}
   );
   gpc1_1 gpc527 (
      {stage2_4[27]},
      {stage3_4[8]}
   );
   gpc1_1 gpc528 (
      {stage2_8[24]},
      {stage3_8[9]}
   );
   gpc1_1 gpc529 (
      {stage2_8[25]},
      {stage3_8[10]}
   );
   gpc1_1 gpc530 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc531 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc532 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc533 (
      {stage2_11[29]},
      {stage3_11[8]}
   );
   gpc1_1 gpc534 (
      {stage2_11[30]},
      {stage3_11[9]}
   );
   gpc1_1 gpc535 (
      {stage2_11[31]},
      {stage3_11[10]}
   );
   gpc1_1 gpc536 (
      {stage2_11[32]},
      {stage3_11[11]}
   );
   gpc1_1 gpc537 (
      {stage2_11[33]},
      {stage3_11[12]}
   );
   gpc1_1 gpc538 (
      {stage2_11[34]},
      {stage3_11[13]}
   );
   gpc1_1 gpc539 (
      {stage2_11[35]},
      {stage3_11[14]}
   );
   gpc1_1 gpc540 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc541 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc542 (
      {stage2_12[27]},
      {stage3_12[12]}
   );
   gpc1_1 gpc543 (
      {stage2_12[28]},
      {stage3_12[13]}
   );
   gpc1_1 gpc544 (
      {stage2_13[18]},
      {stage3_13[11]}
   );
   gpc1_1 gpc545 (
      {stage2_14[27]},
      {stage3_14[8]}
   );
   gpc1_1 gpc546 (
      {stage2_14[28]},
      {stage3_14[9]}
   );
   gpc1_1 gpc547 (
      {stage2_14[29]},
      {stage3_14[10]}
   );
   gpc1_1 gpc548 (
      {stage2_14[30]},
      {stage3_14[11]}
   );
   gpc1_1 gpc549 (
      {stage2_14[31]},
      {stage3_14[12]}
   );
   gpc1_1 gpc550 (
      {stage2_14[32]},
      {stage3_14[13]}
   );
   gpc1_1 gpc551 (
      {stage2_14[33]},
      {stage3_14[14]}
   );
   gpc1_1 gpc552 (
      {stage2_14[34]},
      {stage3_14[15]}
   );
   gpc1_1 gpc553 (
      {stage2_16[10]},
      {stage3_16[10]}
   );
   gpc1_1 gpc554 (
      {stage2_16[11]},
      {stage3_16[11]}
   );
   gpc1_1 gpc555 (
      {stage2_16[12]},
      {stage3_16[12]}
   );
   gpc1_1 gpc556 (
      {stage2_16[13]},
      {stage3_16[13]}
   );
   gpc1_1 gpc557 (
      {stage2_16[14]},
      {stage3_16[14]}
   );
   gpc1_1 gpc558 (
      {stage2_16[15]},
      {stage3_16[15]}
   );
   gpc1_1 gpc559 (
      {stage2_16[16]},
      {stage3_16[16]}
   );
   gpc1_1 gpc560 (
      {stage2_16[17]},
      {stage3_16[17]}
   );
   gpc1_1 gpc561 (
      {stage2_16[18]},
      {stage3_16[18]}
   );
   gpc1_1 gpc562 (
      {stage2_16[19]},
      {stage3_16[19]}
   );
   gpc1_1 gpc563 (
      {stage2_17[19]},
      {stage3_17[6]}
   );
   gpc1_1 gpc564 (
      {stage2_18[6]},
      {stage3_18[5]}
   );
   gpc1_1 gpc565 (
      {stage2_19[0]},
      {stage3_19[4]}
   );
   gpc1_1 gpc566 (
      {stage2_19[1]},
      {stage3_19[5]}
   );
   gpc606_5 gpc567 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc568 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10]},
      {stage3_1[0]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1163_5 gpc569 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc570 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc615_5 gpc571 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc572 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[2],stage4_7[3],stage4_6[3]}
   );
   gpc606_5 gpc573 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[2],stage4_9[3]}
   );
   gpc615_5 gpc574 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[3],stage4_9[4]}
   );
   gpc606_5 gpc575 (
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[4]}
   );
   gpc615_5 gpc576 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16]},
      {stage3_12[6]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc577 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc578 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[5]}
   );
   gpc615_5 gpc579 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[4]}
   );
   gpc615_5 gpc580 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[7]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[5]}
   );
   gpc606_5 gpc581 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4]}
   );
   gpc606_5 gpc582 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[3],stage4_17[4]}
   );
   gpc1_1 gpc583 (
      {stage3_0[11]},
      {stage4_0[2]}
   );
   gpc1_1 gpc584 (
      {stage3_0[12]},
      {stage4_0[3]}
   );
   gpc1_1 gpc585 (
      {stage3_0[13]},
      {stage4_0[4]}
   );
   gpc1_1 gpc586 (
      {stage3_0[14]},
      {stage4_0[5]}
   );
   gpc1_1 gpc587 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc588 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc589 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc590 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc591 (
      {stage3_1[5]},
      {stage4_1[6]}
   );
   gpc1_1 gpc592 (
      {stage3_1[6]},
      {stage4_1[7]}
   );
   gpc1_1 gpc593 (
      {stage3_1[7]},
      {stage4_1[8]}
   );
   gpc1_1 gpc594 (
      {stage3_1[8]},
      {stage4_1[9]}
   );
   gpc1_1 gpc595 (
      {stage3_2[12]},
      {stage4_2[2]}
   );
   gpc1_1 gpc596 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc597 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc598 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc599 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc600 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc601 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc602 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc603 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc604 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc605 (
      {stage3_4[7]},
      {stage4_4[4]}
   );
   gpc1_1 gpc606 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc607 (
      {stage3_5[7]},
      {stage4_5[2]}
   );
   gpc1_1 gpc608 (
      {stage3_5[8]},
      {stage4_5[3]}
   );
   gpc1_1 gpc609 (
      {stage3_5[9]},
      {stage4_5[4]}
   );
   gpc1_1 gpc610 (
      {stage3_7[8]},
      {stage4_7[4]}
   );
   gpc1_1 gpc611 (
      {stage3_8[12]},
      {stage4_8[3]}
   );
   gpc1_1 gpc612 (
      {stage3_8[13]},
      {stage4_8[4]}
   );
   gpc1_1 gpc613 (
      {stage3_9[11]},
      {stage4_9[5]}
   );
   gpc1_1 gpc614 (
      {stage3_9[12]},
      {stage4_9[6]}
   );
   gpc1_1 gpc615 (
      {stage3_10[7]},
      {stage4_10[5]}
   );
   gpc1_1 gpc616 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc617 (
      {stage3_15[8]},
      {stage4_15[5]}
   );
   gpc1_1 gpc618 (
      {stage3_15[9]},
      {stage4_15[6]}
   );
   gpc1_1 gpc619 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc620 (
      {stage3_16[18]},
      {stage4_16[5]}
   );
   gpc1_1 gpc621 (
      {stage3_16[19]},
      {stage4_16[6]}
   );
   gpc1_1 gpc622 (
      {stage3_17[6]},
      {stage4_17[5]}
   );
   gpc1_1 gpc623 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc2135_5 gpc624 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1415_5 gpc625 (
      {stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6], stage4_1[7]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1415_5 gpc626 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc627 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[1]}
   );
   gpc606_5 gpc628 (
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc135_4 gpc629 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1]}
   );
   gpc1343_5 gpc630 (
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0], stage4_19[1], 1'b0, 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1_1 gpc631 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc632 (
      {stage4_1[8]},
      {stage5_1[2]}
   );
   gpc1_1 gpc633 (
      {stage4_1[9]},
      {stage5_1[3]}
   );
   gpc1_1 gpc634 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc635 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc636 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc637 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc638 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc639 (
      {stage4_3[10]},
      {stage5_3[6]}
   );
   gpc1_1 gpc640 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc641 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc642 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc643 (
      {stage4_5[4]},
      {stage5_5[5]}
   );
   gpc1_1 gpc644 (
      {stage4_7[1]},
      {stage5_7[1]}
   );
   gpc1_1 gpc645 (
      {stage4_7[2]},
      {stage5_7[2]}
   );
   gpc1_1 gpc646 (
      {stage4_7[3]},
      {stage5_7[3]}
   );
   gpc1_1 gpc647 (
      {stage4_7[4]},
      {stage5_7[4]}
   );
   gpc1_1 gpc648 (
      {stage4_9[1]},
      {stage5_9[1]}
   );
   gpc1_1 gpc649 (
      {stage4_9[2]},
      {stage5_9[2]}
   );
   gpc1_1 gpc650 (
      {stage4_9[3]},
      {stage5_9[3]}
   );
   gpc1_1 gpc651 (
      {stage4_9[4]},
      {stage5_9[4]}
   );
   gpc1_1 gpc652 (
      {stage4_9[5]},
      {stage5_9[5]}
   );
   gpc1_1 gpc653 (
      {stage4_9[6]},
      {stage5_9[6]}
   );
   gpc1_1 gpc654 (
      {stage4_11[0]},
      {stage5_11[1]}
   );
   gpc1_1 gpc655 (
      {stage4_11[1]},
      {stage5_11[2]}
   );
   gpc1_1 gpc656 (
      {stage4_11[2]},
      {stage5_11[3]}
   );
   gpc1_1 gpc657 (
      {stage4_11[3]},
      {stage5_11[4]}
   );
   gpc1_1 gpc658 (
      {stage4_13[0]},
      {stage5_13[1]}
   );
   gpc1_1 gpc659 (
      {stage4_13[1]},
      {stage5_13[2]}
   );
   gpc1_1 gpc660 (
      {stage4_13[2]},
      {stage5_13[3]}
   );
   gpc1_1 gpc661 (
      {stage4_13[3]},
      {stage5_13[4]}
   );
   gpc1_1 gpc662 (
      {stage4_13[4]},
      {stage5_13[5]}
   );
   gpc1_1 gpc663 (
      {stage4_13[5]},
      {stage5_13[6]}
   );
   gpc1_1 gpc664 (
      {stage4_15[5]},
      {stage5_15[2]}
   );
   gpc1_1 gpc665 (
      {stage4_15[6]},
      {stage5_15[3]}
   );
   gpc1_1 gpc666 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc667 (
      {stage4_16[3]},
      {stage5_16[2]}
   );
   gpc1_1 gpc668 (
      {stage4_16[4]},
      {stage5_16[3]}
   );
   gpc1_1 gpc669 (
      {stage4_16[5]},
      {stage5_16[4]}
   );
   gpc1_1 gpc670 (
      {stage4_16[6]},
      {stage5_16[5]}
   );
   gpc1_1 gpc671 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc672 (
      {stage4_17[2]},
      {stage5_17[2]}
   );
   gpc1_1 gpc673 (
      {stage4_17[3]},
      {stage5_17[3]}
   );
   gpc1_1 gpc674 (
      {stage4_17[4]},
      {stage5_17[4]}
   );
   gpc1_1 gpc675 (
      {stage4_17[5]},
      {stage5_17[5]}
   );
   gpc1_1 gpc676 (
      {stage4_18[3]},
      {stage5_18[2]}
   );
   gpc2223_5 gpc677 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1]},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc678 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc679 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1]}
   );
   gpc615_5 gpc680 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1]}
   );
   gpc615_5 gpc681 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc682 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2], 1'b0},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc1_1 gpc683 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc684 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc685 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc686 (
      {stage5_2[2]},
      {stage6_2[1]}
   );
   gpc1_1 gpc687 (
      {stage5_6[0]},
      {stage6_6[1]}
   );
   gpc1_1 gpc688 (
      {stage5_8[1]},
      {stage6_8[1]}
   );
   gpc1_1 gpc689 (
      {stage5_9[6]},
      {stage6_9[1]}
   );
   gpc1_1 gpc690 (
      {stage5_10[0]},
      {stage6_10[1]}
   );
   gpc1_1 gpc691 (
      {stage5_12[1]},
      {stage6_12[1]}
   );
   gpc1_1 gpc692 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc693 (
      {stage5_14[0]},
      {stage6_14[1]}
   );
   gpc1_1 gpc694 (
      {stage5_20[0]},
      {stage6_20[1]}
   );
   gpc1_1 gpc695 (
      {stage5_21[0]},
      {stage6_21[0]}
   );
   gpc1_1 gpc696 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor_CLA128_16 compressor_CLA128_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2c1b69f3077c2d62b60f822246a572b57ac397ab09bec2afc5d5c507fd9fa8f8243affbc63cb43daa51dce07006d06bc6c795697d4b6e1f1d7489516be973bdd80924e80faeeb6673378a87985382df4502f95bac5969a4fc0637ab9136add3e0b79b73e0392087de6b4a9f51b84c448764c9eeee3eddda8417014204a15de8075bd3be38ff91fba54275b915c6146221225e3d5015231565fcc5053432749b982eed91903a772793dd62b9750bdd98cf9080f1a814fd1c835e9324512a7accbb3f9dea7ecae0ba3f96ce2567972e39bcbe4827ea4026dda717ef809690c84cc1e02bb09a1e130fc9da725c0a237de57d5465ee8370c2339efd9bdee8b1e2661;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdd3ea6e85c5532dbee43284f8e024786da78f9f879ce517c4805d2759e76bda68d53c313265fc6b4f509b54c63eaef99b3211229b867d1fce13e5bc2e2fbe561a9e3621f337b7e8aea427d6bdd1537124867cd9c001ae1a8d9bfe3222673929cb57448191ac7b683f5f9ed748c29087c374112f1dca93c39be5a037cb392121782b68fed5810698516490d385c23f720be6d441348803f7431e3fac1efed3705cc57ab51fe19ed8e292c06f3888a426ef38aed66f66b20ee38c342f7fcf8f44669f757939798c80ebf63e9cb33535593e44355f1c33aa3a3e801ed975ea30d9f645357ec22ad9fb0e594daa7139072d177238e10c4d99f69ef1d9635932851f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf5af18ddc26b1ab04f2d0200f0b1191f5045bddf234750d017e963f7fa5abf26697d8b3d2443b6e8991b628a4e05614576bd8e14e99602bccd9ba7085433f11afb2c687a05306f1cfa0134fd00411ece0aba77f69f2333b3818369e3ffc60cb8ddc69dad0ce13d63eed9bcdcb69a11f5834ae221468cb38fa375459c86ec587c95b623011f0d5a98d231dfdf8de6f0053c6e18b44d6c4fe340ab175a2172cddbfc0a5ecde86860071328fa2243d7f67a856c490b43ddc3e99737c2c2636bdffb4ffa9dc2c74d6659b9fc295526bd0595ec40d07f9f4cd1a5ae0d68e9a519f51966522cb4881af8a4c7fbc894efc6cac6d91fd86d7dc479a7f7a0021ef95f2ff1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha8537aa74e78dd3fffd67f5b1b0467d756060dcc379767aec59d9188a97ea66684df38e20dc4c0f9a7e99fb088938405292914c66d9ac3137a9c424feb2499fffad5800e6fac6abeece6e5408b1d14a3ccf592bb49e3dc53a27612f94840643219577c549358c0ce232bcba9fb26aa8d74015413640f77e15408167a7256314af33152ede37f06abb2bb1d71ebe30444d3589e8458ad8cd87fa11b3f6a99532b43e30be5cc881be33e03ebf23be7c4d82d515a0aa9dd421134512fd39baa5c64510bc7ab24269c9f309e93e80c3617e30b425edeb4990a3d9973acdb9bd3abaeed18b67df819b4e9606948c6c3e436f24b6555574934b59577f2210c5e2c76f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hed71daa6016fe6ef477a35a585ecc5e3de3db659bfd0ec619dceae748fc4393b6dda085eda9d7fda377e8599696d82afd508d1b92a4369fd795e2c219f081bc5be9be94cf1ac5fe6dd68ed96c9df153ab48c50ba9824a093b6d213a5b3a93028b28d9c11470ef1fe15279b7693548ee4c7f46d6d1426e8082ab5c2d3ef2c2fb1a5de8cf9fd49b6af314e7e4e117ab6b93fbc9ab8b5354343042d2fa29ad32e3f6a924ae9914f0c6e833609999abb1d39aa43bc6e8686be76711a9975b30b6668865960c0cb542c962be3e45b43b5fcb1d2ece28c61b5b7246c52caee74d221a0c2182459de6faa0fdd1d8bbb889dd699090f58bacb8dbf9f9ec5352a3e253623;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1faf5cf139ff9f723aa75955c94a3dab73f0a1a5249ff125701bf23b96178fe5a31e908df41df51ae93674610c12183089cb8b78949ea92feea7b0a1bc6f1415a4c652c7f6565d48405911d0ba0bdec5ad2d3fb2b47718e7e29977b691040c310345e9ca7591671049edb08ad8b0cc94af748890c73f8fcd430d79b000f207953a4ca3bd001726e4df2a193f1306b8a60e7718daedf340291a73dfc7aea80f3552ca2a3ea4d31f48036434f0896af11e1f96a151cb0b61edd5e8db23888b1bc46819c3ad734e98f6854bb56d66deac0450b81ae49832f6ad7bf36d2bf77e29bd85c359f11449d6d6ce60a9e83f6e509a61453307ebe8d80ff3727c10e00832c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdeec85a4ee6aecff9576590af67ab23fd3f66dc9840f88fd07cc283054f30ff6521c781af69afc0c7fc2b6191716902400d585f3e0b4c208331f1aac19e2ec737c1d29fbd847f94173c595fe73da4c8fab861930950e67ac0a60a25b39a1e6da0e4fda6a1401f3181034bffaf9e3d84c3c71895a8bcc3980f1c1b960fcbd5bd55de3c3595f4bf95fa5a528055692a13acb502f21c75c2fe46ae7dc64c765d3d4f3fb248c8c6169af52b849c653bdacafb1f62edf7926d706a17bfc6c85873c05eae0ddf267f5b1b12629483d823cd94a084370adcac7465040b1bf221c9e1877f36bb3c8cc43b4592a6b1e3b0dfa5f4a5870d0cd07616358e688755f1fe4f800;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5685b2ff449e6a1fe5c45760629baff0b695b7726490e3e65536137be185f1e2467cf0d451d23f529b0e66848455e66466dd3e8c13fdfa1dd88cd46fa0ec2165dd0d4c0882bb8593fd72171c8718cd04b043e9f29bd2f2eadae6f82cf614aee1c5914b2c2bed69f0cd908277d91e99e445323dec72bb9941d8d281cded1e3dd836a3b0c2f412ff21bebde7fbcd6d0b0f5caad8826a49a61b815a517ee485024c7e056b656f346b5cbb2dfa078d980565e45f2b41ed8c32bef4ec8720e33b4c53229c21d266b29d0d247168e38fa4542b906a4a22430e4e7cb732b5906b6561e1c21f2079861b142965768da1991469e9c7885b9dcd2528eabe08eb8a32e49cf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha688e7da150f88b747bf995f1cb72f00bfbf27b001f27018efd918c358b243a5a597fcb1198075094e90fdae9b288b515ce1db9d28200cff16f7ad2c145ee8a661493db7e5cc5f407b93581d160e89b24fadbea76e403072377afb5c49c059e82653a84a13e9685dfa51ea8c58d698b079ca83465a45a8893342edcd07680f0fbe8ab608184788eb507bb716d85be5d0ad21fc7530308e3b26d52e8e0baba1048056b1a0ac366998e07ac427b69d4c7bea4383d8f235052ee565e2f2b5bb52f94e7d2fcb85d2920456e1ed0572823c3988203b437bc734098ce9bae45067b7875fe6cc32d77f18c292c4c99e2ee701d110bd258a33e6937af678a1e27bd23b96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5300e3f7bd9169c4aaea2ec160ca4c7145214a03226cb950dfa6b03e2196fc6adae3b94c7253e1d06ec3ef1e48ffde946a7cf758a1fe17c518fffaff72dbcfcfaf7916d62bf3605e9e1859d63c930665aff3a6baf192604d8094dc0c1b1b3309b38e64d9607bd9e47df706bc6eaa4b6904d00d0357bafdeabf4d3429364d14d1c087d32425e5c54b11202bad9ed20190d3892b2d0a92b13466c9e21e401abd98351a3978c669ebeb68f642b54d134bb23987cc47694936f6358e8ee85bda151f17aa0f31a21963d695f0503486b6b266652b6a0b6d5173e7f9326f9aea4a59387a004e70ae7d47843174a4f4bc449899fca3503eeb140d627991c4d29240b956;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hef5c2362ac8ce6f9e1840f65be7b1e79bd787caf2583a5cd6d1359a6ccc95499d2273f56d6aa86f18169cd99f4ea21dfa83cc3095f4c986ae2039fb0bea708a18fb565678b9b71d8089aaae3c164ccdd3380f31a7fab270ecd90661293c29f41667c494f72b946e65095afdd9685dcf92fc1a23d5d854d2db4fd987ed10334d3a387da4bd00e635776998e32da3ecc4370d2729c77c9d28666aec75af8ee56b0132d05bed58105d9d3052024b714633e16bab2592efda5ab81833c64936b695384359ad7e16dad11c6152a5983f7292d84a545fc3d272874f4d9453953a5057dc0a5b58d732b4a74103f71b975a69f3d09bd34725718252882583083d6e66862;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h361e80c1415bd83f53f044beaff511dfe38a529cde87e012a2671303c80dc067b80ac646f567722c28ec4f843fbf8d48e17a09cb20508b5c4249cd3e2a252c1b6fb920fe1b9a7a6ef849f57068c0b625aacec5901e1f42eca85f3fa946878614afeda7309e6fb5ec19c065cb5859e792f584671ed0ce2ac3d5deccabe13eb423414f92738c59106b7791686078d13b9cf9ace4621c877d76d51dbc16ffb084cdba8df25b73ba212874583fdc858c18e7baec52bdc01266c3e3c1204b709c5c57a56014d2184963753b2e1ed41b6e3d6738af752aa7c5d575c22c3a0ec499e43e11587959b6f98f3aef1a0d3f76c99fb41a72bf271dbd19cd1ed4b8686aa2ae70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3aa3ee85c165c2739af55b48ed1f8b9a1958bda0e442e8f9021e6d08e9465ba8c1373256241e125bfdc01d559acd21cd30c13f11f603fbf3501f4f83812dd9c64a46aaa3082ba9fa74f507c041fd5ce75b15c48d0632962066414b121034a84940d1d4c5b0ab74d5183e76ef5c548888f20fc06c6bd46feb587eeda72c895b557081f480b8d0149085451fc8bba03c95c897222c6ccf5b10029bf1a606c6a181b055428d140713225fede2535f7f683b913ed8a2eef933463b74aed923c13ed653ce0cde45851e7086552ec3cc68ce980d86f1a2d9b83cdadf69bcbfb6b51d6b91dbc31ef8ef51bcbb1b00d837ede15150acdb04a3dcf15d5a53f3d542c13e3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h38cfb1bd1a3f4654e9d042efa14d81e82d7857a2a1520acb8a6f5779903559984368878ae237ed473fcc6a4adb02136981ea70520ec96ef637a526085fea3a63f7a6bf51bf8d7d515b46b10d75da8c4478bb2bc3708db1b73634b5a98edb8b5160bd8ced1d55640e59ab5d982367907be920c68522ceb9a12dec86dcf3e33e7fbc24a09da5895bb97cdd31ec8259ebcc8ee4cecfc1b9e6b1f2959e5bda113bf0bbea7f23af03d8747757536990e9fd390e59afab61da87f3fa7ad64b753a59669bbdb0bafce3cf031248f91d0f9fd9c87fd7ce95e932aa39fe75056b12fe14902087ae2abb0cb27560794b213246106a40ea38c2da3023b9cacac4697837f309;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9436844ae3cadbc913aae1d7ab96a7d610757de90be461c70e1ea307fec891f4545bfa3e676526e4dacfe215e355c477cf8da2fe1f80a9cc02c2795c3ed038bd17cc7b37861fca01f775aecb44ff996751a5383164afc6b5ca979a411b09429a52bc87d78e15a2bd9bafd2e2f45f8355763c0df290dc392250dff05699fb6d0349a812e809fec0945bb2c34f4f76bd351552f5fda0e78097fe9206da931cf2203bb3fa0a3e495480b55e420b1f7a7f2fa7e3c57a626100fd283f991c68b12b208260e1ed35707d177980902f1cc1eaf1962cac7caae5cd325dfd7ec7ae1b5e16822891f3b1b4b4c4efffff6ab0d888d981265221a96c5ce554f52882b782b18b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h252b44376f89c5b0c5f159de010e2e36a79f37c15eccb118d5e68d9b73b838392bc2c8ec2e27a2a428bc967dfeae0a5fcce4f7a274d48be539d7956df926ffb97a6f8ad19b21d84585384eaef48413b4b5a0a8d5f21178e6eae2b9225eda372899e7a3157aad094ccfc55ca106ee91de4938cf93933723c5c0e4dae8cdad7c7f0b538466d792fc831f47a714095eb4524feff4c5fae15872688cdf208f54ab2c6074be2bd5cabb8acfebfc03b84018983d223e47537455461439923a222e988f285b14331456abed4a04b6d082f85b60bbfc7de6ea0c00d254cc7b0b5091067041a023ed9fb6f8e7dcc2fef33391ad0f296f0dd90957819c58c5a2471f51adb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haf72a8886f2bff177b63f90cd04ef31be1f013bb182a71cff90ccb19ccbadaa3653120da2511fb98e92eef418c53d923f3003707a7a5c06ac1d37a659190f2b882834381237a65b25e83e6bababb132017b044facb8b7145c66e202f47a7e29755b6f6e9a2c4dd566017b2ceff61a50c65a495449843f524996a5eaa81a5c08f2babeeadd1f5dacb6b6a99b81ba37b78fa3dd2413581723c0f444dc00b24901b086571587b407ced8d2f6938a20cc7c34eb27e459bfa11ffb2cdac2132f6cd4873a65fa231aad6521a08bdc0beb84d3eba4bb34fab361185e8e067cc1f6a6b0814a83259f5a32b6c12c95ac2191225d8ca63301e4ff9cb729f6ddbef16a1f1c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbca3e8050b48f8fac807855b59dba44212a93a99d787c2d063be357f485cf0f58873852f6b1018c1624f138eaac538d82e5d85756ee7430728b381b149f83ae386b8b7a91893f18907b7648d661725dfa844251c1a3e071a6bdd538dd872765bba2fddd5875a14f6240c16d8c0743f8399779a253c1e649659051f61895939df96aeab2c9dc77aecac23a2b7127bab0028c113bed5d8ee4ec0a99450777d524df6bd8d5251a62b4913d4015030d5c6685af7f5c67bf830dfd231f0f878a83529101d8b3690b101292a46759247812799947812d5972632d48847bb8d47ddba892b0d9597a0b0ae9a008e9331f630edd00b3d92391b3e527f8430a47acbf5850b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6afd58893270d6afb37e870e6a47f31d4a966d599deab6d270d4541f847561c531b82564c44fb5aabe6bcc849045843d148f90244a28002ab3a20b507e6ff5f93f160400d7dad74df3dcf92e7c5f2e11a526b6869a4049f258b420dedd08af2e07911bdd672675e0deed2f237460fd96ec1c67988150c625e7c8df274a7b3b971a46558e713d47195b3c46133b8009f11b9c8730c93fffbe6b6952e4568b8a63b02eaec8cda8ea5f3aee326a430252164a2a6fe62e613162c70753f117cd09c8956de2ffe307fadfa34d1d7971b68e597f75ad3521f951638db45fae434a6dda142385ddd1a89532d9c9fdb46cb031f794625fe48c1c65213848c641ebdcdb48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hab531cd33d9fdbabd1b0fbd6a737f0cb3d3784177653d517b13a3a4b70a03e8f0cb937982690715e1337f177f4091497e79208b45a11f3ad5322b91d874b228bfc0dd9896605402ef9843f9f8505e13b3fad7fe62f0d17429572b2971fe67d9ba2843515b334c9f593f3a4017d430d6659a58fa24209a9da0b88120596706f9c33965913e4cceae8f05263f373a2a9f3367388cd0fcace18ab055a5b1d9e3a7e7b6c0d8955e31614c50d27936622f13f94c7937587d2815991448e3b41673537a72b6bcf6406530d23584a483115698a62b4271045b1fad13239eff30d0fa396cf6caf7bc2c40e51c3a1bd460a80ed655968b395651697e5883c32f1be7978b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcdce59da0fa5564c87e2d8c1781358868f0ffd035ebe83564ced751283edb1b81884e5c8a6adda8a42920756f29faaacbb556cbebe4dd1be6fc31c39d37698d512bfb6b938a1ede14561027eb867dff6ea0c4c34f73c766fd1e0b58e72d8d32d1c0d3d32ef97f876edca4de754d733f142374ead3759a84a1c4a026fb8b03aa13bc14c982cc86e5135c04ead94dfe2e99acc1960b2502af5da33cacb07c6ddb1512efc19c0df5bc6380264ca19825de4194ebdc2df08291e25a006d39f09557b85effe7923f0173aae354e4b01544e44882a7aa6d96cec6f15130e5feb964161bb52c4d5d5090289f7c448631346c75aabb8c46b52fb33ca9444afb74541657d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h79474616b5ba789ad27f772af7a2065d9486bd0481dbfd99d5844297f426afbc96ea84a67cd667bbbd7125709f3891f08f86af1a52b1446e84d95e969e8355ad6b94b95dd2028d35ba29ba941de6c58399769c5ab5654c11f6318aebd56ad984dfc5a7169c325e113563723cca8f6736d104b97befce29c4f371482f13a4894f0a5a7b3d822b64fa8cadec2127165ac0f0ba562d5dbe15f4fc3d8cc0d2ebe3c2402ae7a26df38444314c6f06fbb40e5b470dda01bb1b5057ebedc5f7c5efb197a3e4727d2b8bf3051743b55a445c36014b1f147221d4e3171b64297d0a8b8b60d1c526b3524186324a930c9f6e007ea25d844555714caf76c024c5c00cdcddd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc0f2a4554e99de6516f28f81e472e29c4695b78f2bf3fe74a14f6fe9b2a38b28891c2edcdeaeb4a98786cf072b76e50c4fbf7016b6eff36652028095578fffb7702f45ba0734c9abfaa2e95ef904fa52cc58d88254c76e82b0d387ec66f67a3678db072d0b60d625b3e1a293bb5c36a2799dde02d5f65b91125ca44baad20d43e7472455ffe5b846942ef66cfd7b41a35b977235199002dec22e4abbbb8b8b23c7d66c3aa5fc94454d18a20d4c7fe9498d15219f00247ea9c4eb135078ffbc74a41b90eeeea0f86f849d4d47b5416251433a02877a518d31b3cb410121667175f2f5855bd4e049a41f6ad521528e7b87e969351f691897e69b17e5dffc1544b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd4a4813293b5e9bb57f997382e887485c0465ee94c63d6002f37c302d05ae563bdc1cfa743d3d25a36a73630eb012419f6c3cd3f7b52246e7f49dccc709ba2eade2c758b2397b5a6d0018d4af8b175812a0a59e1a4f86e7f15cabdb636315e335d282b0c25cc9db9eb0babfa41e120c362f762ec69ff18f211c8c63bfc17f76dd090bf50874ed1e55b0ed4d51f5f6cbb2248e6b791372f2711a043b2c139c66222ccd0788914e24a2d8e50038196fa2432d8e8a2f82dd1de420c72ecf518696f0ecd4a3fdce3b61ca0b3efe91243b2a37019045ce2f0bd4452e3c0361e6bc59a5795551cfee3a833ba8111771c3e4c5c20a1f8499f28c30e728c3f9271851ec8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha22587e08ddb73894ff0a5dabcb41d276444f1d9c2e243a6b939b373510daea963e2f853477a6b1f7ae0fb19a59a4eb0a4231362ca1a411b6b949d3b98296dc74d5aacc6bdfd4ba64db8ccdf855cc01ce2fcbb2ca8f697f002e18e3b1c05123033c763982ce2f18382f5e9638c73f1d2456f8a3a2870d28510289c5f70687015d1d321a51baf0f620cb98e3eb55ca43dea7162e4d8f19be468b3f3db1347370901b89c7d0fe3894a9ab733634cf7a8b1286a81b843775cfa4efe5037c6c999397d480f6f32c29531e522a562e5fb278ed58045f7b590afbdb08b6b3768ef7ae7737a3a3131830e2fcc79478cb8bb606402aabdedbed5d40b97779ffcc49320e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h19c464a90d296e1ac7a89f9371529440fe4f06786f92ac7ef80d18b9bcb2008c94ac949b8cd35c6991d9f7c79f220ee5f937e9100b9a7b0a9b0c8d4cb0cd0eb77bf02aae88b2157fef4b37ebe42356785baf1e5d359a886e4f24b2d86ab606c76ba3aaee68f2f7f94b5cf936468cb3e356c9bea36193350c82b39f7d7aa03fef445a8ef6ee87f9fa4ecd41f8e8b7c6a0d573795f5140ec8e773b08e44f835beeff13e52f6dd3d2840d3eaa98a056108678141312270cb82a35335dd9e8395438b2d793a1b30567d7ec772e8506bf12c5bafe5ccd8ee79a2c76d4944ef965777bdd8ba04a20165631fccdc5555a4c5e5dc67589f029c2a31a21171719079bff4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5d710a98952a150782f10e52c2cb58b187b9cd148f2186761cf5b054ed1d04aa34cb0a673ec8115f87ec98a3421974cec0dc8f82b0d16a04f9ee230ab4557ddf886756ca041f7e580b89ab4624994400a84647017c36f7f18c3bbfccca6fed92f54602e80ef4d49dddc57c132a4403abea3de20dada2fa8f9fe656386f49c22dac17dbe2efcdefffc343a5077b4fed5145143f123a545c556a16ee6fc609ec9f9a5d717be9e6c6333be5ab600cd4a8808e81d166477943a28dbcae1d7faf772e9a7109accaae4550e9bd1608f31d86e5a0964407f0ee1f0396b1b30b2e1564eb67cfb423e37214940219d9f8f99edd1edf3d9f1840ec1957de3fb43ae974bbac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h99eb255b663aedfae6a05e9097ec606cfe3a5b3be21d720958cfbdcb51d9059905e1c88cc39602c0e1619f7d7ca884bdde268ec745f5ee7a257a408d37a1e684abb0bd48b8d9b959378b4bc0b70e366b4ecda078c0c07e3a3f008a7648c88b686a7cee656f8642b5249e0e4b1af1dfe9f66fb67a477b568f106007be8db026690f89584d03bc3702a3b807c1f066da93bc6d34ce98e3614c5e04e677fd21905105dbaafd2d9b541744b0f8b54e88b23e968ab43bd0d8d711263490f642c8f151e360642f1097b3e66b4bb5b2cd19f2b7d429fe1332147932514ec7965e4b54a2c30823ce4a79c942c6515c5c25fa4fce930be8163e353168f00c13e5a7707653;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd86f074704490b788d2dacd0c08acb217d5e69e25399193579ccdac398e9918dc85cd8785f7e7e05713c49f152f0a53b037efecfe0a8af5d0b2c7c36f82991242a5d0ea0841a0818c28716bcf6a731b7da1ae6212d6a488b83d73ac43bc287cb3d6d7751b24ab4050512a8ce0a0f889cbebcea865eb0b3633ec77d95837af062da233df9161c39f96e20e627cce0c5659edeb4d5a1b02fc0e28db6d3d0a6d1867e497424e2a8fff628ecc53208431fe283753c8d4b473b0f795de40be804ccd8a7a19d70bed803ce83bdc4ad9a43a7a4599ae9f75f05498e4becefa26cc5365955028672a268d8f2e5fa25df7bd7266fd7b154591dc1e3afc68164d8b6f3d9eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h37de1261570b47e109599cdcab56084e5bd7b0f3905257ec7da64e7652098617343b53d3247878a95636189c2d8833ea60a941f2e4cc3ce9850ddcd20a3effebffff4303873aa58ac161bad3be19f1c9cd9612975b6d7c476d07ba1bcf5e220854c17243c77ab7b212d75358f1117965e278fac60a494004c02cdec4054df822812d9ecb1c787410d02abecd88665270b973fd6e2c609c2b89c055d5c77410798f4169c59c818796fe5415d1365737d8d9235d77b4dc57106240c6b9051dcc8dc5c0db41466e1443f6feae737006e55cd9017b657b4d96da8b0099427850c1919bfe342b67ed6a97a38451362cddd3daf9294a92904c50ac69e60a6ce236f585;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h94a786480e518fbb09c7ac5e62bdd5d14dd33413ae64c38ab36359e3fd425d969aefc23c3aebdec8d60c3047b8b357bec600f8c2d330bb19a0c854dc58c065c5e3c74b9959ebb1058fecc6b669d331478e52cc043321ae74fabfd44d6e40b92bff9a04008f6173ee531aa5d86e9f9997adc4afe3c995161b45304e6d9bcc3d7168debef32c79bfa5dc5595ac3e0950d6f42ef07a7d6b0f4731c6e5f76a077f58f3064a0b1078ccb62ba4bae8bac8b8e95101b4bb0e89d530cfe62ddc67ca975dbd8293f071c1c482aae8ef20968f79599b512eac0659e78a6f78a22bb013b634ad81729d55338aec0aecb8a3efb7e44a5ebaa8a04c84ba612038743461b18b55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8ba4bcd4d101c73ca50f22151d52488ddea69c1377b2e2aff746801c8fae7b4190b5d968fa4ae41a4a91668e7d51e4df5744fafe0c60cd9882fc1f17081ecea47c93d9299892dc7d1a14ea3c58cae09554483c8e98b673e1981ea54f5dd503d86948fd58e691011745e4a6f254f09857793aae7f8f3bba127b488ceeb16307ca8aa071ad82297295f3d16941e7b94bc948d2f095dd6bfac6024834cec99bf4f4c978438304b0a34ef2bf5f11e559494d10085a1888612f271e975cb9bf62e3f363be02e389279ecbf5873f798d041867e73d39a288422de96ece1a341af4a9e699633435672ccc0623a698b638202d55e8c032bc8a3031e9bb788e7cedb09809;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6e955de27cbc846d5b50ac0195c38b246cf65d4154c7f9e5cf640b93d3c0bd5d127e50e0c2f6177fb09762120b1978f510b63d503a423e498d60fb7e861fa3ed94f5a897fcc35e46e09702378d016b90c5ae6b7d619ada136f07ae0a0fd016aa37310d2b163f045b7a8d1d55fa51423626261c60f0b7e670b8dc1a68dcc3bbfa15eff8e80eccd0c28ffdf11fa5a1f17d4087ebc9a5d90c81e5eee4a8adb36043512a2ef5c18b5fd2c43282f75388b5093cbe1724cce8661c10f60b6c870fd38fd99c66b39260482623205f49b1afc88901b768dd0dea80b6b4147a9f35e5f9320d54a8d63e823556d3cd2418c01ccd93ef9851438fde06bbad7da4719b9d1b30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'heebd1e095464313bed762ef049d4a5fd1bbfb4dbd201e07ceebef68e6ee1e569d313ba01023612c21d66d59915b97350e118544902aefea5ea4e506ab9a07b060d8ad9ff32a034834305d9902d531c3503964c3c88d1af23982de9358c8a17fa42a46f81c85f1f034898ad6abf5ff1adfb0f3b2a0748349699d6b8f2c9850b9b233a2d7535a57e1433926c1e1f6e2b9679e68326484f465ee7ec4d5e0eeab1247b4ce424c8ea52c05ec066339ab8f5ef3d54dcd942404bf6c8f615fd897f87278bbe0909d724ee20e35073a7837d2598de453d78cdbf1e7206186de55ac5828470c5e6fd07ae5bd436583c46525944300728465bccef732208af54779d7728f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4ba78e4055fb028ee2913614539ace1cb8cb3460b3f9ce40abf443ba4821563e0c43efb6deb23083da488c9109033540040c24d9272d562d1eab4233123bee11ccb0b37c8fa8023310cc4eb892686e7129ddf46cc40c19501130b5737cceed23bdbd9b44f7b3c9b68104b40f480fc44a030716559364649552418d6fcea16f9f1d96a05bab1198f2211ecfb75d03ef266be9925c56256fa7a854bde987669e08a4ba0328680e5fc87d73cb5a16ce12923ff17a4ee1a8da526fda72bb2da408d2b917637cb863500dd85b02e22bd8ac4782c2a24bfbca86af9f7ba0c031006d7af92a2dae74dad0689c5b6db8bc63d244b8d3350fe5d9d355c2d945879199e1c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd418c6e4c846da777121c3ba6dc0f5cb0d4c2a3674911fe3b85a69ed95785a57aebbf93f319d0cfb306994e41aeaad6d6a10e02e8ff32e09ed3adade37c6615a61d397051308a6c8ef456949993477d274e8739a8360ce90b7f987fe92c7e21c5100497f6516ec58ab905b921bca10356b322d0087bb4706a04c72237d0b7b2c358e7f38df852559ebd80dfbb9791217d76468e349ae4a65795e7b1c4adae54c60dfd2ebe326dacd6a9c7b784f240b879527eaa11a1cccccffe181b88189cee1d45f9e5affcfbeb139efe2691e119a3f17d7f4264c4ab0b2a1f57419cd080df63ce648bcc1172e7609046c19492efabca45b08aea55ae0fc061a86075603f3ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h138f850a55b5de1a5588762cab8850aaf45606b5a78f0837f1940270fab0398dc9cbfe945fd319b07a35208ff0169c5a38ae5b82bbdee3db482933dde94f65904fdac4d4ad57f85c518d65d37dba29714038d4b56ec3f3aa0f6b0698e93210d6842f01b9d75f49b3981c484cf27474dc594ecc7781a0363595086e5fc0f2dcc3d9df551dc17f3840a61af196008a234975052631ca92e6cee9611ac60465425b717676c26848b91a6c1e779b36e4ec559f4cd9a681f77a07f849580d66bca01a968907293917f7fe2b4396b2f373ba4b13eb05a17ffd71ace1621ae2faee54edb5c97b8b1b5c636b8207640b7e02e58eca8798f503faf74997eab1c972ccec94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd9a98a0b587dc60e842ab564f353b92d3515dbf2745345645865f357cdadba8ba149c4206b43f66aee8e7b6eba3185c59e2b74e2f68fbadb598d26dcdb5589bea5be529050466c5486ab5f3c0df09f8db727b464094703a746cb107e7625585c1ad51f8658e2adc5c288d48f0d1b0dda5b063514d23a4fec0b61a260cc34db6118a09b18a1fa7fca7ff5d469fdb17ae8049e5a9fdefeaab41238fd139179fb2396b8e56c3153120c7f11a07391d92e896b1e14e799797011c876d3210e11e4d25355620172470642a9ac71b6ddb322af86c0677d8258f9221a20238a9add453c89b5874857bd728d8054e4796be217d197936e7185fff30e9f2c1e7591b9758b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha1ae1db848a638e1c98b0baa1e231bc9c8599988c1304681fc576b3bbbaf43da4217c7223126c7bebe0e7d2c0b45872aa1145bdb0f6e1fbdc6a2c6739d917eb043b20d47c9113540292ac66682aaabda0e9afee30cea0b17725532eb451151fbae805ab32ffe927db36fb318eab1f8261e25ac908c6f7acada1f15bbc804f82c23475cca66a24ed5f7de378ef84c61fff29bc05511072e98113c0e94fc2a95b93ae496ab9d8c3bdc494c010191924f6ff392977c6715364db813591be9552b6227d3e96dd3cd82a5d32f67dc1167e47abf3189e5c5fe615f4b65ff25b1f7d47e1792eb59fc4065553ad74daff4b771695a6bd8dc4b9b1662101fc4bda5dfca0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hac68bbe8a8313d279abe6278a88d964b1699e607cb22b5cc92cc12f6ea53d1b04ea1792c7430fba949828c7498b1081875a769acb405e14dac9465034fdab898ef861cbc0febeffc71232f0bf371a1e2e4a78b21c4e0f9b4d0dfa26e57959bcc5944ea199f4df29dd5bb720e2380c17cea9349458edcddbbde4e9325e0eff92cdb3463d94738c8eb98ed40c7501a61f7157072e670c1cff3a343982806c4dd5bc272df9928893770010dad97e87aaccc64844ff144d3aafa1e1654486efd97ef417546e0afce37dab0ce0995be54665ebd5ca7b064597d951be213f64b61472d0638058257b350cc2305c693dffa390f6cff1ef74462d77a68be5399784fa54f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2697a26b02c75caddcfc3d61e74e0e72064164e26209e65937a4222dfe919dc5f9416e3d13e557bc521461eebef86a42838e89b93806d21f3e4c665b5fdc4c8697920076179b63285117ea230b212424269116f77cd66d2f0e0812941bcc6de0c4d542c8c5e70880290e50a25b5a35e5dc7eb352e9727ef255d6170f11cb818df5407ed680958d9570ae19b029730f8b93767305804bef0bdf0b2adafe6ac47e5dc1e57cda10863c3eef9113958c8ef07ed7cf3c20d860e66d6f202c59050f07dbb2da1c01cc5c14b7493b1dcbf428b534d0fff937438e68403bfebadd6c041b0b23279c4d3cece1e19bcd322c276b07abc57e4aabe70d819f2018dc09a1b8b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3d201936f6036d8024a9067410662bf7e3a0a1348749c3e5342d98246e4ee4c5563e42bdec8d0554ea47586c6f0a35a1e79b60f7a0cc50ef38bb005163e8301d7b3a4965ac7eaf13c27ad44273325f36923274c05921fa9af6f42c9ded071a5ea61fc4ba7e7f5ae51d0aaaecfe796087582a2fb46fe5b425311c9d0026747348273ef95d168729ea6c306486a75fb723054c3bb47fdc61c81a5a856614885348305853854fa81914101ecd7bc6fa255b48c1fdd5813756a027c1b33d389a301dfd05a0c3fccca4da5f02c7c4ac92722ea3dd5aabfdc4fd7bcb773d06a86a50d58d1982fc19ba8e62acfd131924a6f31b16fedfb89e92cec013df4f6fc551a976;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h24f9e9e5d2cdc9feffa1699ba589985eeed85f4259b2cc599255035ecde15e2ff313450e994fdfd291211819a5b8dae8a8cfaa52853089402e37ac2debd2e004fc38546e1266381b898965b149df0462c228efe17f34d280069101c9ccde8590d939549b65b40d9e1c55f0e46921c0810e276bf297bc70f4c20002ab706d1ffcd481050e3ce0909f108fa466d84ae2d22c476757a6a5a6812d8a7d84051500be91f192f726991f80b53fd82d0dc63f6f89a9f614029afe74e3814989df6b0a18981318f4c76cf9706c7c234473e5938ab61b6c712907923ff779fa19ceeaa26b79fb00fcbab07ea780aa121fc1fb7719edd089ebd6d8e469ba560c6992f3659d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h918e948c46b1fca3726530839d20f209a0b745355ddd26a140d9fdcda9dee441641e35622fad026fc4eaa6d403c5f11429c40066deeb98cf9f5ce772c160c470171d0c25e5e53d0034f8be6e48d1a3d66ac18ec3421f1ef7dda60b0f75903a57962631d8052a4c7e132d03ebac188ce3fe49f91161f9f880bdbb78acefd1fccfb94b5cbab6cd13b968456e7452f6ef0c97eda7c81349de4c52f6fcef66dd4e605a911e70759d6635e988b21ac73fa50fcc654eea19468a734559d83975252302eaea5bc73b053912d3b64d391aada5e70acf233ba14219bb11e32ab3ebab21a8a0fd14c5ced566dbf0165f094a7dd67afe4629aabb9618e1c73339dd09a6da3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7b762d4da4fbd52cab652bc218b037b4466da1dda23b9bd47e512940b5e8ff937cfddb6bc4e2cfd5e988a742c6d4aebfe9764b6ce05adb4e5ede6c460fe5298ab3a1c6841eed4687bcd5d4a4d7e051b0952e3f161b4093be6c1d3a00ad2cb420f3afbd96bcbde2af6c4aecb61b2167ed932e97626a11d1f54c3ec4f799c085f4330ca150bbe5a425ea6a092f164f6e18515d915a66f366dde7117a5a9126193d2360e0d670ef010edf84b1820834c2d6d7042ddd02aa138b5ecb1f841e8d6de0701099594bd901890c3664aeb8d0404671d3192bdd249e263c3a954c23133bef650fe9b5f38cd681442b34736e25a2cfd38812e8a1abbc5d214655103808645;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7ce9e43c7aa345a95ca552db21272457870eafb7af779fc6ee058c469a8aa5eda035876fd3bbedbde89f794027ca5214986f8182c429e8029bbac6a3b434ae22baaac38174d11b8c13f7f5462913f5e61b86e884c21c9d8fe3b0a2c289a8d2bb850ab478aee2797faf29aa4055040dbb139b0814a01586d0ec41d8696fe365618e2570064048b2ebe83259eabc1aded588a01406930387bf21e0e1c5eea8ed9a157630eb4f40946f986b0d17e7493cac19b3bbf24da5964c778c67b3bcf79f4783e0e3a643cc5a55ceeeafac0400e6867a50856649a5ba806078abf2806f05560f5a76612728adef53e3751ac772f60a3dc59b106dc1565d566796c51c7c21c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8adf4f9ac0e4df88370354ea5e754d39f19f8c49db5e2809c19ae579dd00b5b6a66e147d0dcb704a45d7d37573054abba0371a10a3b6b9eb32bf78af0b1091534170ab7bde249cb3f0a282565378a1c588bfac0daf88ab8eece26627f04b3da5bcfd9c066194516ae59becef101db41bb1990c41bb342f62eac821deaafa4b78a506c4b29923a38554111c7aa0ca4187aaa45b9ac493579bbe334d9a4f9caf197f8e9f6958417648327412dc32bae2f4488a5c584e1e77e712f7efc079236155f71e41657e78a7e35327da0d1bfe68333d528d61bd5cb90f1bbe008dc501dffaf1f8d4734b37b093e1743564514b85b6fea077dd7745994ca7537b7d92081ac7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2481ee01deaa5cb2b5fcf14dcccfc174083216ab3524d4c48902accb6d30f2ad83ddd651779dc7e92128d76d75ef4cc2d4480591ce2e1ff55888f3c6c1ed4213cd54e82dd47bac8e57843e8f5b64b871ab20970e8be0e0be56c83d9c805cdbde3486daab68f2040b4b7e5998907ad7edfdcc2a1d392b87a6f484ea2c9e639a4dcc70ecbc7a67c894455ec06183c49d9dffd332574362eafcb98c404b9a6f1e04dabd465f3685b06916da8883cb48063cf5769b162f2b3227f2d5ecffe542029ccd482fbe3654497cbedaafcf1e388529c984433f4e636792116e77726d20544892c00854da96ea001c9d006599ec61181444182cf2f2bc326132fad00ca40b07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2a57143787861a04044513ff25e17edace3a7a3617139314046999bdb0f32a214b20246e295ca3dbf720d6b89991f5646b85bff719cfdbba46da66cdbbc007121216b5b502f571251102eccaba5d6ad1cd297247ecd180ab366b91f58fd4021f80143059a6606225248f354bacfc8b3fcc7221c6e846fc3c58bad11933493ded0c12869bef34d6a7c18b7d4107c688669112b4da4a8836beaf7d52ce67d25643aeae28abb229ed7107435cb25906eddf5e9ca7c930d75c85375b7a9484ccd60b328d986a0864830d67e89898bf567a4480a5c932582f8a9f460194e5b16d3e884ea5787c93cd5555c5226ef54c2803172a3f1466a2fa1067d0b8c09b7ab95a74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h170d2cd712d6e697abe3d3b059a5348d3a65bde233cd04facfbffeea962543eddd18a49f8cc37fae5351c25cf25d2b2fcb56f063a1b4492788d2e7870e9f94da6e8017c791c803a586316c48568275014734d9872e186066e897a131eb839cddeb50cd02bc2b4a315a39ce82414c80664d51478660effc183ce60d779e142cb8827493e30f66359f67a9104cbd383a7b26db32b7343b614f3f1a8093fda09d41a658e921e63dfb315855a531baab544d2cb95b04247ad877dd9302dc324cd5fb2badb8d2d96c8c6f3b69d1f6ba54126f692d79d78bd08cd022bfc6d462c6c8f56634e7dfd2b5b5ba5232eaedaee6f8e7dc40878de1af9267a389d17011665146;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5fd2e2f191ca4e83494266a944e1193cb40168647e0c370c8494ce2f2bba671bbf69c9457b4d4f167eca6cc8b07ef96f179b3be081ab8c175c269f38c66267a3a46060a61f83073c720f342a64b27c073e4f0df41274fde00e35105645a8086e9641d3fe3773e2507969af0f85a73e5219ab9c1df555b2db3cce1325c1834612ff0ae2b4f86f988e80d68df289bcbeab47b9bdc8ff232080c4fe004ab05218c517d5735be252903800c3f2a1c7bdb87d3e6efd09edab5a1aa8a203aeb4f898f4fda0e091a0ef31c97e5d635c1069357a63d9d36da7bea54ca374068088304a210cfce5aeb5190b6849ef6191be82b25c923257eae2d1115a4646e37f02f12e83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9a97f9bb774171a66e0cc151ff018b002ee1062402fad28f094ab78828fa8b94b52c7e4f65ecf26322c6bbc41d92dc8c466b686a22c5ca74a084173da63fc4307d0d949d4075fd22dd3c8908c0b28085a8e04f12b4e31ca69027d9caa76be2340ebf1806454d9ef186db7c5093549dd4be42d8e4e26c906cc0cd94047b1023b1a51484cdab378d79c3b140833a8536fee5aa2809e349b2969d7a6cd7d4202d1830b2cd1676214a9a7df1ca6e36de5c8eae274ab343ae8a7a41a103f4565aa629e15e83cdc67210d316aded4527d7ffdf51917123df6c187b64278d4d8b305033eb848282161bc12b3ffccd76db464a821b8e15472001072ed220749e6ba56eca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8e607c6551372a4b9eef902c7a81580795c57d9ef67952accb68f0b75de08e0e07720ac7d84cffb0740e8176f7547cd69cf68ec3fe679f270b5d16c812697fb22be0142801e6812b6776b12ea0607c9a0f779d7edcbc6ef22837db4fcdc885752899768d97b00f143735980a56548804079bfa22e1cf83b498650c695a3c0f847eb67223be51703c3244df11091268300658b75ebdfb5262a8a68e5aab9c00d9b4a047e0760dba7c58b634b29491d7d6b7731b75518b26394a967bdb620a0d5001b94e92aa769f6cb7a9903bdd52e6fa116ae7839580161b0b5e833e2de7e84d225359695d289ccf9c0c52a78fb42157e42aaad01038f39f499d9fe294306007;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1d79da58a77b44b20a9d689a4855fb823a35196de504f6eb442d8270100973c38b1f93e0a8a7748364ea8fcb9787f005fd3615cf07c85763191bb3c76884de4b0ab3688f425ffe18897274c6a797ce7c8b8c9dbfc58e71ff822056e7ded4fb36914a380bed664b824e71aeb1407dbf83bf70b8c9bbb2d36ece18fd9b798c38627ee524337ef7ba65e9c69993c3ee2c1dcf46895a37f6309ed20edede4cf034bd161f05f938e11fad8c5952f1cb0c110f982feac5c26dc076cdbc2a6cd32de03d1de491f5bf071b23ee297e375b5ecbb994be7fa65b925aa8e5dc478f6a5e28e77a652808cb3d641a5a5d5d243bebf8514d5765c3a210c141f98473fe4c6a7ad5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd726aaab604013b9385fc6aaf5411c998a3e76378770da629c76cc016db513899f50c57b843d42a95e84e2a6864720b211a8c3c6a36545fc638d0af88891cf892bef6a9cc63fbcab8b5e74d99767a3f1ed22197f9e7de1593d9d13644ad36104510e3469ba65a57bb4cce1c948fdede737f2e507f2fd234be3516fd9046f3401cb7c43610799d4b9df44afad06019c734c83ecfa048c14345b210ae391fc918da4ce5b2875019d50c25fda0c52c85aceeff81dfd3a7e479f04cd0ca1757cdcb170b943dc87c03ab7a8cdd4603a36067b868bc321585698ec7b9840e44147109a4a5841fb94ce1e28515a1c96a6c93be08efbf0d5cb3c4ba75f3fed9f700aa952;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h13802f2d2df188c17cc94ba17ea970cbf572ff5bc3c956631b1b6ee2396d1be265d28db88022a2399ad848ecdccb9e84a1d0ce5b2cfbb0d5c6866a79d9793376282b5d620d65c812e76b5db34f1c397ccde349b00e866d3af8b80ad9876f7acf69164b8dd52a849bc067c44eaf9e9e300f6312f4a6aa515885f1df88e9fac41a26c51e1c5e0e4369091ca1cce6e0cc77e8957751464779053e31ee374aeb2dbbac751fd08db0f5fecb6ac53de812a16fd541d6d3830c2c4d9c31fbb27f202f8c61533b1cd8d7ea1f4be9d08a052eaae96b6a928360a392e067a19544a91b28692d4c4ca02a021b1b849c75ca213b72298439253b11856230028af225ccc21e41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h733fa5ed9f500625d9052b5cda258aa9ef3238be88b501c7afc2ceed89678e5f9cf8b5bd051a01da50a0304c20d7289ff21274fda1a193c8620729f0d371743d76b1d460db29efac19eb62ca7d08cbf1f175e7b063c8e4160030f96f78161c2f479112ef083c562e6a4a2f243c9f89296c919778ec5400119a433b4061f4e5551f5af6730fd48360fb8d622e643fcdbb2af251ab4640c34af36b39677206d7074849e0c55f9cd10043ac4778720cd0c84282ab6bf6fd9c6e8bb35997e783deb5b52a655bfeb2b867751c25a0d64ea206e73bf5fb0965289131d7138efce8a162dec5142b4f56def8a2695071637681455d8f1259fc8e07023bbe2ab81cc1fd54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5855ba4a73a8f883155edb02d69c0a3249c44d8f7ba7576b9558f7dfb7b46a574bf99f0acf269b7ab8792f5ee62b64ffc9abf7718f47739639ecea387c4fac98c0a46bde2e112a451cd665b2fbc7f17434a1c060a83962a48d40981f6d28847cbe5dfeac789f6a78c018417f36059c2e040576caebb477b9710f052ea28976af83f52e84f473951fc73c7541f0d6407f40cee242fa1f4650c772bc33debc1270ae17939b962e5f1f14a47f1edba2d03833d05ab53a35ce511dfea9ca32270f363f180a61e8232b9d3d55df93c8e15cfee768176f384aeb4136995ca6f7780252552d37c9099efc57c74ff668c50a47a1b417a8ee6057f96d7967e0d1b0c8102a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc9fd9e62ba18b7ba576eb3346bab611a9e237e73b4d4551112bfa3495f65507c867ea924fcde428585914cfde03a70944704ada3dc6c3ac29b8f0ab8a823aa78f2e3d20d1d0eb2ba1be2e47f622662e0f0da32f44d9a613a50f770b54b1b2f61c516247d6bc59c66e84d68aae3103de53ac6a13fecc50489958de8cdc7122a32c25bb604e301d47368f1695e991c767bb66b06a02e3a27b4ee8c48d11c0ab8283c1f1f128c145d9db3fb67e5e1c748b33bb2e01541ce19dc6c0b15be5387d863d7d1077b76503f970fa1d1e7111d5810399fc1f38878c95930ccb366a52b3b690078eb04c08c64da0d612cc907b449af45395669ab32aad86d4d7a3399c5eca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he3fa89353f1309983a4fcfe122f5c4ca20386763af684caf70b7ce77ffb6c0144ec58d2701d0c4214b472f0402e8bb49d2a360fdb4a1bbcebec9ac846c4e1e29e875a43920865f9bbb9d5c413ced26843c632a3471d71061ca99b3967664732a3bef9b275b98beec6c7647639a71cdba01484ea226a37acbc487bfe58f586c05449000a63b157d7ef86eac9df331dc5b62d55bc543c2a18d1d2b219aca20a69a8e8bcbc4b621168b670c6e6678899e59994b4e84d2ad9a3daaa39b8205ff9d36a287816ec7c0deb977f0ac7483ca274790fa27f92930eba741a2747b1ef6bfa8934bf3e53522d5b85966cbcd92df87a77a03b9caa14930be0d2386c9c7c5a461;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea3792211dd9890c5b9f4fa488729a5e383f0df3196444b0aad6949ba111691bb698a2b810d167d7c19e9929598e59991f474f30bbd9d7d154634a2c138a5c61a919d529faff6ac673709cec83c7e233fee8f0260bf5af4e5e04d7f49b6ba8ab92933a47173ff557e80a189aeac5e35183314a913e1e76a1a71266476a7d003eda3b6765c3cae9e43364c688c9ec4b7c8b9419106b5c9bd41468604b09a3d2b422285ecdecf5333eeb2040e10e3bba3b5a23c0a5a3476f655cfe1b133a79e0084b8c82055c7f096da41196e3b54fa6c621d8252190e99d48d076af7eebb5ed448e053feaf4b27c694175a27540d50d8fe17818bcffaa9ac73dc7d6cfb62a6ddf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h961535e881b5d01e69038d6c98a7e276c6fb025a199818d6682c6dbcf544d1f2e70194b62d6853f3e01147b18add1c3b8845a7fc281007f46af6049f17bf4bd689400bbdd6623bc7348aba7257bb175a359d39043e670696ed642fb9d795565caacad59abd899044fc9da87c3a5a84ac133b0e7da08a4128cc5a479be6e9207babbf243239d992a79f497ec9fb384d45837412526378892a4f54b20642121d92f292718506fcf4cf5fead596684792a21b08016c72422645ecc3752af93f339ea8304b645a30e3ba71dce86efc914536b6308a314b1e503b81de36788267f36b02feb83a68fc01c2bafb51a599cb0254703bc78774803bd52965007d77808fe0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9bc7c550c021d8239b4edf32e173ace98d7b6a400af3193688007a2719adbc730a7d15acb8116e0eac2a04099a93156709ca1fad0f950791cc82b7874aeba260106726950c329203d40609f774e7de8f48faee3a73f521be518e3faf6dce7553f8cf78ecafd8cdb5234f969acf91e7dd3ef7aefcbe1e21f2f911ba0f7ffad7261d57c61cb18eb93aad9a6726f0be82b0d340cb9edb553457bf5b50fb8dd1d6cb7b08c4868d665d24f2ab35ab1a57903a36e76733a85e94e443e30d27cd7460a251ed546ef5bd9cb801129e8785af19cd38077204201458c52a591d8ee8e5838babb8c2211597b0632fb713c6428a0971455570f50fd38966c28251ad47d7d7e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h102dda752ebdd9d98de963fc7106ba94475dfe428a9fb204acb34f612459fc8efb78be806090aa46594654431aeb5d9ff7048ea823d2e5adbb702919b1bd79f9beb9873bdca53d71ce6bc9d12349962517eb03ab406163694a9a9f8bc2e5f0fe761eff45d7fd9af5e23e7732ef6063531046fc40424671cd5d2d751f18829d0c6e43ffd50a07aea0057e604cb0f159b1b8f12e890fdad45b608a27e3aab654d6625b50f797fa2f379c3f265eeeb89259b8fded95c1f628df56f7628d71bfc83fec25ececdfdbeeb0efac96cd7f601d22c7f612a194416ae7fe71765f7489a1adf60154268481a15f0c6c4ab2afdea78480b1631afa375a7efe8f472cb8da704b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfed50f68129317a3f9927aa820b3971cd7023be225d5159426b4dec3eaf54cf881b8ea51fc609f83a734e51b75eac53a587621b3b325e7f6a9aa8d7399f286f0deed421d9f78fcc496c763105056f553a7df2a58ac24e182147c998ae7e42bd96d3428419c0ac771553d83b556182d4769de54de7ddee7024580a1f2ec70a80c5be9895f59f273928fe9b35f3c83b55d173b6eba6e2e26b17c6c961f97e60b6442e07bdf44ce2fbe1722566d5af3378ee35e138ba9cc833e0ab7fb38487b258dc654d332d9863d5f69b6bda7cceeb8cb9f889aec3a52be46c84d4b39f5b8e84db77d9e709fbe1faff028e0d54567443714ddfb0c4c5a49124c10b3127d4d6936;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hca7faf50dc8b808b23252e2f3dd356c21bb766cd5b1eb2a4bf187c03b4c6c55c36a107354e147bc3d240e28cb9c477610ef6a44720ccec45ec0ba742e85d143f9a423d71d1c80c2dfffa3e814bbb2eb4bc7378ce3af85594aa867a50a27e845ac7317beb19b9ecd04decc1b2ccf645ea2e3e48570940aae94968c02d2f4cd39366c8864150818f504ba14386a6e2b3584a28e8dc83da412be7af70b748f41e892417163ade3b12b72e7d03479067b0588f2576b5af34cb52f73162e46a9bebbefc3ec597c0ae6b6b7d33ce8b871de326d4f80d657a8e87214b563d662302fac654a5656707ab7c5509aaf3da5001fa2aaed65f6baf953bcd243bb59ad77b7804;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7f44c4ecd8bd483828689ebdb23dc83fa01868810fde588dbe0fb1d7c8fc5f2e0cf114805981ff634e705c4e1d0ca4da50fd8c000aeb7e80d57a1b8c224f778da2f09540b8ba88cfdabdf0c530ddd70a5e500310a6ef782b5d372924bdaecf5a114aa54f263ed43921ac5f9ccd0a8f4c7c292e1df72e6c3c516b20090197c9ba20f298ac8219da2408684a9ce3612b812e23858207c70ba20d09b9bf40cba573b00d1881c9a7ff09dbac15c2457bbf334f0597b6e63303d74925b853a38c8b47e08f54997d143a836e8741535371bb49b0fe870cac04d907ce3138c34ff474e9e6ecf47ddfcdbb9dec1410f82c943a81a106ab5f6e1f7a8d0fcf0b4b5255b39b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcf805c19677ccce3a8f12121cc2f3e9121c5771c5effcec5112eb3d7f9b1fa4c36dec68306f00702fa6464d6b3e7356dc5aca98b748d3fa9dbd1f92442cf540145065ac314daa9cc1073dd9911b8d7278eaf2d230a1edd11757101fcb7d707a3e15165910ec1c6d210d35c9f4f5d823d32e9886cf8f812e829802e794a7425a367bec63ecc0d444286cc1b993ca634454c571d1f361f112f7ed9fe9cb52964d1e8c4aebf935fa2a81ddb7efa681551bd36ceef2a4a89db5b32cc5a43721edfda608a47dbeeaab384fcf515088101198a6befb4daeb1dac5acd1ffb3d08f717ca6bc8bbd629f6f9b88967cb40cce2e0036f55d53105668d6dd0d70aa81842e96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2f806a549742bf4ecddfa05335a5ab0b8085757357318b1724d9ae22d923dd65104f5ccec799c4311ff406f7916e9a9e63947aad0b5f6d187f1d9e73e0a620625d89009f3964cc0f13122d7f333b91dc73152617d02cb68357233aa744247ee1271a34cf15d78c22094ac88cef4f2727bc5321591d8a9ea6372ca8ff9328a917a63e4766ff919b116944d2cc821433e0dae4cf182fef5a39e53908463f8ee6cb5e2baeb202e54c17fd99a34aef759a50901f848cb69beba94b44ed92a2b115a398df09a5a67adb3e6e0cb24c463b6fc294e5fa40d5a7dcb6abf35181233d65eb413e8af1d69e6e30d947d115ff145588355681a015b1c2c19cb24845b19ab68e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h82cb6e9fc3b9d389b1fe426b9509a671ccf945f9f16a1cf9e181c7bb747719bda2d2addd2ff046220f3b881c4b2a3d0f99779dc4c41c94869f6ac70f0b32edd081b7a98ed365062f765b7799cd8486f4a05ed05ba4c6f13425a68497b30caa56860e68dc290422364848530cbc1ba0fe91a96a5ac3d196845779b805636f659db207db3fa3d31c3c60047b30e83c6e61972950d78fc923ef32a0bd1f91d0a95a17668dc400933e127107616cbfb9b119c2fc702bfe1ebc50400d1a41942400aae9f36efb5c693ca8292878dc599c4379b36d1c5f74bfd37330183496760a275c4faac57cfe168fd9e867fa8eaff290e46bedb4926c4ca305d379666dc00d2fb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h951a11b5e7a56d3269d12370c3caf18ea6d8f2033989eb2791e5c6f09105a39fe47b05026564b7ab4d6f6f989a593f01541f7ba5ef395a03806aad36906e8d8ec68dcf34b8df42a8e27a6f34052e6568f7ce25ad4ff45cbf16136f8279bc3ba0db5e9b1fa2f4d9103a46f88b3e8d990649b06472dcdb3644f2368b3e7d11b0ca65bd6a1514d582da37ed8a57b53f280ddda2e30712820974f8692c206437e06c0dfceaf8522d52b847733d0e522182f1821817d0946fee2c00bab76bee25f415880557a954d9e6709f1fba0c3a0613db3d30472e4ce25cceaa8892a38525bf4d2dbd49ef610141340f6d7296f7f87eafd882970891dccb5ebc4749c723a82b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc3016953b82a736e9ad589430cc4013f1dd6149d8d0123a560ea1274840c66a371360558093161814a6ea941330ff8dc9f6e0762563919814e493f62290481fac7ec7870109957526e06a21e02f4496106d1407c43b2c7c0c41b6ad8c3451af5c21f6df26d73a02cbd65a25affe05073f2cbe2ae4381dade49a65cd915c4f61d7303f1a1faf9764b74f5ca40b714daace6baddb4d43497c6c032d726d7ed1644ef5828bdd2e1fc8dfa212b6a26cdb7270be1ddc28359fde043ac7b0e1851363f8031e21c360c12f0d5849b1273f6e5e2aa69e6bac8e9834dc1a9b7ce433e9d2f7037e108c0698131fe8d48b8f5983e2a037ae8447fdded64914f9a0dc69e3256;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he595415f1e5d3413fdd18df0936b62c9cfdc869b408dbef87cd07998791489eb506d729a432d63f0630802546e23e965eaa4fa0e9798535ae13e4de971d43799d670c169c442c0177d1cfc0734eb29fd100909c190660ca38c715a699d6efd94832c4de47a36c2f2f70490b02f1ef02ca041c47ce9be2cef11b17b9d2d5860949f2950d86eaa477417b6aa1e84590ab710905d6639753e5a61900d5f592d5210eb8619971bba9e26dd7de9ff321162e040f38516794e7e27f4b7be736ef1e49834ba5226caf1f69790e8cd9eee5e8e39c1145ff974592182142732e2d73721ebcd42dab5cc9f21f36e49890dace69e230dfa3c24532d881479e56fb85bcf2f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4e55fd01b28f12f69295858c7d9bbe66a16d49ba76ecce312640eea918f2f1b215bea8e99a13b6442856af78f0d726e3b391c728667f4cefc3ad95268a226227c2d8ca89f294cc291c1f5dec8395f937a0c7774d8f7a2f9a4b4b6894fa090cc92ab9947c17ab9b2c6c8e12f29da024f613f0e4f3877b5193bf9584ea4ca5441094902b6cd64de79f5fd8d2a414d8f3e3c27daed657e8f0e42c8bc544c508014cb5391eb5f0ea4d437edb6efde8bc12829207d4f5a296ca225145454a7564e12158df6b73a8b0e146a5aa67b79b8504062ccfa6db86e825cb60f9d2bb1367524cfa8a0e644548e7553a43dbc54b6c11a220480b580a0a0046041568d0549cb25d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfb506255dcb4b321709f91343beb7048a1513d7e3e31ce3c397d9c5586480698e7b56023aa9ca54ac6b93de7f03dec309ec9e732c297158cdc5bd988e1fef0112a5e2f8752710191ae0c286ef227bb8a32508bd19ca0f88e015d58c1114803fff435e5f76c15fc4e21bb5bfe764429347ad51cdef889ef9cef588592f1ac0a956a3731b0bd07befa8afb6d3cfb967db350a84a3cfb49e8ccff081c019cbec3a0aebd6e80d8fbd51e4ffb57a3cc680bfc615f4d2f25d9d0a6968aed9b24a78c5be451efb8292179228a472c0fc432a8475acf5eaabcdea9106589496e9d4d0e154e36fc477d395884ef16a01349e389ebe26267a8b1c3a30bf33c2604b344e8df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he97bfe4ce9849d450025d2ff3872148be19df4156ef5b0fcbfd467d926e8574343fc034caa96c169e7d5ad783f36518f97f87cbde2e50927532a72c74a5260fb8c65a3a592038f5b2fd19bbd8635a00007df0df33df67a58df9358c463947cc60b921110683f63df5e3e4e9918ffe054a410c89ba723d57e05ef4d338ef4fc59951cf31ab2eaef023b685df53ec03946c245cde3380c809de3e8d7cac5fd1e7e51ddf63565c698f3de63e3a1d73ff944cb4c89eb5ad2b39eacadec1b7982da7211f01d8bde76d663ac28c11faeebaad858fc268b2d8a75fe78bff377dd753f75a75d8119ac739d00550ae72235e5d3d9967396db5a7300abcb66314817f1edaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h568deebbea64de662c47c37f97672b44be7e1823bd4a9cb2418f2fdd89bc2b5969ead894242b1a229f9b4b1578b2f3ddd687776a8b94f80fde2d099758213fe4bba18d1f818c927b3566f6110b8b5884b46b1b0867d3e9ddfee90a244c49a70c90b1e14883182965c025db6074b4541c34a12e264538eb1d2df4c35e7fcae1f704a788cf4fd0f3c0232ed8e80c900741ebe7f1962fa95f74c2e0abd208462b957cfe18a72fa5416fdfaedb480dd432e0940fe19a3412842c77c88302af3b8928c6144d3180ccf138998cc8ebaf76fd303a010fc0a54be7e7987d42704905190470eab326577d2f075b49368daf28dea98fa7ff02b83961d1c0f61e19200784a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he6b837bcbe628e91c848dac681283fe32ebb97a21b1bdd8398c23e580167afafa66125754db81bd155019542a8aa027c8db083a9595276a3df7c821b1e8f7fbf82cb14be6ace2756b16e99f71ea86a8ede1e0fa3a13199710c200670917ed88b32f7cbd63e569bf5e0e20c5071cf08a832aac3712dad7f66b0ed9cbcd1b2d74a9bc52b048033e0b66633c8877df07cef27bbb209d0de0dc6eabb9a2748dd55cb01c373f6f446ddf934f2edd8db33f5373ff9df895196367ee03422421885caaf324c02c2d52aab1765da8f212d1985d9160f565eb01d94056f447edb9347a47fcbba5569e30a1d4835f17e40f80545682a3334aa80252b1c17744633e05d46d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h15a2bf56bd26b3b8f38cdbf85b3ef28055586ca2af4add6ba98b829568e7da1bf00b83b65e8cb1099a1c131d1292b73da0f4b712a855a4768b4efead98256160ad2abe03927bb364761f294ab51ba2c06eb85887eea8f6935a44c15556c32fff7aa3bba6bb649d895258ac4e9bc4c1b752c7a0b8c4725a36f1b9992f56484a1c092461fe7d4fc4d266297dfd2dda334bd40ea13da075089f7287846b2c4d87c2a6be739aa5caff16f382fa8965b86bb4fb6eabb599c161914c36eb07fac9d2191af0658160101128a9283fb2db43ceb349f65f1d9d9c87a2c11ba7292b1763a70150d9d1e98eaec10c0b94fd3aac5a5eb7f6f79e77f17b849f284764bb1c7360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h480064afc62f465347eb2cc08f0a122c9b2909ba94139f3fb8b276ac4566a9e7ea85d72c3378d4bcdf3dabc0f1ea70961730a9ecf2d8c76e2325513d438978b4d57b094097b03637695410e2222644fcdebf2ad82926b05195c12b8b9231c232884bee054ef558711b49079bd67a661a8340011a38110db3575be67271c35cef8345178cd9be64ca344b1e951d4e69f6eb1309daf13f283369ebd6c68c975e02c8b3021806ee3c2ed7cc937ee3e8c8b228d0cc673498c73738b85d4c2567f46af2cf1b100f3aedad875624349510f2811237eaa955c77a68727f567a82d637dd7abe5d3a5c87e10ba6031ebf9fd7fec4e19fa54d57139d379c9ac4e421fa5602;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h63ebc701d07091f86197d573692a8bb0ac87abd16b6ef19e514eea556755d2d91ad34ebf853d476557c5e3f55376abfbc5ac19f63570a3fb39196524fa8790be4c518b03c910fa311a357cf5620bc04dd6e473a9351a9212a27e1bdd67bd586c882657420314b6ac6884939ee2fc4acc5d18bca8bb27c7d1238bb43a01ae476ffa5a03fd0e7a6972a30afc7b1ab594d29818592b04f8e9dff0e20adb2fb46063eeec3c1cd282e6b7b983046f321dbfb731b1e735a575e70e70013ae1a6154dcdeb17d91ed94ba44acc9558ce19bdefa91edd3ce40595a557aa123ff25080860b7655640f03655cb21b57097bc09efb840997c9152a3bd5fc6c3e161ca06d0968;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h486e33280685cffaf35309f15188a33c9b60911b843f147f98b857cdb7c221a8a4a04361b5bff433e00fadfaddf8090fd5aa1075207f8807e63d25b4c5cef25f9059a503baa4501168fb8674bc62bd00d65c764793c57ce8ebb6b5f25d1c46e12e4766ce17629388fd3a230fb0724b29e815faf406316646c2f65898af3b5999944e10fb15a780705b6091963f49e2edf6eb859f2d904156fe5ef72266d1bcf7bcad7779bbe17cc0271d3a5b5421bccf7a61def9134ec7fbfbd6530d622af02eb17c1fa27e865ba8c1285d3a906ba6653eb759563f393f31472e6f3b58426ca60bf8ac4919de8eeb4c8e4e33b254160af7b18c65f9d78d86ef73ec47cf366796;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hacb2771c55166ee50c4111d5cdf5781f7b2d38032c9a360bc8ff9ff1bc60e05fee113914a08dffeab4543176b4b26bddb57f8972a848c83f71d4379ee27d1a6231b0ce5de3b17ae7450beed81c954275203c551edd0b9b5b6413845ca159bc0a832d07e9040f438dc43c54fb8e8cfd512094fec9afb2deab4a14be5d8784d1a41d094c71fb86f0dcb295a1cc2a35977566c9470800c66566023274dbadd98fee162dea5deb7c6de581fa3074bf072266cee878eb9e2fa7db166542606d17efe7c390646148cda5eb8c5e3fba5f5c2de2c7d6295cfe9a3d17f41df14515b3f3cf4c893dc95d720e786d8fbef1132e5feff5a9c29edb16ae14ce71c1bc08d9d7ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hba9bcb4a0fec581c2560565593e281b3be13ded32dddfc78edc7263f7a515b5303ec644eb2e8b94598baf393f00befabd2798a14ab12fe2a1a6497cf88d1c358101190b5f1f491a38e0c3cf0e0891d5171cd6b5f7239e985e16b0570fe4fa5ef3a2bf84a798b385d2015a44005f6187ac2b4548a11dca447c872dbb3c821e32e1f50cf7eeb2e1144f6e166d551ac41a38e787b34bc3861592cd3bd97447c1346e4fffc2d13b863552d0b4fa7f4cfe3e86bcd634c29a26e2f3de245c56b0258528df3426297129a3f6dd733a905e02de287d0d8bfbd02618b1cd4eba163c0e3e30b8a14ba47342d0e1bf283658d44bd21c1dafbc45b6c5e7d93959917e433940f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h98bbab19fe3cb2d3e5150325abd1bf9dc11d50a2bf25f2bb3d1907f314a250d65e92db6ecb368b9f3aa395db85c0e3ee54bf1bdcc83c6ed2c59e78478a0db48eccf142691f46c2ec465eca362aee3ea6cbf427cb6cf0de3d61b9cd111cfaa0750b2b144c079971a7230323af51abfc5ea3fbb679119d2a7369c886bb6222365e2a4aceab12e60df95f0f7de74708806abd957ddec9b8cb6892cd0cb818f040f34c9f73d0d6b57507be50113db71cac8263ea25d3eb872a67d98c41d3bf2c4bdc6a15a44899000f9cfed09ecb38e309681796b8fe6594b0c105a0e155691dbd25fcdc633891c785717a6cc42d33dc8753a76862953c8384f9b1e214bc72f10292;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfe1ab4a66605fbd536aa29d90390f17d40dcfcf0bfdbe5d9f13e8a34050370c9530d9158ecc53d8af5e886399403b14798a0d01207152dae859020fc02dcda52657806d73831575846e195a9eddbcfdc423526fadee0f684f6eb7d1b28726e97fb4ef552dd8564cac75d441ce6567bb831b2f5bce94665a87dc34e54bd6b82b65754856f030ef9dd46f07783a0fac5e91e6b0c4d73fe46ac5910fcc77659f3c64a967dda4fb404e7fe6da4d95d002d5050ea70eebdd71ad90644733c26af04608dabc8da8632afdfb2d1f8c49ab4aad9b688d0302468c31320350a6c56b8d2c032acebc21a5087fd5853ab258df2f322cbc386779d7219c9a5396d696298b696;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha84438d06c5746123787f89f003b0824e98fdc1f799272fafc3396eb3ebb4fc1a2b7c36ad1afd6e5a907b1c5f68aa4a29c4d2246011a95a3da2b7d1a3482b7ae11d9ed800aa79fe9c60b9df9ce8c774fc359b6d31b96571947429d1c3f61cecaee1d05c1f6ad70d280845fed1aa5bf9adc4c66f9e7b06028ff09b338e6fc39604e329d677592247e44de0279b04ab37b7274704c249d97adcf38845bd5cadd1faf0733fab3091789c8e45cf57af92e5003882c90977f77523f40339ce95217b08189782836bb663897abe5cd48496630b0ecca62ee7a7e1a86a31cf6a407aba35f5a84df173ac950aa377b20ef0bbb1143bfc0511e6952ee91deae253f200e6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he5796d17ea62f5ceef87aac41f372af05ddea66ab762a908fbd50dc197711999629e2a6976dd21646f155e0bf88ba120c2041be51a59b10859092e1ac4b311d09f625c7a70ba8429df1aad1d1373356c05688403ebe1cea7997899fa2f9d04244ec5a4e19ed491ec41d89edec057d571b9b104639162e911cbeec477cc2294fc509974a89a762067cfef66a3b8bc998e99c96279e29cd5241371872a7ec202cb9883d80e35f5722122276f1be79e3ff4748ce0d5f5710c35d0050b689d0b8e13f0c766dc6f33e5ce964021e09ce106254b733c8504d3423b77bd90671853053441e61619f0c9dc233baee892f58b9a7975a381630df7dc4ee0de340139e29745;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hed6aa52142cdd66b05b15bf6708908d3af23be06fae88ab9e6e403c746f00be40f1f20b40021243a2e39605534b37ca9f7acd22846358c8f94608807bf83766d6f42c43d34882c1f01a93a7a457d8e3a812171ad2ce29160f57621b57c2c3e99ffdc5f00d79b7f4d7ab78333a93b454cba8b4a794174a5ade085cab2caf68e8f899a1756d57f55b0e593a7496c2c9e74b86d9d95d160319c2f7f58797a354c3ca3be30d6bd3789bf582badf35b6c154ee885f7ad900eba1bf04c5f5e78331f5452b95c6cb5e18b6bbfb9b8c9aad55ddf70fd0d5d38fd128910960620ad963096e4c626099c017b2a58d1c766b94698c436c9fedfee3cd49189b4c955669cc3c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h313a6a114e6e1a8c9f36cbda2090be62de18979f75ef88424d9dcacde363f1274a117f89697f77257ceab39f9fd33d91caf693688e88495291d7bb3f129526561aa059ea28a7663b8a2c7786b3ca1f495e22b443e527022929e8cf08cff63057be166ec341f83e85311e0e82c3618ea3a1f211344d49c2b81547b3bad2ffea9cdec2eb5a2f20e87b07d12273ac2a359e0dd084c922b7aca308c7f30b4141e18aeb7b749c036f73f4f69295837bd4524da122c32114eab37eab56fc98e57a20d80e76a9db5e458e8ad5c7dc39cad786f3af88b8b5221c52e1ddeafe32fa5f7ab39b7da73d21592ea0aeded0da2a30a4702f9f43d8a762b2d83bd6008917e95408;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5877d43113a04d5135d6d2fedb86effce8c293ffbae56a4f417cb55b71b2fca0af7a9a0514564125fc9260df733029d08e9ca222f0833f5db5cfad30ff38a77afebed858c6080340226377c78cf92810288f464978fd7630c55c4977941407e673fc6b7a1ac80cc6e01dc97278d0cf8e15890334abd49f4812e0ee73f7b30a7c377af79c45e82421b6e7e53d61eecf212bec000a6d149eececbf0fa786b49e193258ce7c7d87c8ada7bff74d03954c5ca02d5cdbe4c42365963865b41e40295de098eb7bd78cfa5cfb88be0ff8d8c59a1dcf41ef6dba14b7c5e27b0e719836b69ab72b4b3c54ec2969dda3b64911ab416be0d224e17074452108b720dccd462;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8aaebdeed84c78eb8e4549e2a503e2bd18beb9f19ee4c55b374430358ca32a0d71ce7b493321a806a20416389dedb90e82f8caff3ac7b6a8db4ed6a1b7fed2992cbf494ff4ec458370e96a58546f3a8fd6e3bbc54a581a408334175e7033ef9abbd12ded6bacced10e1d834488a21af2b410fe3f016aaa7153c02c6a6deb69a30cdb5af8b5bbbd2fe237e605fd71a3ebf22a1695c62e973e9bef29f93564080ee78a08ec57e49b5ea39dd443c0bb566ba98cafbf37b5bca5900041db43ed7c169372a8036b5dea1ed92da460c25f8b92c5a99f9b21189adb8f465ef0a6f0c2c0a31b9894ec03cceb052cf0f08fcc52b4311285507f43ca372d1c78d64a50e126;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfd62a37a3159f0361da28a9e549aa61f5194af231ad768ab9d857046a48460e5024432343cd066efab157f3dfb09e9c44f7d48d114c70939c542c99f233b993aff66dee616baf10bb86369f73ee5f97169eecd33904d5a7d5cd09d0f94659e8c9d8bd1905743b0980e72eb26686b1ee01f3604dd5c6e084072facdbddcc4e59869e2530ec497b122720e57697963c8faf3942943c37f4888c481b2479f150d23279fb4598b66c0d129ede262470bae75dc24105f2bebc3b6af1dde0d7c146bc4eaac1599d9827bd7479db7d549be5d8beec887f1d3e697e7426a313cbebf4fde5ae589ad07f27ae5d4d548d91d20be0a5d6d3bbfda567b57cb289d7489f7f5f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h18d33eaea05f343b5c587e3f520f58630698566a147d7cbf79dc1c81112f9e77fc88544afe350920744da514e470225d62d539cdbfa0804a53269830f62fb09c133dbcb4a97ca4cd3dcb2528948e30dd8bfa5db0a01fd0e44f4ee72d86e3c744a37782b11b93257607b5f1185b18c1350c785d667dfd4355897cc7f69887bbbdc57323dfdf9f5f25d7512b520fa95f05de75b81d2dc17a8e3a3bad994be341341a653cd6e6e99b47cc23f069ecf85b2353c5af9c40ae4661331b428f9bc443ca4f73dc4a0e9c9edac1b8947e6c561842eba034d95bbc9dd1cfb6552b93b7f7406bc335a228b550751f2da9a015b4dfb4b21d5ce42da346f07bf810a37546c41e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h751e4a579b83d4a36d9bdf9d31e6844f9fed09e4a5c1d42235e955f9f22f08979aca85a72bdc431fb2e30d31b2b02a6f9c5417649e05236e08347ced9b31726748aff3c27199c4bb5fa65678f19628923a7e1bee9baa20084b9c22abcf348c7c0f33afa2ec66bf834ce4e64ef1c30eae15ced69c904a6ab9567c4ac75c7d17d536e9c9838f2a38da1122f38f174eb866f26a1d5aab40ca1cf601be594b2dffcc48c1126d06cff9acab0f03b46e998f772df7f2c8c9784690f059045b819fc130df70d8436ca0b238b1ef3d96d23b33cff2fd1896d5cdab2c87091fa0254f726429d769960b2d172e7aa6d80b432913b5336e09182106de30c0c0b051cebad0e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9c68aba3b75ab77acc024c32b0ad0f8b5913f70c64e42c7c0dc9a8322bfe9a6396d468632307ea05458eb02d0189135686ca569cf5bf72cb20a81aa54545cdce300e9b7ed0e828de4249e7a95b8725f63a960176844f5f7797b7f8e0bc373bd69cf1c40bce5a0547a7bf1e5c87f1d8bf1337c8ea5f2ebeb8c28f47434b5b0917501516ff7798dec610fe4e11c372d10ecd9a18bd699182812a2c4e84cfd16318a6bb4be0f5b2f600d8f3d5948ddb8ebcc8aa2d9aa05d52563cf3ef4c4986840dd660e16d280d0c79e678f5fe78e6947b6345aed7e81de02dc49d793277a54f84c2f0d7064f697f30568ebd4d1246945b1afaa08f63a738f358850697319d792d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8668a70a5035c40302182916799dea779cbbdeb91dfe6fb0c052dc7d8dc9ab4e2d57812342cd9eb1978f4ef7321d0dc3373e6e493ae4b03165959f5a82572e8e3e55fcea91794b52fc358d439104c77d68e69f7c433e103f72773dcc82ccef8f08223eed8168600e32c731a491ee99f7431525e99b09ed072ad42a923f7aab8f2e1eae0e7237d858410bb726839b9ceaf0042dfec1a63080eefbcdd6acc5cfa052b415f630e86744772ea97301dfcbfc82403c6c865664ce05b410b09b11c4877ee24d1f074184dc37c7d8d11f76c7eed95ace45d3a770b771f88f2c3e2e69164dc4f260a69dd90a96a9085fa3f506f46f0b3a63c9a2b334e5d9ce547827f32b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb04f7bc9985d4b9a813b4746ff84e719f6389389d8ec34e1a9cc4ebd63fef0961107e9c0305f00d1a5f32e2ee17f5086d8cc60ce4b8625365b4c5019c19d068f863a297c635b55bd9910c095a9cf3685a67db7849b9aa67928d322e636ec6354873e4d8f28aed1b674e53fd01e7064c6324ee35c528188e0d46f78793cbc4ff5ed1138a476ecad22e3b885ac2e9b0d32f02ecbc66301612b8dc39031f26d07996e0ecd51156fb9a9f3823d0ccb394b230c2ef0f97c71c4622216be2acabbeb27b3200fc5431b39c82f18fad6d65a1adc1cf175484121b5a32573520db32a550a43302965f2b9d37b392cd88fee0c305998893788f4ae8ecf84749650e898b2cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hae1a1ba3a9c279e6fa762c97f5848deb435ce853a8e6f4f8c2977757d910d93204147871bb551589e2c9be05a63e27c50e891ba1bb4c4d2124daa2bf101fc9e280b3207383b6a0f36e4bf2cae1c92bf39d5e41dc63f1759479300a768f9ec74b779c8486ccfe163d837b5d4d99f565f0a8a78c9e35130585007c694d68d578b81bd0f327ba4bcf9ef3695d24fb4158d6e5803f7fe9690cf2dafd783e05f87ac8787907371e1da5c2eb164bc72a064513fc8d27100fc91af8e89f0a6a16907db997b87be596d78c6f29d34f178a95f8624f0a953626e3d413c2ef238ba5441aeedd5087c59b0ca9708c3de3c50d6cb2d44dbf02613833cfed3de0e2c0acdbb9c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7622e71a107b56e9a45181d1fc45fafa63eca1564831d788effc726334bbb7d45632a2f2906c811e6324c2fb39dabbc3cee2b9666476c58a594152f0f6b65f58f36c30bf1e438b21c1a83609741fb823b82e5445d5c5da92f8184fe55a607988279e757ecdf46bde98985e42263e4849bb208e7d53e6014d5f8d8c3775a93525ca9af3d04b306670bdead050cbc97d3d350b0b60c021fd8bb7f1563cf358d5b298f31a569a0b013cdf5588708873e33d0ef3f503bee92710ed839723ef0fd7fa4514e490a22e851296d89151fadf52a716d0a2e73ae1a90675d087a3659612ea792c4acce757fd1519e72795a1fa65f4fa03d5d34fd213279f43c17044d4c264;
        #1
        $finish();
    end
endmodule
