module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1100e81b88d979916b383;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h430ca8dcb043cb524089;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b917f7af61de6c41c00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb171858fa33eaf410f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b3217241e5d9226e238;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff96d8724e00489dcd35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1893d3a7a3a58cd4d18d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heddf9f15e10cd93527ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160183e7badab4a12ee56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fde7c3b9e2d676e2d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c90261400d6a6c30520;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e91e0f76cdda29a73a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19298526bb0d664a24ec9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173b72fccdbd9a591da28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h618e28e6fbcaeaa97a11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2e516a6ff33d951d980;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c1376cb70e5d22d1e9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf31915d63406f1a366d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15187184f6e789c6b2a79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he19834d6620f634c174b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0c1cefc2894ddd06577;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124fc625603ca0c1cd020;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf21c713ef07c61b7fc2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112db3ac1fc6223f52dff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2104af94f2a71e2b88a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f42befaf6556b319a75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e8e63d2c2a19de06b13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148534cdd65498e958dc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11bf611b5a81cb78bb44f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e658e5b99bdc6d2de3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b5beb46c92c9429e36c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb588059b66196f255151;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d280dc4e0d27516a875;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6767263bcca62af47e59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ede1fbf96a34083e97c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcbb8a874c2422f765698;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11173df25b75e7ca9811b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1587841f13c52e7d96e34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d3e9917522e09476103;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f10729550fef9d90c71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ab393f1e6432de2b84c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hecd0ace1970e3a5cf4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133e41555c0de704c68d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7d0835beb39ffb2b9be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a38302ff5ee73e745a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f558efeb1051e48682c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1742d496cbab5a497ab3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16848d98641f079820ce4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2eb9b2e538c82fb2956;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a370e9cdf9b3a80f1179;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5b9a5d45b3c4f6f4770;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47f99251f502302d1ce9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17250ac461284bdda1d50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec3065402f6e656cf93e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1b5df0b01bb4191e062;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14850b8e9ad01a1bd2fd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cc4e7b4074655932ac1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12523c09b026d4fc25daa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b5fc636cbf8fa94a135;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4697e10f2ab9024cae9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26b890eff6a8236f0b53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a62b05aae5b8de76d83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a9a3282b560cfb94892;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hace45f8bde044d9a784c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3aeec5762fdf21c95140;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8541db222755beeacc3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14bd2af5501ec1b79a79e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a790ee8f112f49f0f7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h971adecb8bed97a00253;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf8e9c5ee246d9dd9c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7282b08dd4cca8304da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c824a6efa8645cc303b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e871814f17c7dd7feb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50cae953a85934e4abd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf00345f6b1f0e308c1e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41b70170935c1fd07198;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc62137249b50799f4472;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b166f857e9200c9bf321;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fd7d77b58cac7f56d6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148d4e8dd732580c02eac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa041ab63f7b1b19ddb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164fbd291e85b9c6251c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1150b6d98ad36c8fa4485;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d1e70b7b5157adc3946;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ca2c7f64afe8340d55e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6e7fb224975440d2a89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha357e7bbe5c21f9f52de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0c5b2659a8fa27ae42e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf39d3ed8f1542bb35076;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc7f01159e188b94cd5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee2b2b3effa28e9f6864;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1439a780ac29fe84c3409;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf7bb8c421c159f6c7e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f93e8e3c9c566c19f799;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ef42de7bb54fc508550;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9fbaf14f490d0cd0669d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hada34b3f794a8cf30e0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1736f40f1659d62c5e3d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112e1def9a127d90fe668;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e0783ca328c78e682a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea44ca695dbb9d6f9ce7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h577c53ba7d69ceb6352c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae0fa84bac6cdf55f6b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147056b86b17e086c1c5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddbd200bb5cb9a902a8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b01789d49725b4356d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f11cc15572d0323eb327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b34d0e3852784a14766;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172784e3c1eb2dfcb70b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1992dcd342e8984bb6016;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h980771de6847a6c64165;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cb51984f3ea2862c83b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173a0033d79c3a5cfb9d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10722f06649f0db68500;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15481f780c0e9d5c1ee9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1745b5fd709e70c489710;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44fb7949387461d3f0f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17880ece4417f7920cc4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157358b7f86f84d024b2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8eadf002f08f5d104cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbeeab15c9b759f61a9eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d0b4bba73b7e01f32c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a547a442824566e7418;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9df409e0d81287dc498;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe8bf16223bec26ec995;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae8f734ef63ccf4aaf3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39f11562adc96887dd1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f537dc312c8695c67add;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3d45ee1f89f3ceb7f80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha21ca8db0bf0f93ac7aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7aa81fc412f602d6319;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10672ca459e78227de58f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49a342f8ebc4fab2b709;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d98f04ce3c8283a6ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88544c2dba76baf5fad6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf57b125a74079d552ece;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147687e4f39a8999c5aef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9875ca0b7f5f69757cb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7f6482bf8831b52f57c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105b2e17913a02b143a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9672a68362b5e27665e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa6d38f26d52765676b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d9f86b07bda74d68c25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f0bf9c1543cd63c7883;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0caaef25a40009402c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5634e400b002387224f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf87012abba1e6ef9cfa9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1810c6748e1fe01a37377;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b7ce97ff2be4f7dbec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1426c719c16f64a608e8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ff53e30d293287f542e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1313ed91470eb153da662;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5841e8ebf6c631c524f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0285b918cc6359eaa1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1699afedc290aecee8afd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bf2c1b384690950bf03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ac1e30b9d1b0e273ad4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17892f5457ce789073cd5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d83dfbf884165ea0ee5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95688ebb2f68b8e481e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83914f0417dec14d9510;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1137b874914039a5b5f95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he85b06af285b42e2bb54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c29ea0529fa12d37b4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11974abe3f72426d3776c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4aac9b2a4e33fea0042;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f883f292ca67febc8fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3299efafc07133e9e9b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8221822e353ffbb51fc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ce350054c015be8d3ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16db1eecf591e056c8a47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e87d70560f3d59386dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h926a1b7790cf26f68c20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d5f47b23134f8418558;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc868a09f11610bc40a00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde5d35fe178f5659d428;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d81a6d8c2db1d97a1677;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b0ed11b9572563f15dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8084833e25aff1bb6b04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf8a17434c3df3037ac7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7bd96a1af6d32a28a0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b19b2c98b7e0a04a635e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h46203a56933ee0fe79f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc4ddd42f4c10ba77cd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140eb9addcdfb22e5749;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e4256b5002cc963ab6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4353a5f5a168c79eb031;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd716b7d8838a93de8a2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11dab1787a3ec72f15287;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194f98c6e1bcfe600dce8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5099bbb965d43f77ec34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b44da3e9d9963362e83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f8e67fb3ba7f42251af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55da718fbbc686206971;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ef8017716af4044739a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd87202b354e8254892bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158d100343d5a8a87eff2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbdd20788b706385db59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53dd5a3d5bcfc6da54ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb8ad1b06fec597ac632;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c0cef0b7e40c3e3fa8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11036ebe7c8d8a6f5eb65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11346807acf304cc47727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31558fb3ee3689b70aa5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fcda47396bfa2cb0760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1633537227bf8e85e7a86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h438e614154e47fd5ba47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c628e7937c27a6b65d54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8e57c82452dd1550ec8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26761f86b2365cd32a10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d4a710b6a3cfaa31267;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b5961674116b4176f2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88ef52004c427895c94d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133f4aa6c09c2b786d97c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefdd4b61c9fbc610d72e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1544f6be442960324f932;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1624f0208344db9386a09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h357b1094ee4b3eea0179;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94d01e5a9da7df435e78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he841bef501d5ad36c99c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd86d26241e5be0b37024;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a68d795dce3a374774a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he54b11212088eeb92074;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he19fab916074d23f9172;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140ae266a7447da46e440;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b384991d7647ade0b1d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88febd74df754e163199;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ee572c91b1fd6858789;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197bb4e4a578d185e9f27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98833f0b3fedad4fe3f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h980c739b13dd62275936;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116e7d7bcbb107b91d1f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc698636bed4002d94d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1089864b88add912c8b41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da5c7336a8285836d5ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184359f9bfbecaebdfe18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175e67f4d19ff1cdc25a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6b80d047b4ea7644288;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f3e8241aeadb540848e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6ffe0062249a25ee689;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc923504d86a1b1e8f476;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe59f18bdc6a7c84d4c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35269ac7a298b73547ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a6e04a9c74f06eb5beb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7168ff978c72763f474;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d9604ef59e7f5446fa8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f2398d53609600bbf0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16205a4cd4b11212aaa82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51d653fc575157376b7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141a44a60f0d5efddf47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c037feb200c330ab456a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176d17a5b1deffe4932aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5de9150c601eca267726;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0f250f2a116d2de1ecc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2cd1061b38b91ff0899;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a03419a7bbe2f90c7d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0c0094ad51dc4b24df2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff678d94e1977bc586de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ab26c5c98bbfbe16fb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf770a496fedc1e690717;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h864673ff1d0e56da88ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1adaff55ea615989596;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c49466fe4fc8424d826;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2c3b452d3800a8d51a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32740803acee2fa55834;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc843faf09aaa33c1e699;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb07205743d3ee8cabd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c94e91acc25bb27d8254;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe4df4fe4f5bf368796;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h381bb2c692745c82e951;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e7eaefbe489165c380c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd36b65e14d9c3b4b3d9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ad651e8c234f87c3d2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dff21eb052aa31f1f2d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8c388dd73fd6fe04904;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he925138e40e8c1d3cc6c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8dc7d8097d738398e335;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f63774f80e5580d100;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14605b3acbb86ae78c56b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hece04e7f56cf73c2f2d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8cc225b5184f2cf65e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5bfc0121c4bfe66ea09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1671ef0d9ab38de102d3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e1e81fd6b1f5e0b4e0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbec97b646cc6bd426808;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1253b69b45a6fd929d536;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15973eb6b3524810ce0c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8a68f0a241207f036c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54dce486876e3595db1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c02420cc225bfb3e61e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e5c43d2d5482bea15cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3bfbcc0573b233c055c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16da84b58e0343779788f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111a303cb5fcc0b243c97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd13685b243f91fd4b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151fdda5f3280a8f34bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9e41daadb138ff5a5b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba75e9e7c7b3469e345e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2b5da0dd9e7cbb629be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1700375b3f37d933daf1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb69cc568fb661ba585fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7884792a376f36081f7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189ff78015635c4d4c07f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188561bc0d389020d6035;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d33a07e7170e3adfdfb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116d7f94195a536f5db3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he51fbcbc73ef9c93686f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1577d183cd941f2e3d0ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ac087b7cd59f32ed3da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h814e55127405c22e6372;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c3af0706013251ad2c72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e46abc0745767ba757d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88c9dcaac30b9864f301;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a73c89eecd283fe05f53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2f30b51daac0104bbb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f491aa140154a8d4d2ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11558431ef44cc64ed7aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb10ac99caf6b5fb462d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he845e28f5a5eec4fce82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d3dce669db4d0edd56d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1985533028753a584d260;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ab19bfaf362636182c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb01bbe55569465f53d1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1698ae6ccf9b19fb7351e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135543a793e9352bb9f41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95ac62f0ea60f94a8cf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1789c9fd1d149ecc74dfe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1400ee0fd203cdb2fb136;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f819b602066b100ffd8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81cf6596a32222c6f11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104d71a37f105d7c097a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb5a29575a41d94225f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9636bab4135547a7f539;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ccffd23d659abd6d096;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179d4d5fabbf1b095e3a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heabda602a7c35457b528;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddf26bdb493535758712;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b31da1d72d47f42c466;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1362f0495e94eb7fbed4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10faf30748c6cf4c6b6cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c7f0f8b45a588580d16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d810b4e77735df8c33d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5447915137463324aa1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b610be87bca9ae7a0f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1974c4a46af94bb4f4c01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52b7c3e296483f9efe8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3905c591f13bc8b44d6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54865fb797bf1b0a72ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59cf9e4a35d1a8940972;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1083eb49e0dce30643e61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ecadaad1a10f73d52ae3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fbafeb81bcc2c96d0b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4d00d941230483ddb77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1587eee9648ff85e32571;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9977fbdb5c1bbe31584;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bf8ce26619b3d5487fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b4c803be2826dfede2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1691b9e089e1e4b304fc6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4015b60b6ef10e6fb0b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd6d89bde7de8ccda78e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe141b217b4bd4ddc583;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadbf8d507e65d445f2a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16582d93b02491f669b8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b1f8fac1732c425be63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196682433c7685a60c740;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fae4d609c2e08e48614;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38e649250e021fb5e04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc91a5fbf583f6605272;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b76d7f8ce5b451af5dd2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd76c6801d43760e9929e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d46970fdda604d191fa7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188e10b264267830777b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4510eccc8d1205c5542;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4835faed713e2768983c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d30ec9c4ba65881cdff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3512f391ba7e9c4effb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167037d1b970682632adc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17349db1877a5f145ba39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19779ba44794e324f399;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1b34a53b8d8d722fc6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7e3c188d24421cfde17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1e552691da1201c005;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha541ea1afb2ad91942cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd5de2fa6229eb4069fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9e803c65308572b7fc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h871fb0db39c5fc366a7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4f4b2800f7b3d04c67b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1534e35f665fd4a36c232;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb55c6847533c8f7bee09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e39df39b7116c1dba88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e108f8413cec7fc9594;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13837b98836dbba0e6098;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee4fa3432a87c672bf76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d377c2263e43b3dbb930;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc0fde3ecf64abac5878;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea716a06902bd502e7f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154e743c56ef7d6b1e1a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3820fa93e7168d37a28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf44eb76314288feddaf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30696ca92fd2f8325d79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114209fa77082061878cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1fd97a3922ded098f79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84e7f481d742e1980011;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h710e54352cb1c88d34ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfb66b5a79e70baba6d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1196c1fb53f065abe0ee7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68dec13f1982f1913a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100516675166338af39ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1413ae2b26b00954295d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5deb5a7b91cc79785724;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8de5dd3b8b1318312423;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc25301e43759edca2448;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe2150b3b63c0110c52c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1144692569323ef6fadfb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13eb79ce3afc9a369b480;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18dd55816d2bbdaf3f7f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h333531ee2f3e77fd3e1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edf2a4fef23361cd0c0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8155a450d310517e1365;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2482917f122ded3a8e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18878053dc233c7ca3203;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h979098cf731b2017905;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7da62cfb4bd595de8524;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191395367e437517b1e61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9c2e20bc4a6cef763c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145cc78bda525c34923c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61c2a5d00f6455622d46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7a750e5d994d78cfc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4be85e2445010ab528b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11dd6d7e32aecb21ba0ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b5ba149182ab0dfa50e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf6cb079808ba1269489;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6ac8ab551052b0d12e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78636f881799da2687c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119ee10bdc75330dc7a46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c4d517a93661e89fa2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed83d18249456273d1d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1375a5a13443271a5661c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c1e938e738496aa97b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1761f23b95ed80beeb2bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c9678f259b36e0b0c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9b2b29925d6718d0258;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff89608efb6737646080;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc67bcfefffe5c2fa1b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9f5aca60089375dcedc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9939db6dbb1cd5c19e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be03826e4d2540b9cd99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d59e49d4cc5f9e8cfef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a658ed4af568be633ed9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f9007b07ebb15197086;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21993e5413cdfd1bfa3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdb45030eb31ee640828;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1366f168c7c30c10cbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115ae6ba9ae8a747245ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfddf5efb87c5c8e200c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc06fb7c0cc644b7cd83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0d7b76913e6d9ddff81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1230927af37b3772d245b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ee84be8d629d3173f5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e5439df9415f4f161da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ed15251d878b066f584;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf340f77555b4e15a29d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14409fc282a7d7e9b9d57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e5f17b0364cb98876b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c03f94316c6670e1bd21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h686f2d19d8a07b46f948;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7acf2b433bdbe7d0073;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc6f1c1e9f8a5ead63f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dcfa94c7bf884d16679;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a8f8399be1fd124e162;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e19353c6fede22a8adc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1827c864b12d4495c86c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178c68b1c60610ba19f6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67a2d6238369b84dff87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea2b2bb7eeb18238b80b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h201d2f69cd412f3aeab0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4685a895943f756af1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d789a8f4184df698be7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65c5c2d7638dbea13703;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec3be049845b48a74680;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1326a8195c0c1802dd329;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1fad804708dcabcbdc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf11517eaefff28cff8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a957a45947f6c1b0c55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h589fbb5aea98c2a16b74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h767683db6fd930ed7576;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc539e34559c6014ef589;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199a015f7b582e100ac89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c182eeef0871dd62f85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3843bb90162cdf5b054a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e05fe22644d869e8d58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa61256cebe99cc0a354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1bfc9f80c19e5fb7503;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2da26baa7a3d5d6b5e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afdfd1fcba20a26eaafa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd8e6b7e412803b81f91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5027663313f5308684aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1426d8f68eed97cca47e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36f4e2e5fb78e1acbefc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10bc64401041d9b24343;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d4238e89be2f65de159;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hacbb31aeeb0d2ea1cc60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he055fb4ffb3311362cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h216bd806f1be4d375507;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124a53c17d95c1d29c4f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf4c4b2bfe4f6671613d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a4e8efa5065aae0a2e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d190973adbc798af19fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f56a25902ca91e7511c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f91db45edb0dbe3b3dc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c61963b2faa17a01430f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac4e32295b39b9c78d4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1235520256f9456e82147;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ec8746cf5d412f4cb4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a14c3e621aa596d0b6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bd277911d7387777a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c307ec8cec4dd841b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115204503aeaa261f6e32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a935177a4970b0f9a48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1accf5d9044312d2122ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cdb213c46ee32c7749d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc50d2bfca6923622799;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307e784ef1fec2f06564;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had7fa0f3d398c3377bd4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb59a004a8c6f2b73ecc9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1155293c154bbf1f48c70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70f2713dedaccb98e411;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0208e9d4e161223a27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22418c20a7c454736006;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4bcd6ee6d489a55db12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdf6bff26eb2ccfbc8a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158261af211525ba9266e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf33a825fba2260306e15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1119a41a51c70548e6a5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h458303539d246cf950cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16881cbaf0cd2eed49bcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b32e7c7508329642e91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdca6d3bedfc75cdb88bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6097cbc30ed6f18e77c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be4f429288c503d8d4ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd23a6ba469c82606693;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8793a4a552d149f45a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121e860a21797f07a375c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51ce435c361d897a2fff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f275ee12d74cfd287be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dea3c55a6428f438fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca69304ec12c0c0bf677;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d401a97c0c0710495314;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ed421a3abbfd0163183;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9bda5d4bf9700285afc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he313b3c0eeace18951d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3abffe009103b7bd5721;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1025bba39d0a62ed19083;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6f059cc62046d72a89d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h601d2b930b54df0a543a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f2baa78c7a8c69e424a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h768a0066583dbbfd530c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1915588235a2d28adf30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfebf26e8201a81386d68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1471f6ecaea8f8c35a940;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138e00e452804109d5a3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb23e9a8a017b644124e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf75dc8d0a4d7380a22fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d75831004fd4c194be96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18992c36ed8925ddc4628;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hacd1f14f89442c04d821;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8fae5e430a2c15b0e16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d08043b28376017330d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15983584f5e865a39c101;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d46e0962b589112b96e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb8e8363fa885e1e386e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a63ed6ce04f0326ee5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24329ee134a305f47e32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1c9597625b18f406433;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5e14ecc29839f7e5b27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e898c87e88367c5ae4bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h91a88b10124f9b995046;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9c305e31ee2902deeeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18dcd0274fcf82e4cdabd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb967f8fe2d3387753e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4ba75640621ee9a61a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e6ab6e6032d2408da30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f819f54e4875d6994b28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fca48889fb5b0b7270;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d333631ad4849c5bf2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f61eb829ab9fb4c58793;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11253ed65763d043d221a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60a15b45671e6bceddb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176e1d2d36f7e9ee0f07b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec6baadf48bae70c7d2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b9ef4a6dde25e39982d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5568af4f9a442bf2153;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc068ae94fae85033f1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22f9189d4e5695c276c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b81d2e57a4f6fe7b757;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd43d8b18b7ba51455c10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9a346277534d404cd9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ee57d15a56c1ac0a221;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1158f48764a3d1279fe47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h77e82a93b619242d6a96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9a078718bc0240eb969;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142de05c0daf1f9e3f941;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0bdd8e9ae05699a027f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hecc2c39f3c0637817ea7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d13263d064c8cde49e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181ea1b2db86d6a80b1b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe8b0f7748a64b40cadd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf971f401e516c643219;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2bcdb185e4ea225681a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da91326f2c25dd20191e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1942afe3973a1b227cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b7fea4e1c608dc858d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f540bb039592830e99d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1345bafc9f7e9f150e533;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fdfe9c5a419d7904d3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11cc6e47342a8d5ec20ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'head1424daa68f7bca18e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5209fc22988e9f72c7ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc9d80a274dc2a806690;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ed30c9f0797ea30c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h122aba7d53c2069f71a88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d725217e87a5525f004c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f80a6cb3cee655430c0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e4b78c07f44fb00e073;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d059f6eef903345f134;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16143eea42a88166009e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99fc83afcea0285d8249;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1819db25109e7c38f9444;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5475657b7a491542d20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h402c35c9d04f0d3c04df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182cdb38903469add8c92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfcfc2e4d53387242e250;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be1346246d99c9e48e99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfc5d90360e015ab34c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1425afe24bf1d987f28dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab5e7bd56ccfa577358c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f77e102bbfa2a8c47436;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha97ef2686c12149f54ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2196b55e78e319285562;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d663152f39d20980cb90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h316b030467f5fe4c1b07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha318dc653224c1525668;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e61eab529472ceb77b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f93bc96acb65ad78cca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131267f5671f0f7c058eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ba8cb7f6b6696006892;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cebdbfbd3bdd51094ffa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ed515d2520b5bb89815;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb4023a4eed83e904a21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d28179401ab30505809;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f79bd40a928fd6a4d90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd90b84ee52d390c4d59e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14af0eba50448fb9f717a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce3f868a5c848473dc71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13eb35426ce3db8bdfa39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8e309803587d531f2e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0c25554f38930942ef9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6cb1f19f2750cdc0dcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5591349a6562e7fec13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bd5aa83b0619b5c7f1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda95c3d293e1813ff07f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9668846e57f5b8d8af6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9318b39e90f7b8f50eaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0855167440dfe8fe43f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16953d0278b055633bfb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfae1303ff99b5dfffe58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1decda1559f5f69df8076;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf59025fbe42ad8546549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83d43c066e68d3d8143e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191622980949fbfa60305;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af9f9c9f4fc5bfaa5218;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198e2f17b522b3d3d7ec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb9eca2534b9d68c78ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he676b26e5815b372dc49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ea715fd0b9f9290959b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfab65c3062f0ac3ca71d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187826549d8227736fff3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afab0ce2679f42253e80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90a2e391c2015e66b3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca7bfd5b0d470c558c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111fa9c2c47b6ffdef848;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed0868da640a9727ed9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf77cd07e71c53ae1632a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc318327463939c3de85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9792e6db9c33f0d1640;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1996ddcb2a15bb2d01494;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbe9a3ac2b89b4c75b88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bfe8289afddfafedc46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc72754b7f51150a1ef50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb333853edc72f1e2548;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a5c6339139c8d0811d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2f65244f03ced4b2b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40315cc2b44022b95689;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92980375d28938e9fb8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2430586c6efcc24eb5c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1284005e69877026c1df1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h311b6781bd0def65adc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3373abda02cec664a009;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68dab5a7c13753fb703c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186563c97aa2c8d203fa1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d52e205bb972902202e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d29426a63410830dcb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae6d1a9e638320997558;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17cdbb22fd32e45a94179;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15147b00126d550e7badf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1982abf1ee968d91eaea6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf6c407a7333984ed00a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1769b0a5db2d00544e053;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134dca0fcc5a7422f3903;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125f27160b60fdf28702b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199032fc4c8a89dac45db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7f1b1db15bef4bce73f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165b6e3d82352e02995a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfedc648b34e225545ee5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcff25c69ec9dd33a105f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102ee54c6fbe7f76d0bd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ddf4d456eb1e67902d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1345ae0b07bb0d7be48c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfb49be38a1119a8f69a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0c089cc16e2202921d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca66923b3264cbccbe48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1402fc2deec73fa581012;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha15a11081931b15636fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c0bfee32277b6ed7f0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8279d28597113f06f2df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b116cc93280da5fb7981;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14360ed226c7454c11b87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f38d1a930b00d6886e01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7adee567930d06806186;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5b8216cd2289ead4145;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc272d79dbb2f4ba49efd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b587a5c099f752a00d64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa570563c7976e41dce9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f157f90c624bbd7e0489;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c6f58773a7239598aeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f27389fb266afaac1893;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16003e24409bde60c526c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h482f870a40b83f8d5f66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0ac8e8ab10f5133847a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0e0e84c676fc21ca6aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12982c6306270dac271d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15157b1bbd9028a737652;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcbbda8f93b0286757ec3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8a0f6120ba41a8a8c50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198ac7e5d07a18643e7c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9f52d6f831551b3a946;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11fead743204a5daf022;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h418b917516995f7460dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1e55b16b757d7256d08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b03d0ca267077850e73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1bcd97f2e1e4545db49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdcef79bdf90257278ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96da14ec80b0b80c01b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc565a3141096f14eda44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197ee2201f63b143371c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8f40e3327808912364d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187435aef8a2c4f08a0d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb7a4578a0852810322b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4307b1f000a8ca577fae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191f71f7fccb18a0d022f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a7566b3885e8e540a2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4cf021ff045342b69ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bbcf0039da180831cfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0c3743e2c5603ec4487;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9778730c7428add98578;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff8390b4ff7dbdd60896;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1e5f41de03bb0f6a48b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148b0c599639e73785b10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1102a9f3b6bca96212116;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb6a4242ea2d94a74d61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h91cc98b25b171cd71915;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbcb4548460ad65a1720;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb1307c6cc7d34adf37b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e532d798acbc134886f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2e6e90e324a28efc6fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7ca73d2ce0e347fee4b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51d0cf5bc6aecf715313;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c124b3ac282dffc4e5e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e2b16cb85aecfa9773e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6af9e1141a423ecc1e94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h574966988895d41f0242;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191618e47eee8e8df7cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c2271c4395b072b85af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7330be860fc11e1b6b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4748752bc84495999e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8e9d9eae8d9fd9f3087;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7b8bd62d969f909653f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he56f847b1cd4d59d8f37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19da8bd1c9c4f609ba1d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15169848c60d363f2c09d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5e22560960e15b582f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146de46356a18bfd71001;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd27775e244fd1faf133;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ec3df2d3388ebe1b3d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c54184fa446cf64a6a19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ff308b6ac9dd9e9836a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c308dd918b01451280a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1582a9fe566e9bf35bba5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14642099cc3647174d1a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae84d98404ff76359e22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1951d7c8130f6b004de6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1fcb1b00f01897debdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5bf604848e90ceaf5fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f33b461b8c6d7867d835;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125b3cebd7f353d4a7134;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1053a89862ba1271f7d87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbc7b2a5f34a8e4b2e2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d1dea007a7f790ea0a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1007962b962eaf8292991;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9315fe73e920ff6a196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a7cbe17f86520089bbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124f95d9d90cc31444281;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b8004c23b5cadac137ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb98aa75b76954291f03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd0e3dfddf24c30b5af2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70b02334287d8a1ce591;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4cdef81b5d321c23f19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbef7f7635fffe830e27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24cd7c7e36fd20747cdf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1001acd8722be0ca84552;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heed37bed4a55213782ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a53ad7f2d148f8be736;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ccc5254b4600b31c26a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedac2a82126b8bd99ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h77ceb2af02580754cf11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159cb237cc2de27c0416;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a59f2312a552f5f5f067;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b0fde53ebc71a33236b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbac6e40fe8a1b5298a5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1641623e41c86b71cd690;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170bfa8c63c2e7ef52755;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cf3ce5e6017497d60a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b8c8259a70e4ca62b0a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa4217537c8e1d9e4d45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ecf5a31f819b65a7290;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125397a1cfa8309c18972;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee9457d8ee6d01d8f4ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfa049465d0b67e5ba42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1857bb1500ac28499edae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f65ec052603b12446fa1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4de107acd0c23653750d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c4af4f14319b3be91a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12861735b48f7d1345516;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1716d8500ded0e05a26cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a0468a29620c6fc8261;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he716e77d1844883c41fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b84e62db94d51e90497;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be734c60b1c5c8287159;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f366724d95908e74e0d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9bc751d63d44c426c76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd0c4f86129cfbcfc1db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e225a8f8dd0017c6d14f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28dcae474f1c3b5edda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf5ad5043c9f355f30d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7870a0584c76044d7bef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fe3d102e32a09e1fcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f1d776adbbf6ceb8cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e04748e94909ecbaf60f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7734693b405d82ba16c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h122bdcad50b846820c2fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had1f9a08b7937889c635;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1121c9ad7d5f29c83ea3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha94704d3448c111e9291;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d39b9e5d294b1144452;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134bc4cacd6809fb0be9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e3c528548bcd6c42149;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1313f9b844ebedfaf5b26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b02c5968e9887bd8254;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce840025b61cc004c7b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4dbe27273514eee4533;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9528919af0530f6fdd3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54517ddb0d1bf1acc75c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d675c6c6160ab60a6a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h901e00893bfebd23629d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1876448d12127f10c66c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40a4bb7f2e55d2849c31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a031a20e1356517e1583;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddfc584b6f1eb986a204;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192e368c56943dbed5a10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b20f0a2ea240ab2fa25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h233df089b9c6ffc9afb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e2f0638a2efbaeea64d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3805ca6409642ffb5d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14dd4192abc3e06019f9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd289152802169ea338f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa655f24e922a84395cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1beaed6479df7aa3de70c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c61d95f75bfcf6264ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1053633b523a25fca07f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7086e3f4c5263e05b02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d74c06eb8a1a1db36a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d64a4b2bada38caa2f9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be19f656b8dead216a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9dedc8ea8e37a62a690c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17398ae6586a38ef113;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h601c8d9161ed70309607;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24efffedfc2fc8a6f0af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e7df488d2f78728ddfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7114165581f5754944b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c5232812e15cde93bcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170caf337db6638c73b23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bae16139bbfc0ebe4f7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89a289d19bd5ae5bd5fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb270d5a46894f02adbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ec8d44681cbf0e24823;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0b50d0b3f6434bdd3ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha708814b78cb36f479dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde74534e524da0c602c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e8876fdd9df7fe5e8d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3ae423d8c6bcda166c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7fb465d0fe13dd13e226;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16391dc627023441aede6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e749e479ebe027489483;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h763f2f183ec4013b5d21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he16dcc11f17a3a617644;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13416f22ea500c0be6fb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cb130d52c4f16d0878e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1236cb86af99bacefa50c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h387ad01821c49986bc3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc041e9c1a6fe44f36133;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf23e029c2abc6274f88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52ffff77ad6a727af3f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1094d28aba5a22e48060b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddddfa6218002a56a395;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10483f0752caf95d3b826;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81f99b621aa26701635;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10194c1451f1538c4287e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c56e7fa4a2e3053656e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11daac7dfbf591e4f8b13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc39081493bec052936b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35ded389a0a07cbcd9ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefe636ef8333a008a153;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a2fa7d0e4f9d7db0576;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d8e1de911fa804dc549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb980c234bfc9199d833c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha355ba04b27266caba4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a68de3402e8f576936b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd627db1e508b60b1602;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36a1fdfdb30708d07214;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e89a8d5473a9c0b636e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h528f4d2df9e9768408f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28fbddea690c2f633d52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c697c476a352397dd27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h261705071e9e9a98a276;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he80bf1bd33775dcdc882;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cc0b58bc266e5d70ae1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac856c3a9d853e864527;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8037de15333844c5a01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ac12f0e12c8ef60f666;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc84897432938ea00480;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d30b729e03dea74bb01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f312c5a8bdebc49d859;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190afe857074e9c55a49f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb060e159f3ee1c13eec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b8fa8817660bfd81f2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed48c421b6f1cfcf8ba9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af092621e8856b9f2b0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bc51adacc4c3cf21479;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156926fcee7d891d0b0d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a16df98df53d6dd3107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc118660cb02af1f7875;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1134f7b3ae7e556649d07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7cd66ccc3ae479e07e49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e02ec369b002389f3273;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8f424bb0c7d20324ff1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14be4abda2faebd42b10b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55b25b16700954e0bbc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ef62aeccc080a9030b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f606c6b411eee7bf285;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab715e7889e54d44fb86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a110187a6d952042d94f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h195a20e6115dc24e67a8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h476e579fceea2d4d50e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1606fd2f262ea60881694;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdbef18c1bacc6badbbbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha92655f94afbb1c4b68a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1561e1f348b6782bd66a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbb9deb5f72395cb6d0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbde70c2775045e55e7df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105a2f83c39d9970c9b53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dae87be33b4307cd7517;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bda5b31cb8ed566a5ffd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3d5a077f53ac4ddf2a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c6d1a0f9e4b09bc9008;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h668508655bf495e6602d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1d9dbfd968b198d6f8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14df41e72a69a064c0038;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f76e90ed60b5804862fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf431dd1524e6f9054130;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf2014154238ffc54e95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e597587d49c984d0306;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1761af3160e17d4d34016;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1586800f874bedef8eaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188b63b629a578afda991;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9a1df3322ef055d69c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b538f0c6210fd84486de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a06902c7e0cc380c9125;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0f0ffba562f3ccaa6dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d04e91968a203fc9617;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1237ef0d0355d9d9db672;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac25557611f986ee749a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e7b4aa5228e30709abe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140132eff35eac511fcf8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc4cfe057369dc11faf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175cd2a435edc107ba53b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174d91c164ecc48557fd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139f43601265fc6fdcea4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha279b1be6d90a5f4be1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ec4c6570f285b1514a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8819dcf417b2fe3641d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180ca4bee90c823b38163;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d897a429e86e2f18f5e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54e5a7d157da7511403d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9b4a42299a187ead673;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2fa897348c5fc1591b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h963fc38d6e0bb922ee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d4eab02f3fc5264fb6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2bdbc3a24e3cb3c96479;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44f751ba67b4fcc5e16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4904e6e413f57227cbe0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181aa8f6598cadcf0e1ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef534e8696eefed10533;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f47b047765b869de3d21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124a05ed009aa294cf3d3;
        #1
        $finish();
    end
endmodule
