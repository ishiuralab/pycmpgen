module compressor2_1_189_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, input in_data128, input in_data129, input in_data130, input in_data131, input in_data132, input in_data133, input in_data134, input in_data135, input in_data136, input in_data137, input in_data138, input in_data139, input in_data140, input in_data141, input in_data142, input in_data143, input in_data144, input in_data145, input in_data146, input in_data147, input in_data148, input in_data149, input in_data150, input in_data151, input in_data152, input in_data153, input in_data154, input in_data155, input in_data156, input in_data157, input in_data158, input in_data159, input in_data160, input in_data161, input in_data162, input in_data163, input in_data164, input in_data165, input in_data166, input in_data167, input in_data168, input in_data169, input in_data170, input in_data171, input in_data172, input in_data173, input in_data174, input in_data175, input in_data176, input in_data177, input in_data178, input in_data179, input in_data180, input in_data181, input in_data182, input in_data183, input in_data184, input in_data185, input in_data186, input in_data187, input in_data188, output [19:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    reg [11:0] src128;
    reg [11:0] src129;
    reg [11:0] src130;
    reg [11:0] src131;
    reg [11:0] src132;
    reg [11:0] src133;
    reg [11:0] src134;
    reg [11:0] src135;
    reg [11:0] src136;
    reg [11:0] src137;
    reg [11:0] src138;
    reg [11:0] src139;
    reg [11:0] src140;
    reg [11:0] src141;
    reg [11:0] src142;
    reg [11:0] src143;
    reg [11:0] src144;
    reg [11:0] src145;
    reg [11:0] src146;
    reg [11:0] src147;
    reg [11:0] src148;
    reg [11:0] src149;
    reg [11:0] src150;
    reg [11:0] src151;
    reg [11:0] src152;
    reg [11:0] src153;
    reg [11:0] src154;
    reg [11:0] src155;
    reg [11:0] src156;
    reg [11:0] src157;
    reg [11:0] src158;
    reg [11:0] src159;
    reg [11:0] src160;
    reg [11:0] src161;
    reg [11:0] src162;
    reg [11:0] src163;
    reg [11:0] src164;
    reg [11:0] src165;
    reg [11:0] src166;
    reg [11:0] src167;
    reg [11:0] src168;
    reg [11:0] src169;
    reg [11:0] src170;
    reg [11:0] src171;
    reg [11:0] src172;
    reg [11:0] src173;
    reg [11:0] src174;
    reg [11:0] src175;
    reg [11:0] src176;
    reg [11:0] src177;
    reg [11:0] src178;
    reg [11:0] src179;
    reg [11:0] src180;
    reg [11:0] src181;
    reg [11:0] src182;
    reg [11:0] src183;
    reg [11:0] src184;
    reg [11:0] src185;
    reg [11:0] src186;
    reg [11:0] src187;
    reg [11:0] src188;
    compressor2_1_189_12 compressor2_1_189_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .src128(src128), .src129(src129), .src130(src130), .src131(src131), .src132(src132), .src133(src133), .src134(src134), .src135(src135), .src136(src136), .src137(src137), .src138(src138), .src139(src139), .src140(src140), .src141(src141), .src142(src142), .src143(src143), .src144(src144), .src145(src145), .src146(src146), .src147(src147), .src148(src148), .src149(src149), .src150(src150), .src151(src151), .src152(src152), .src153(src153), .src154(src154), .src155(src155), .src156(src156), .src157(src157), .src158(src158), .src159(src159), .src160(src160), .src161(src161), .src162(src162), .src163(src163), .src164(src164), .src165(src165), .src166(src166), .src167(src167), .src168(src168), .src169(src169), .src170(src170), .src171(src171), .src172(src172), .src173(src173), .src174(src174), .src175(src175), .src176(src176), .src177(src177), .src178(src178), .src179(src179), .src180(src180), .src181(src181), .src182(src182), .src183(src183), .src184(src184), .src185(src185), .src186(src186), .src187(src187), .src188(src188), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
        src128 <= 0;
        src129 <= 0;
        src130 <= 0;
        src131 <= 0;
        src132 <= 0;
        src133 <= 0;
        src134 <= 0;
        src135 <= 0;
        src136 <= 0;
        src137 <= 0;
        src138 <= 0;
        src139 <= 0;
        src140 <= 0;
        src141 <= 0;
        src142 <= 0;
        src143 <= 0;
        src144 <= 0;
        src145 <= 0;
        src146 <= 0;
        src147 <= 0;
        src148 <= 0;
        src149 <= 0;
        src150 <= 0;
        src151 <= 0;
        src152 <= 0;
        src153 <= 0;
        src154 <= 0;
        src155 <= 0;
        src156 <= 0;
        src157 <= 0;
        src158 <= 0;
        src159 <= 0;
        src160 <= 0;
        src161 <= 0;
        src162 <= 0;
        src163 <= 0;
        src164 <= 0;
        src165 <= 0;
        src166 <= 0;
        src167 <= 0;
        src168 <= 0;
        src169 <= 0;
        src170 <= 0;
        src171 <= 0;
        src172 <= 0;
        src173 <= 0;
        src174 <= 0;
        src175 <= 0;
        src176 <= 0;
        src177 <= 0;
        src178 <= 0;
        src179 <= 0;
        src180 <= 0;
        src181 <= 0;
        src182 <= 0;
        src183 <= 0;
        src184 <= 0;
        src185 <= 0;
        src186 <= 0;
        src187 <= 0;
        src188 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
        src32 <= {src32[10:0], in_data32};
        src33 <= {src33[10:0], in_data33};
        src34 <= {src34[10:0], in_data34};
        src35 <= {src35[10:0], in_data35};
        src36 <= {src36[10:0], in_data36};
        src37 <= {src37[10:0], in_data37};
        src38 <= {src38[10:0], in_data38};
        src39 <= {src39[10:0], in_data39};
        src40 <= {src40[10:0], in_data40};
        src41 <= {src41[10:0], in_data41};
        src42 <= {src42[10:0], in_data42};
        src43 <= {src43[10:0], in_data43};
        src44 <= {src44[10:0], in_data44};
        src45 <= {src45[10:0], in_data45};
        src46 <= {src46[10:0], in_data46};
        src47 <= {src47[10:0], in_data47};
        src48 <= {src48[10:0], in_data48};
        src49 <= {src49[10:0], in_data49};
        src50 <= {src50[10:0], in_data50};
        src51 <= {src51[10:0], in_data51};
        src52 <= {src52[10:0], in_data52};
        src53 <= {src53[10:0], in_data53};
        src54 <= {src54[10:0], in_data54};
        src55 <= {src55[10:0], in_data55};
        src56 <= {src56[10:0], in_data56};
        src57 <= {src57[10:0], in_data57};
        src58 <= {src58[10:0], in_data58};
        src59 <= {src59[10:0], in_data59};
        src60 <= {src60[10:0], in_data60};
        src61 <= {src61[10:0], in_data61};
        src62 <= {src62[10:0], in_data62};
        src63 <= {src63[10:0], in_data63};
        src64 <= {src64[10:0], in_data64};
        src65 <= {src65[10:0], in_data65};
        src66 <= {src66[10:0], in_data66};
        src67 <= {src67[10:0], in_data67};
        src68 <= {src68[10:0], in_data68};
        src69 <= {src69[10:0], in_data69};
        src70 <= {src70[10:0], in_data70};
        src71 <= {src71[10:0], in_data71};
        src72 <= {src72[10:0], in_data72};
        src73 <= {src73[10:0], in_data73};
        src74 <= {src74[10:0], in_data74};
        src75 <= {src75[10:0], in_data75};
        src76 <= {src76[10:0], in_data76};
        src77 <= {src77[10:0], in_data77};
        src78 <= {src78[10:0], in_data78};
        src79 <= {src79[10:0], in_data79};
        src80 <= {src80[10:0], in_data80};
        src81 <= {src81[10:0], in_data81};
        src82 <= {src82[10:0], in_data82};
        src83 <= {src83[10:0], in_data83};
        src84 <= {src84[10:0], in_data84};
        src85 <= {src85[10:0], in_data85};
        src86 <= {src86[10:0], in_data86};
        src87 <= {src87[10:0], in_data87};
        src88 <= {src88[10:0], in_data88};
        src89 <= {src89[10:0], in_data89};
        src90 <= {src90[10:0], in_data90};
        src91 <= {src91[10:0], in_data91};
        src92 <= {src92[10:0], in_data92};
        src93 <= {src93[10:0], in_data93};
        src94 <= {src94[10:0], in_data94};
        src95 <= {src95[10:0], in_data95};
        src96 <= {src96[10:0], in_data96};
        src97 <= {src97[10:0], in_data97};
        src98 <= {src98[10:0], in_data98};
        src99 <= {src99[10:0], in_data99};
        src100 <= {src100[10:0], in_data100};
        src101 <= {src101[10:0], in_data101};
        src102 <= {src102[10:0], in_data102};
        src103 <= {src103[10:0], in_data103};
        src104 <= {src104[10:0], in_data104};
        src105 <= {src105[10:0], in_data105};
        src106 <= {src106[10:0], in_data106};
        src107 <= {src107[10:0], in_data107};
        src108 <= {src108[10:0], in_data108};
        src109 <= {src109[10:0], in_data109};
        src110 <= {src110[10:0], in_data110};
        src111 <= {src111[10:0], in_data111};
        src112 <= {src112[10:0], in_data112};
        src113 <= {src113[10:0], in_data113};
        src114 <= {src114[10:0], in_data114};
        src115 <= {src115[10:0], in_data115};
        src116 <= {src116[10:0], in_data116};
        src117 <= {src117[10:0], in_data117};
        src118 <= {src118[10:0], in_data118};
        src119 <= {src119[10:0], in_data119};
        src120 <= {src120[10:0], in_data120};
        src121 <= {src121[10:0], in_data121};
        src122 <= {src122[10:0], in_data122};
        src123 <= {src123[10:0], in_data123};
        src124 <= {src124[10:0], in_data124};
        src125 <= {src125[10:0], in_data125};
        src126 <= {src126[10:0], in_data126};
        src127 <= {src127[10:0], in_data127};
        src128 <= {src128[10:0], in_data128};
        src129 <= {src129[10:0], in_data129};
        src130 <= {src130[10:0], in_data130};
        src131 <= {src131[10:0], in_data131};
        src132 <= {src132[10:0], in_data132};
        src133 <= {src133[10:0], in_data133};
        src134 <= {src134[10:0], in_data134};
        src135 <= {src135[10:0], in_data135};
        src136 <= {src136[10:0], in_data136};
        src137 <= {src137[10:0], in_data137};
        src138 <= {src138[10:0], in_data138};
        src139 <= {src139[10:0], in_data139};
        src140 <= {src140[10:0], in_data140};
        src141 <= {src141[10:0], in_data141};
        src142 <= {src142[10:0], in_data142};
        src143 <= {src143[10:0], in_data143};
        src144 <= {src144[10:0], in_data144};
        src145 <= {src145[10:0], in_data145};
        src146 <= {src146[10:0], in_data146};
        src147 <= {src147[10:0], in_data147};
        src148 <= {src148[10:0], in_data148};
        src149 <= {src149[10:0], in_data149};
        src150 <= {src150[10:0], in_data150};
        src151 <= {src151[10:0], in_data151};
        src152 <= {src152[10:0], in_data152};
        src153 <= {src153[10:0], in_data153};
        src154 <= {src154[10:0], in_data154};
        src155 <= {src155[10:0], in_data155};
        src156 <= {src156[10:0], in_data156};
        src157 <= {src157[10:0], in_data157};
        src158 <= {src158[10:0], in_data158};
        src159 <= {src159[10:0], in_data159};
        src160 <= {src160[10:0], in_data160};
        src161 <= {src161[10:0], in_data161};
        src162 <= {src162[10:0], in_data162};
        src163 <= {src163[10:0], in_data163};
        src164 <= {src164[10:0], in_data164};
        src165 <= {src165[10:0], in_data165};
        src166 <= {src166[10:0], in_data166};
        src167 <= {src167[10:0], in_data167};
        src168 <= {src168[10:0], in_data168};
        src169 <= {src169[10:0], in_data169};
        src170 <= {src170[10:0], in_data170};
        src171 <= {src171[10:0], in_data171};
        src172 <= {src172[10:0], in_data172};
        src173 <= {src173[10:0], in_data173};
        src174 <= {src174[10:0], in_data174};
        src175 <= {src175[10:0], in_data175};
        src176 <= {src176[10:0], in_data176};
        src177 <= {src177[10:0], in_data177};
        src178 <= {src178[10:0], in_data178};
        src179 <= {src179[10:0], in_data179};
        src180 <= {src180[10:0], in_data180};
        src181 <= {src181[10:0], in_data181};
        src182 <= {src182[10:0], in_data182};
        src183 <= {src183[10:0], in_data183};
        src184 <= {src184[10:0], in_data184};
        src185 <= {src185[10:0], in_data185};
        src186 <= {src186[10:0], in_data186};
        src187 <= {src187[10:0], in_data187};
        src188 <= {src188[10:0], in_data188};
    end
endmodule

module compressor2_1_189_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    input [11:0]src32,
    input [11:0]src33,
    input [11:0]src34,
    input [11:0]src35,
    input [11:0]src36,
    input [11:0]src37,
    input [11:0]src38,
    input [11:0]src39,
    input [11:0]src40,
    input [11:0]src41,
    input [11:0]src42,
    input [11:0]src43,
    input [11:0]src44,
    input [11:0]src45,
    input [11:0]src46,
    input [11:0]src47,
    input [11:0]src48,
    input [11:0]src49,
    input [11:0]src50,
    input [11:0]src51,
    input [11:0]src52,
    input [11:0]src53,
    input [11:0]src54,
    input [11:0]src55,
    input [11:0]src56,
    input [11:0]src57,
    input [11:0]src58,
    input [11:0]src59,
    input [11:0]src60,
    input [11:0]src61,
    input [11:0]src62,
    input [11:0]src63,
    input [11:0]src64,
    input [11:0]src65,
    input [11:0]src66,
    input [11:0]src67,
    input [11:0]src68,
    input [11:0]src69,
    input [11:0]src70,
    input [11:0]src71,
    input [11:0]src72,
    input [11:0]src73,
    input [11:0]src74,
    input [11:0]src75,
    input [11:0]src76,
    input [11:0]src77,
    input [11:0]src78,
    input [11:0]src79,
    input [11:0]src80,
    input [11:0]src81,
    input [11:0]src82,
    input [11:0]src83,
    input [11:0]src84,
    input [11:0]src85,
    input [11:0]src86,
    input [11:0]src87,
    input [11:0]src88,
    input [11:0]src89,
    input [11:0]src90,
    input [11:0]src91,
    input [11:0]src92,
    input [11:0]src93,
    input [11:0]src94,
    input [11:0]src95,
    input [11:0]src96,
    input [11:0]src97,
    input [11:0]src98,
    input [11:0]src99,
    input [11:0]src100,
    input [11:0]src101,
    input [11:0]src102,
    input [11:0]src103,
    input [11:0]src104,
    input [11:0]src105,
    input [11:0]src106,
    input [11:0]src107,
    input [11:0]src108,
    input [11:0]src109,
    input [11:0]src110,
    input [11:0]src111,
    input [11:0]src112,
    input [11:0]src113,
    input [11:0]src114,
    input [11:0]src115,
    input [11:0]src116,
    input [11:0]src117,
    input [11:0]src118,
    input [11:0]src119,
    input [11:0]src120,
    input [11:0]src121,
    input [11:0]src122,
    input [11:0]src123,
    input [11:0]src124,
    input [11:0]src125,
    input [11:0]src126,
    input [11:0]src127,
    input [11:0]src128,
    input [11:0]src129,
    input [11:0]src130,
    input [11:0]src131,
    input [11:0]src132,
    input [11:0]src133,
    input [11:0]src134,
    input [11:0]src135,
    input [11:0]src136,
    input [11:0]src137,
    input [11:0]src138,
    input [11:0]src139,
    input [11:0]src140,
    input [11:0]src141,
    input [11:0]src142,
    input [11:0]src143,
    input [11:0]src144,
    input [11:0]src145,
    input [11:0]src146,
    input [11:0]src147,
    input [11:0]src148,
    input [11:0]src149,
    input [11:0]src150,
    input [11:0]src151,
    input [11:0]src152,
    input [11:0]src153,
    input [11:0]src154,
    input [11:0]src155,
    input [11:0]src156,
    input [11:0]src157,
    input [11:0]src158,
    input [11:0]src159,
    input [11:0]src160,
    input [11:0]src161,
    input [11:0]src162,
    input [11:0]src163,
    input [11:0]src164,
    input [11:0]src165,
    input [11:0]src166,
    input [11:0]src167,
    input [11:0]src168,
    input [11:0]src169,
    input [11:0]src170,
    input [11:0]src171,
    input [11:0]src172,
    input [11:0]src173,
    input [11:0]src174,
    input [11:0]src175,
    input [11:0]src176,
    input [11:0]src177,
    input [11:0]src178,
    input [11:0]src179,
    input [11:0]src180,
    input [11:0]src181,
    input [11:0]src182,
    input [11:0]src183,
    input [11:0]src184,
    input [11:0]src185,
    input [11:0]src186,
    input [11:0]src187,
    input [11:0]src188,
    output [19:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [0:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [0:0] comp_out18;
    wire [0:0] comp_out19;
    wire [20:0] out;
    compressor compressor_inst(
        .src0({src188[0], src187[0], src186[0], src185[0], src184[0], src183[0], src182[0], src181[0], src180[0], src179[0], src178[0], src177[0], src176[0], src175[0], src174[0], src173[0], src172[0], src171[0], src170[0], src169[0], src168[0], src167[0], src166[0], src165[0], src164[0], src163[0], src162[0], src161[0], src160[0], src159[0], src158[0], src157[0], src156[0], src155[0], src154[0], src153[0], src152[0], src151[0], src150[0], src149[0], src148[0], src147[0], src146[0], src145[0], src144[0], src143[0], src142[0], src141[0], src140[0], src139[0], src138[0], src137[0], src136[0], src135[0], src134[0], src133[0], src132[0], src131[0], src130[0], src129[0], src128[0], src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src188[1], src187[1], src186[1], src185[1], src184[1], src183[1], src182[1], src181[1], src180[1], src179[1], src178[1], src177[1], src176[1], src175[1], src174[1], src173[1], src172[1], src171[1], src170[1], src169[1], src168[1], src167[1], src166[1], src165[1], src164[1], src163[1], src162[1], src161[1], src160[1], src159[1], src158[1], src157[1], src156[1], src155[1], src154[1], src153[1], src152[1], src151[1], src150[1], src149[1], src148[1], src147[1], src146[1], src145[1], src144[1], src143[1], src142[1], src141[1], src140[1], src139[1], src138[1], src137[1], src136[1], src135[1], src134[1], src133[1], src132[1], src131[1], src130[1], src129[1], src128[1], src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src188[2], src187[2], src186[2], src185[2], src184[2], src183[2], src182[2], src181[2], src180[2], src179[2], src178[2], src177[2], src176[2], src175[2], src174[2], src173[2], src172[2], src171[2], src170[2], src169[2], src168[2], src167[2], src166[2], src165[2], src164[2], src163[2], src162[2], src161[2], src160[2], src159[2], src158[2], src157[2], src156[2], src155[2], src154[2], src153[2], src152[2], src151[2], src150[2], src149[2], src148[2], src147[2], src146[2], src145[2], src144[2], src143[2], src142[2], src141[2], src140[2], src139[2], src138[2], src137[2], src136[2], src135[2], src134[2], src133[2], src132[2], src131[2], src130[2], src129[2], src128[2], src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src188[3], src187[3], src186[3], src185[3], src184[3], src183[3], src182[3], src181[3], src180[3], src179[3], src178[3], src177[3], src176[3], src175[3], src174[3], src173[3], src172[3], src171[3], src170[3], src169[3], src168[3], src167[3], src166[3], src165[3], src164[3], src163[3], src162[3], src161[3], src160[3], src159[3], src158[3], src157[3], src156[3], src155[3], src154[3], src153[3], src152[3], src151[3], src150[3], src149[3], src148[3], src147[3], src146[3], src145[3], src144[3], src143[3], src142[3], src141[3], src140[3], src139[3], src138[3], src137[3], src136[3], src135[3], src134[3], src133[3], src132[3], src131[3], src130[3], src129[3], src128[3], src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src188[4], src187[4], src186[4], src185[4], src184[4], src183[4], src182[4], src181[4], src180[4], src179[4], src178[4], src177[4], src176[4], src175[4], src174[4], src173[4], src172[4], src171[4], src170[4], src169[4], src168[4], src167[4], src166[4], src165[4], src164[4], src163[4], src162[4], src161[4], src160[4], src159[4], src158[4], src157[4], src156[4], src155[4], src154[4], src153[4], src152[4], src151[4], src150[4], src149[4], src148[4], src147[4], src146[4], src145[4], src144[4], src143[4], src142[4], src141[4], src140[4], src139[4], src138[4], src137[4], src136[4], src135[4], src134[4], src133[4], src132[4], src131[4], src130[4], src129[4], src128[4], src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src188[5], src187[5], src186[5], src185[5], src184[5], src183[5], src182[5], src181[5], src180[5], src179[5], src178[5], src177[5], src176[5], src175[5], src174[5], src173[5], src172[5], src171[5], src170[5], src169[5], src168[5], src167[5], src166[5], src165[5], src164[5], src163[5], src162[5], src161[5], src160[5], src159[5], src158[5], src157[5], src156[5], src155[5], src154[5], src153[5], src152[5], src151[5], src150[5], src149[5], src148[5], src147[5], src146[5], src145[5], src144[5], src143[5], src142[5], src141[5], src140[5], src139[5], src138[5], src137[5], src136[5], src135[5], src134[5], src133[5], src132[5], src131[5], src130[5], src129[5], src128[5], src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src188[6], src187[6], src186[6], src185[6], src184[6], src183[6], src182[6], src181[6], src180[6], src179[6], src178[6], src177[6], src176[6], src175[6], src174[6], src173[6], src172[6], src171[6], src170[6], src169[6], src168[6], src167[6], src166[6], src165[6], src164[6], src163[6], src162[6], src161[6], src160[6], src159[6], src158[6], src157[6], src156[6], src155[6], src154[6], src153[6], src152[6], src151[6], src150[6], src149[6], src148[6], src147[6], src146[6], src145[6], src144[6], src143[6], src142[6], src141[6], src140[6], src139[6], src138[6], src137[6], src136[6], src135[6], src134[6], src133[6], src132[6], src131[6], src130[6], src129[6], src128[6], src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src188[7], src187[7], src186[7], src185[7], src184[7], src183[7], src182[7], src181[7], src180[7], src179[7], src178[7], src177[7], src176[7], src175[7], src174[7], src173[7], src172[7], src171[7], src170[7], src169[7], src168[7], src167[7], src166[7], src165[7], src164[7], src163[7], src162[7], src161[7], src160[7], src159[7], src158[7], src157[7], src156[7], src155[7], src154[7], src153[7], src152[7], src151[7], src150[7], src149[7], src148[7], src147[7], src146[7], src145[7], src144[7], src143[7], src142[7], src141[7], src140[7], src139[7], src138[7], src137[7], src136[7], src135[7], src134[7], src133[7], src132[7], src131[7], src130[7], src129[7], src128[7], src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src188[8], src187[8], src186[8], src185[8], src184[8], src183[8], src182[8], src181[8], src180[8], src179[8], src178[8], src177[8], src176[8], src175[8], src174[8], src173[8], src172[8], src171[8], src170[8], src169[8], src168[8], src167[8], src166[8], src165[8], src164[8], src163[8], src162[8], src161[8], src160[8], src159[8], src158[8], src157[8], src156[8], src155[8], src154[8], src153[8], src152[8], src151[8], src150[8], src149[8], src148[8], src147[8], src146[8], src145[8], src144[8], src143[8], src142[8], src141[8], src140[8], src139[8], src138[8], src137[8], src136[8], src135[8], src134[8], src133[8], src132[8], src131[8], src130[8], src129[8], src128[8], src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src188[9], src187[9], src186[9], src185[9], src184[9], src183[9], src182[9], src181[9], src180[9], src179[9], src178[9], src177[9], src176[9], src175[9], src174[9], src173[9], src172[9], src171[9], src170[9], src169[9], src168[9], src167[9], src166[9], src165[9], src164[9], src163[9], src162[9], src161[9], src160[9], src159[9], src158[9], src157[9], src156[9], src155[9], src154[9], src153[9], src152[9], src151[9], src150[9], src149[9], src148[9], src147[9], src146[9], src145[9], src144[9], src143[9], src142[9], src141[9], src140[9], src139[9], src138[9], src137[9], src136[9], src135[9], src134[9], src133[9], src132[9], src131[9], src130[9], src129[9], src128[9], src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src188[10], src187[10], src186[10], src185[10], src184[10], src183[10], src182[10], src181[10], src180[10], src179[10], src178[10], src177[10], src176[10], src175[10], src174[10], src173[10], src172[10], src171[10], src170[10], src169[10], src168[10], src167[10], src166[10], src165[10], src164[10], src163[10], src162[10], src161[10], src160[10], src159[10], src158[10], src157[10], src156[10], src155[10], src154[10], src153[10], src152[10], src151[10], src150[10], src149[10], src148[10], src147[10], src146[10], src145[10], src144[10], src143[10], src142[10], src141[10], src140[10], src139[10], src138[10], src137[10], src136[10], src135[10], src134[10], src133[10], src132[10], src131[10], src130[10], src129[10], src128[10], src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src188[11], src187[11], src186[11], src185[11], src184[11], src183[11], src182[11], src181[11], src180[11], src179[11], src178[11], src177[11], src176[11], src175[11], src174[11], src173[11], src172[11], src171[11], src170[11], src169[11], src168[11], src167[11], src166[11], src165[11], src164[11], src163[11], src162[11], src161[11], src160[11], src159[11], src158[11], src157[11], src156[11], src155[11], src154[11], src153[11], src152[11], src151[11], src150[11], src149[11], src148[11], src147[11], src146[11], src145[11], src144[11], src143[11], src142[11], src141[11], src140[11], src139[11], src138[11], src137[11], src136[11], src135[11], src134[11], src133[11], src132[11], src131[11], src130[11], src129[11], src128[11], src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    rowadder2_1_20 rowadder2_1inst(
        .src0({comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], 1'h0, comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[19:0];
endmodule
module compressor (
      input wire [188:0] src0,
      input wire [188:0] src1,
      input wire [188:0] src2,
      input wire [188:0] src3,
      input wire [188:0] src4,
      input wire [188:0] src5,
      input wire [188:0] src6,
      input wire [188:0] src7,
      input wire [188:0] src8,
      input wire [188:0] src9,
      input wire [188:0] src10,
      input wire [188:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [0:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [0:0] dst18,
      output wire [0:0] dst19);

   wire [188:0] stage0_0;
   wire [188:0] stage0_1;
   wire [188:0] stage0_2;
   wire [188:0] stage0_3;
   wire [188:0] stage0_4;
   wire [188:0] stage0_5;
   wire [188:0] stage0_6;
   wire [188:0] stage0_7;
   wire [188:0] stage0_8;
   wire [188:0] stage0_9;
   wire [188:0] stage0_10;
   wire [188:0] stage0_11;
   wire [37:0] stage1_0;
   wire [71:0] stage1_1;
   wire [73:0] stage1_2;
   wire [64:0] stage1_3;
   wire [94:0] stage1_4;
   wire [85:0] stage1_5;
   wire [70:0] stage1_6;
   wire [77:0] stage1_7;
   wire [96:0] stage1_8;
   wire [89:0] stage1_9;
   wire [67:0] stage1_10;
   wire [110:0] stage1_11;
   wire [52:0] stage1_12;
   wire [22:0] stage1_13;
   wire [15:0] stage2_0;
   wire [23:0] stage2_1;
   wire [23:0] stage2_2;
   wire [30:0] stage2_3;
   wire [31:0] stage2_4;
   wire [35:0] stage2_5;
   wire [38:0] stage2_6;
   wire [27:0] stage2_7;
   wire [30:0] stage2_8;
   wire [41:0] stage2_9;
   wire [37:0] stage2_10;
   wire [48:0] stage2_11;
   wire [47:0] stage2_12;
   wire [36:0] stage2_13;
   wire [5:0] stage2_14;
   wire [0:0] stage2_15;
   wire [6:0] stage3_0;
   wire [14:0] stage3_1;
   wire [5:0] stage3_2;
   wire [12:0] stage3_3;
   wire [12:0] stage3_4;
   wire [25:0] stage3_5;
   wire [12:0] stage3_6;
   wire [17:0] stage3_7;
   wire [11:0] stage3_8;
   wire [10:0] stage3_9;
   wire [22:0] stage3_10;
   wire [17:0] stage3_11;
   wire [26:0] stage3_12;
   wire [14:0] stage3_13;
   wire [11:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [10:0] stage4_1;
   wire [1:0] stage4_2;
   wire [4:0] stage4_3;
   wire [4:0] stage4_4;
   wire [9:0] stage4_5;
   wire [5:0] stage4_6;
   wire [5:0] stage4_7;
   wire [6:0] stage4_8;
   wire [11:0] stage4_9;
   wire [4:0] stage4_10;
   wire [6:0] stage4_11;
   wire [10:0] stage4_12;
   wire [9:0] stage4_13;
   wire [5:0] stage4_14;
   wire [11:0] stage4_15;
   wire [2:0] stage4_16;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [3:0] stage5_4;
   wire [6:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [2:0] stage5_8;
   wire [4:0] stage5_9;
   wire [4:0] stage5_10;
   wire [1:0] stage5_11;
   wire [5:0] stage5_12;
   wire [4:0] stage5_13;
   wire [2:0] stage5_14;
   wire [2:0] stage5_15;
   wire [5:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [0:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [0:0] stage6_18;
   wire [0:0] stage6_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[5]},
      {stage0_3[7]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[12],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[13],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[14],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[15],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[16],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[17],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[18],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[19],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[20],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[21],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[22],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[23],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc615_5 gpc57 (
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172]},
      {stage0_3[152]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[24],stage1_4[57],stage1_3[57],stage1_2[57]}
   );
   gpc606_5 gpc58 (
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[25],stage1_4[58],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163]},
      {stage0_4[6]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[2],stage1_5[26],stage1_4[59],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage0_4[7]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[3],stage1_5[27],stage1_4[60],stage1_3[60]}
   );
   gpc615_5 gpc61 (
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173]},
      {stage0_4[8]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[4],stage1_5[28],stage1_4[61],stage1_3[61]}
   );
   gpc615_5 gpc62 (
      {stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage0_4[9]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[5],stage1_5[29],stage1_4[62],stage1_3[62]}
   );
   gpc615_5 gpc63 (
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183]},
      {stage0_4[10]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[6],stage1_5[30],stage1_4[63],stage1_3[63]}
   );
   gpc615_5 gpc64 (
      {stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage0_4[11]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[7],stage1_5[31],stage1_4[64],stage1_3[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[7],stage1_6[8],stage1_5[32],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[8],stage1_6[9],stage1_5[33],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[9],stage1_6[10],stage1_5[34],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[10],stage1_6[11],stage1_5[35],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[11],stage1_6[12],stage1_5[36],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[12],stage1_6[13],stage1_5[37],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[13],stage1_6[14],stage1_5[38],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[14],stage1_6[15],stage1_5[39],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[15],stage1_6[16],stage1_5[40],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[16],stage1_6[17],stage1_5[41],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[17],stage1_6[18],stage1_5[42],stage1_4[75]}
   );
   gpc606_5 gpc76 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[18],stage1_6[19],stage1_5[43],stage1_4[76]}
   );
   gpc606_5 gpc77 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[19],stage1_6[20],stage1_5[44],stage1_4[77]}
   );
   gpc606_5 gpc78 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[20],stage1_6[21],stage1_5[45],stage1_4[78]}
   );
   gpc606_5 gpc79 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[21],stage1_6[22],stage1_5[46],stage1_4[79]}
   );
   gpc606_5 gpc80 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[22],stage1_6[23],stage1_5[47],stage1_4[80]}
   );
   gpc606_5 gpc81 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[23],stage1_6[24],stage1_5[48],stage1_4[81]}
   );
   gpc606_5 gpc82 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[24],stage1_6[25],stage1_5[49],stage1_4[82]}
   );
   gpc606_5 gpc83 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[25],stage1_6[26],stage1_5[50],stage1_4[83]}
   );
   gpc606_5 gpc84 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[26],stage1_6[27],stage1_5[51],stage1_4[84]}
   );
   gpc606_5 gpc85 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[27],stage1_6[28],stage1_5[52],stage1_4[85]}
   );
   gpc606_5 gpc86 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[28],stage1_6[29],stage1_5[53],stage1_4[86]}
   );
   gpc606_5 gpc87 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[29],stage1_6[30],stage1_5[54],stage1_4[87]}
   );
   gpc606_5 gpc88 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[30],stage1_6[31],stage1_5[55],stage1_4[88]}
   );
   gpc606_5 gpc89 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[31],stage1_6[32],stage1_5[56],stage1_4[89]}
   );
   gpc606_5 gpc90 (
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[32],stage1_6[33],stage1_5[57],stage1_4[90]}
   );
   gpc606_5 gpc91 (
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[33],stage1_6[34],stage1_5[58],stage1_4[91]}
   );
   gpc615_5 gpc92 (
      {stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_5[42]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[34],stage1_6[35],stage1_5[59],stage1_4[92]}
   );
   gpc615_5 gpc93 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_5[43]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[35],stage1_6[36],stage1_5[60],stage1_4[93]}
   );
   gpc615_5 gpc94 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188]},
      {stage0_5[44]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[36],stage1_6[37],stage1_5[61],stage1_4[94]}
   );
   gpc606_5 gpc95 (
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[30],stage1_7[37],stage1_6[38],stage1_5[62]}
   );
   gpc606_5 gpc96 (
      {stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[31],stage1_7[38],stage1_6[39],stage1_5[63]}
   );
   gpc606_5 gpc97 (
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[32],stage1_7[39],stage1_6[40],stage1_5[64]}
   );
   gpc606_5 gpc98 (
      {stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67], stage0_5[68]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[33],stage1_7[40],stage1_6[41],stage1_5[65]}
   );
   gpc606_5 gpc99 (
      {stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73], stage0_5[74]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[34],stage1_7[41],stage1_6[42],stage1_5[66]}
   );
   gpc606_5 gpc100 (
      {stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79], stage0_5[80]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[35],stage1_7[42],stage1_6[43],stage1_5[67]}
   );
   gpc606_5 gpc101 (
      {stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85], stage0_5[86]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[36],stage1_7[43],stage1_6[44],stage1_5[68]}
   );
   gpc606_5 gpc102 (
      {stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91], stage0_5[92]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[37],stage1_7[44],stage1_6[45],stage1_5[69]}
   );
   gpc606_5 gpc103 (
      {stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97], stage0_5[98]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[38],stage1_7[45],stage1_6[46],stage1_5[70]}
   );
   gpc606_5 gpc104 (
      {stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103], stage0_5[104]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[39],stage1_7[46],stage1_6[47],stage1_5[71]}
   );
   gpc606_5 gpc105 (
      {stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109], stage0_5[110]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[40],stage1_7[47],stage1_6[48],stage1_5[72]}
   );
   gpc606_5 gpc106 (
      {stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[41],stage1_7[48],stage1_6[49],stage1_5[73]}
   );
   gpc606_5 gpc107 (
      {stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[42],stage1_7[49],stage1_6[50],stage1_5[74]}
   );
   gpc606_5 gpc108 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127], stage0_5[128]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[43],stage1_7[50],stage1_6[51],stage1_5[75]}
   );
   gpc606_5 gpc109 (
      {stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133], stage0_5[134]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[44],stage1_7[51],stage1_6[52],stage1_5[76]}
   );
   gpc606_5 gpc110 (
      {stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139], stage0_5[140]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[45],stage1_7[52],stage1_6[53],stage1_5[77]}
   );
   gpc606_5 gpc111 (
      {stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145], stage0_5[146]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[46],stage1_7[53],stage1_6[54],stage1_5[78]}
   );
   gpc606_5 gpc112 (
      {stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151], stage0_5[152]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[47],stage1_7[54],stage1_6[55],stage1_5[79]}
   );
   gpc606_5 gpc113 (
      {stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[48],stage1_7[55],stage1_6[56],stage1_5[80]}
   );
   gpc606_5 gpc114 (
      {stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163], stage0_5[164]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[49],stage1_7[56],stage1_6[57],stage1_5[81]}
   );
   gpc606_5 gpc115 (
      {stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169], stage0_5[170]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[50],stage1_7[57],stage1_6[58],stage1_5[82]}
   );
   gpc606_5 gpc116 (
      {stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175], stage0_5[176]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[51],stage1_7[58],stage1_6[59],stage1_5[83]}
   );
   gpc606_5 gpc117 (
      {stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181], stage0_5[182]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[52],stage1_7[59],stage1_6[60],stage1_5[84]}
   );
   gpc606_5 gpc118 (
      {stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187], stage0_5[188]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[53],stage1_7[60],stage1_6[61],stage1_5[85]}
   );
   gpc615_5 gpc119 (
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148]},
      {stage0_8[0]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[24],stage1_8[54],stage1_7[61]}
   );
   gpc615_5 gpc120 (
      {stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153]},
      {stage0_8[1]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[1],stage1_9[25],stage1_8[55],stage1_7[62]}
   );
   gpc615_5 gpc121 (
      {stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157], stage0_7[158]},
      {stage0_8[2]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[2],stage1_9[26],stage1_8[56],stage1_7[63]}
   );
   gpc615_5 gpc122 (
      {stage0_7[159], stage0_7[160], stage0_7[161], stage0_7[162], stage0_7[163]},
      {stage0_8[3]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[3],stage1_9[27],stage1_8[57],stage1_7[64]}
   );
   gpc615_5 gpc123 (
      {stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167], stage0_7[168]},
      {stage0_8[4]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[4],stage1_9[28],stage1_8[58],stage1_7[65]}
   );
   gpc615_5 gpc124 (
      {stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage0_8[5]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[5],stage1_9[29],stage1_8[59],stage1_7[66]}
   );
   gpc615_5 gpc125 (
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178]},
      {stage0_8[6]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[6],stage1_9[30],stage1_8[60],stage1_7[67]}
   );
   gpc606_5 gpc126 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[7],stage1_10[7],stage1_9[31],stage1_8[61]}
   );
   gpc606_5 gpc127 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[8],stage1_10[8],stage1_9[32],stage1_8[62]}
   );
   gpc606_5 gpc128 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[9],stage1_10[9],stage1_9[33],stage1_8[63]}
   );
   gpc606_5 gpc129 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[10],stage1_10[10],stage1_9[34],stage1_8[64]}
   );
   gpc606_5 gpc130 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[11],stage1_10[11],stage1_9[35],stage1_8[65]}
   );
   gpc606_5 gpc131 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[12],stage1_10[12],stage1_9[36],stage1_8[66]}
   );
   gpc606_5 gpc132 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[13],stage1_10[13],stage1_9[37],stage1_8[67]}
   );
   gpc606_5 gpc133 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[14],stage1_10[14],stage1_9[38],stage1_8[68]}
   );
   gpc606_5 gpc134 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[15],stage1_10[15],stage1_9[39],stage1_8[69]}
   );
   gpc606_5 gpc135 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[16],stage1_10[16],stage1_9[40],stage1_8[70]}
   );
   gpc606_5 gpc136 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[17],stage1_10[17],stage1_9[41],stage1_8[71]}
   );
   gpc606_5 gpc137 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[18],stage1_10[18],stage1_9[42],stage1_8[72]}
   );
   gpc606_5 gpc138 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[19],stage1_10[19],stage1_9[43],stage1_8[73]}
   );
   gpc606_5 gpc139 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[20],stage1_10[20],stage1_9[44],stage1_8[74]}
   );
   gpc606_5 gpc140 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[21],stage1_10[21],stage1_9[45],stage1_8[75]}
   );
   gpc606_5 gpc141 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[22],stage1_10[22],stage1_9[46],stage1_8[76]}
   );
   gpc606_5 gpc142 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[23],stage1_10[23],stage1_9[47],stage1_8[77]}
   );
   gpc606_5 gpc143 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[24],stage1_10[24],stage1_9[48],stage1_8[78]}
   );
   gpc606_5 gpc144 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[25],stage1_10[25],stage1_9[49],stage1_8[79]}
   );
   gpc606_5 gpc145 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[26],stage1_10[26],stage1_9[50],stage1_8[80]}
   );
   gpc606_5 gpc146 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[27],stage1_10[27],stage1_9[51],stage1_8[81]}
   );
   gpc606_5 gpc147 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[28],stage1_10[28],stage1_9[52],stage1_8[82]}
   );
   gpc606_5 gpc148 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[29],stage1_10[29],stage1_9[53],stage1_8[83]}
   );
   gpc606_5 gpc149 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[30],stage1_10[30],stage1_9[54],stage1_8[84]}
   );
   gpc606_5 gpc150 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[31],stage1_10[31],stage1_9[55],stage1_8[85]}
   );
   gpc606_5 gpc151 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[32],stage1_10[32],stage1_9[56],stage1_8[86]}
   );
   gpc615_5 gpc152 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_9[42]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[33],stage1_10[33],stage1_9[57],stage1_8[87]}
   );
   gpc615_5 gpc153 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172]},
      {stage0_9[43]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[34],stage1_10[34],stage1_9[58],stage1_8[88]}
   );
   gpc615_5 gpc154 (
      {stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_9[44]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[35],stage1_10[35],stage1_9[59],stage1_8[89]}
   );
   gpc615_5 gpc155 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_9[45]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[36],stage1_10[36],stage1_9[60],stage1_8[90]}
   );
   gpc606_5 gpc156 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[30],stage1_11[37],stage1_10[37],stage1_9[61]}
   );
   gpc606_5 gpc157 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[31],stage1_11[38],stage1_10[38],stage1_9[62]}
   );
   gpc606_5 gpc158 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[32],stage1_11[39],stage1_10[39],stage1_9[63]}
   );
   gpc606_5 gpc159 (
      {stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[33],stage1_11[40],stage1_10[40],stage1_9[64]}
   );
   gpc606_5 gpc160 (
      {stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[34],stage1_11[41],stage1_10[41],stage1_9[65]}
   );
   gpc606_5 gpc161 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[35],stage1_11[42],stage1_10[42],stage1_9[66]}
   );
   gpc606_5 gpc162 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[36],stage1_11[43],stage1_10[43],stage1_9[67]}
   );
   gpc606_5 gpc163 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[37],stage1_11[44],stage1_10[44],stage1_9[68]}
   );
   gpc606_5 gpc164 (
      {stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[38],stage1_11[45],stage1_10[45],stage1_9[69]}
   );
   gpc606_5 gpc165 (
      {stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[39],stage1_11[46],stage1_10[46],stage1_9[70]}
   );
   gpc606_5 gpc166 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[40],stage1_11[47],stage1_10[47],stage1_9[71]}
   );
   gpc606_5 gpc167 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[41],stage1_11[48],stage1_10[48],stage1_9[72]}
   );
   gpc606_5 gpc168 (
      {stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[42],stage1_11[49],stage1_10[49],stage1_9[73]}
   );
   gpc606_5 gpc169 (
      {stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[43],stage1_11[50],stage1_10[50],stage1_9[74]}
   );
   gpc606_5 gpc170 (
      {stage0_9[130], stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[44],stage1_11[51],stage1_10[51],stage1_9[75]}
   );
   gpc606_5 gpc171 (
      {stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[45],stage1_11[52],stage1_10[52],stage1_9[76]}
   );
   gpc606_5 gpc172 (
      {stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[46],stage1_11[53],stage1_10[53],stage1_9[77]}
   );
   gpc606_5 gpc173 (
      {stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[47],stage1_11[54],stage1_10[54],stage1_9[78]}
   );
   gpc606_5 gpc174 (
      {stage0_9[154], stage0_9[155], stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[48],stage1_11[55],stage1_10[55],stage1_9[79]}
   );
   gpc606_5 gpc175 (
      {stage0_9[160], stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[49],stage1_11[56],stage1_10[56],stage1_9[80]}
   );
   gpc606_5 gpc176 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[50],stage1_11[57],stage1_10[57],stage1_9[81]}
   );
   gpc606_5 gpc177 (
      {stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[51],stage1_11[58],stage1_10[58],stage1_9[82]}
   );
   gpc615_5 gpc178 (
      {stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182]},
      {stage0_10[180]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[52],stage1_11[59],stage1_10[59],stage1_9[83]}
   );
   gpc1_1 gpc179 (
      {stage0_0[184]},
      {stage1_0[33]}
   );
   gpc1_1 gpc180 (
      {stage0_0[185]},
      {stage1_0[34]}
   );
   gpc1_1 gpc181 (
      {stage0_0[186]},
      {stage1_0[35]}
   );
   gpc1_1 gpc182 (
      {stage0_0[187]},
      {stage1_0[36]}
   );
   gpc1_1 gpc183 (
      {stage0_0[188]},
      {stage1_0[37]}
   );
   gpc1_1 gpc184 (
      {stage0_1[174]},
      {stage1_1[57]}
   );
   gpc1_1 gpc185 (
      {stage0_1[175]},
      {stage1_1[58]}
   );
   gpc1_1 gpc186 (
      {stage0_1[176]},
      {stage1_1[59]}
   );
   gpc1_1 gpc187 (
      {stage0_1[177]},
      {stage1_1[60]}
   );
   gpc1_1 gpc188 (
      {stage0_1[178]},
      {stage1_1[61]}
   );
   gpc1_1 gpc189 (
      {stage0_1[179]},
      {stage1_1[62]}
   );
   gpc1_1 gpc190 (
      {stage0_1[180]},
      {stage1_1[63]}
   );
   gpc1_1 gpc191 (
      {stage0_1[181]},
      {stage1_1[64]}
   );
   gpc1_1 gpc192 (
      {stage0_1[182]},
      {stage1_1[65]}
   );
   gpc1_1 gpc193 (
      {stage0_1[183]},
      {stage1_1[66]}
   );
   gpc1_1 gpc194 (
      {stage0_1[184]},
      {stage1_1[67]}
   );
   gpc1_1 gpc195 (
      {stage0_1[185]},
      {stage1_1[68]}
   );
   gpc1_1 gpc196 (
      {stage0_1[186]},
      {stage1_1[69]}
   );
   gpc1_1 gpc197 (
      {stage0_1[187]},
      {stage1_1[70]}
   );
   gpc1_1 gpc198 (
      {stage0_1[188]},
      {stage1_1[71]}
   );
   gpc1_1 gpc199 (
      {stage0_2[173]},
      {stage1_2[58]}
   );
   gpc1_1 gpc200 (
      {stage0_2[174]},
      {stage1_2[59]}
   );
   gpc1_1 gpc201 (
      {stage0_2[175]},
      {stage1_2[60]}
   );
   gpc1_1 gpc202 (
      {stage0_2[176]},
      {stage1_2[61]}
   );
   gpc1_1 gpc203 (
      {stage0_2[177]},
      {stage1_2[62]}
   );
   gpc1_1 gpc204 (
      {stage0_2[178]},
      {stage1_2[63]}
   );
   gpc1_1 gpc205 (
      {stage0_2[179]},
      {stage1_2[64]}
   );
   gpc1_1 gpc206 (
      {stage0_2[180]},
      {stage1_2[65]}
   );
   gpc1_1 gpc207 (
      {stage0_2[181]},
      {stage1_2[66]}
   );
   gpc1_1 gpc208 (
      {stage0_2[182]},
      {stage1_2[67]}
   );
   gpc1_1 gpc209 (
      {stage0_2[183]},
      {stage1_2[68]}
   );
   gpc1_1 gpc210 (
      {stage0_2[184]},
      {stage1_2[69]}
   );
   gpc1_1 gpc211 (
      {stage0_2[185]},
      {stage1_2[70]}
   );
   gpc1_1 gpc212 (
      {stage0_2[186]},
      {stage1_2[71]}
   );
   gpc1_1 gpc213 (
      {stage0_2[187]},
      {stage1_2[72]}
   );
   gpc1_1 gpc214 (
      {stage0_2[188]},
      {stage1_2[73]}
   );
   gpc1_1 gpc215 (
      {stage0_6[180]},
      {stage1_6[62]}
   );
   gpc1_1 gpc216 (
      {stage0_6[181]},
      {stage1_6[63]}
   );
   gpc1_1 gpc217 (
      {stage0_6[182]},
      {stage1_6[64]}
   );
   gpc1_1 gpc218 (
      {stage0_6[183]},
      {stage1_6[65]}
   );
   gpc1_1 gpc219 (
      {stage0_6[184]},
      {stage1_6[66]}
   );
   gpc1_1 gpc220 (
      {stage0_6[185]},
      {stage1_6[67]}
   );
   gpc1_1 gpc221 (
      {stage0_6[186]},
      {stage1_6[68]}
   );
   gpc1_1 gpc222 (
      {stage0_6[187]},
      {stage1_6[69]}
   );
   gpc1_1 gpc223 (
      {stage0_6[188]},
      {stage1_6[70]}
   );
   gpc1_1 gpc224 (
      {stage0_7[179]},
      {stage1_7[68]}
   );
   gpc1_1 gpc225 (
      {stage0_7[180]},
      {stage1_7[69]}
   );
   gpc1_1 gpc226 (
      {stage0_7[181]},
      {stage1_7[70]}
   );
   gpc1_1 gpc227 (
      {stage0_7[182]},
      {stage1_7[71]}
   );
   gpc1_1 gpc228 (
      {stage0_7[183]},
      {stage1_7[72]}
   );
   gpc1_1 gpc229 (
      {stage0_7[184]},
      {stage1_7[73]}
   );
   gpc1_1 gpc230 (
      {stage0_7[185]},
      {stage1_7[74]}
   );
   gpc1_1 gpc231 (
      {stage0_7[186]},
      {stage1_7[75]}
   );
   gpc1_1 gpc232 (
      {stage0_7[187]},
      {stage1_7[76]}
   );
   gpc1_1 gpc233 (
      {stage0_7[188]},
      {stage1_7[77]}
   );
   gpc1_1 gpc234 (
      {stage0_8[183]},
      {stage1_8[91]}
   );
   gpc1_1 gpc235 (
      {stage0_8[184]},
      {stage1_8[92]}
   );
   gpc1_1 gpc236 (
      {stage0_8[185]},
      {stage1_8[93]}
   );
   gpc1_1 gpc237 (
      {stage0_8[186]},
      {stage1_8[94]}
   );
   gpc1_1 gpc238 (
      {stage0_8[187]},
      {stage1_8[95]}
   );
   gpc1_1 gpc239 (
      {stage0_8[188]},
      {stage1_8[96]}
   );
   gpc1_1 gpc240 (
      {stage0_9[183]},
      {stage1_9[84]}
   );
   gpc1_1 gpc241 (
      {stage0_9[184]},
      {stage1_9[85]}
   );
   gpc1_1 gpc242 (
      {stage0_9[185]},
      {stage1_9[86]}
   );
   gpc1_1 gpc243 (
      {stage0_9[186]},
      {stage1_9[87]}
   );
   gpc1_1 gpc244 (
      {stage0_9[187]},
      {stage1_9[88]}
   );
   gpc1_1 gpc245 (
      {stage0_9[188]},
      {stage1_9[89]}
   );
   gpc1_1 gpc246 (
      {stage0_10[181]},
      {stage1_10[60]}
   );
   gpc1_1 gpc247 (
      {stage0_10[182]},
      {stage1_10[61]}
   );
   gpc1_1 gpc248 (
      {stage0_10[183]},
      {stage1_10[62]}
   );
   gpc1_1 gpc249 (
      {stage0_10[184]},
      {stage1_10[63]}
   );
   gpc1_1 gpc250 (
      {stage0_10[185]},
      {stage1_10[64]}
   );
   gpc1_1 gpc251 (
      {stage0_10[186]},
      {stage1_10[65]}
   );
   gpc1_1 gpc252 (
      {stage0_10[187]},
      {stage1_10[66]}
   );
   gpc1_1 gpc253 (
      {stage0_10[188]},
      {stage1_10[67]}
   );
   gpc1_1 gpc254 (
      {stage0_11[138]},
      {stage1_11[60]}
   );
   gpc1_1 gpc255 (
      {stage0_11[139]},
      {stage1_11[61]}
   );
   gpc1_1 gpc256 (
      {stage0_11[140]},
      {stage1_11[62]}
   );
   gpc1_1 gpc257 (
      {stage0_11[141]},
      {stage1_11[63]}
   );
   gpc1_1 gpc258 (
      {stage0_11[142]},
      {stage1_11[64]}
   );
   gpc1_1 gpc259 (
      {stage0_11[143]},
      {stage1_11[65]}
   );
   gpc1_1 gpc260 (
      {stage0_11[144]},
      {stage1_11[66]}
   );
   gpc1_1 gpc261 (
      {stage0_11[145]},
      {stage1_11[67]}
   );
   gpc1_1 gpc262 (
      {stage0_11[146]},
      {stage1_11[68]}
   );
   gpc1_1 gpc263 (
      {stage0_11[147]},
      {stage1_11[69]}
   );
   gpc1_1 gpc264 (
      {stage0_11[148]},
      {stage1_11[70]}
   );
   gpc1_1 gpc265 (
      {stage0_11[149]},
      {stage1_11[71]}
   );
   gpc1_1 gpc266 (
      {stage0_11[150]},
      {stage1_11[72]}
   );
   gpc1_1 gpc267 (
      {stage0_11[151]},
      {stage1_11[73]}
   );
   gpc1_1 gpc268 (
      {stage0_11[152]},
      {stage1_11[74]}
   );
   gpc1_1 gpc269 (
      {stage0_11[153]},
      {stage1_11[75]}
   );
   gpc1_1 gpc270 (
      {stage0_11[154]},
      {stage1_11[76]}
   );
   gpc1_1 gpc271 (
      {stage0_11[155]},
      {stage1_11[77]}
   );
   gpc1_1 gpc272 (
      {stage0_11[156]},
      {stage1_11[78]}
   );
   gpc1_1 gpc273 (
      {stage0_11[157]},
      {stage1_11[79]}
   );
   gpc1_1 gpc274 (
      {stage0_11[158]},
      {stage1_11[80]}
   );
   gpc1_1 gpc275 (
      {stage0_11[159]},
      {stage1_11[81]}
   );
   gpc1_1 gpc276 (
      {stage0_11[160]},
      {stage1_11[82]}
   );
   gpc1_1 gpc277 (
      {stage0_11[161]},
      {stage1_11[83]}
   );
   gpc1_1 gpc278 (
      {stage0_11[162]},
      {stage1_11[84]}
   );
   gpc1_1 gpc279 (
      {stage0_11[163]},
      {stage1_11[85]}
   );
   gpc1_1 gpc280 (
      {stage0_11[164]},
      {stage1_11[86]}
   );
   gpc1_1 gpc281 (
      {stage0_11[165]},
      {stage1_11[87]}
   );
   gpc1_1 gpc282 (
      {stage0_11[166]},
      {stage1_11[88]}
   );
   gpc1_1 gpc283 (
      {stage0_11[167]},
      {stage1_11[89]}
   );
   gpc1_1 gpc284 (
      {stage0_11[168]},
      {stage1_11[90]}
   );
   gpc1_1 gpc285 (
      {stage0_11[169]},
      {stage1_11[91]}
   );
   gpc1_1 gpc286 (
      {stage0_11[170]},
      {stage1_11[92]}
   );
   gpc1_1 gpc287 (
      {stage0_11[171]},
      {stage1_11[93]}
   );
   gpc1_1 gpc288 (
      {stage0_11[172]},
      {stage1_11[94]}
   );
   gpc1_1 gpc289 (
      {stage0_11[173]},
      {stage1_11[95]}
   );
   gpc1_1 gpc290 (
      {stage0_11[174]},
      {stage1_11[96]}
   );
   gpc1_1 gpc291 (
      {stage0_11[175]},
      {stage1_11[97]}
   );
   gpc1_1 gpc292 (
      {stage0_11[176]},
      {stage1_11[98]}
   );
   gpc1_1 gpc293 (
      {stage0_11[177]},
      {stage1_11[99]}
   );
   gpc1_1 gpc294 (
      {stage0_11[178]},
      {stage1_11[100]}
   );
   gpc1_1 gpc295 (
      {stage0_11[179]},
      {stage1_11[101]}
   );
   gpc1_1 gpc296 (
      {stage0_11[180]},
      {stage1_11[102]}
   );
   gpc1_1 gpc297 (
      {stage0_11[181]},
      {stage1_11[103]}
   );
   gpc1_1 gpc298 (
      {stage0_11[182]},
      {stage1_11[104]}
   );
   gpc1_1 gpc299 (
      {stage0_11[183]},
      {stage1_11[105]}
   );
   gpc1_1 gpc300 (
      {stage0_11[184]},
      {stage1_11[106]}
   );
   gpc1_1 gpc301 (
      {stage0_11[185]},
      {stage1_11[107]}
   );
   gpc1_1 gpc302 (
      {stage0_11[186]},
      {stage1_11[108]}
   );
   gpc1_1 gpc303 (
      {stage0_11[187]},
      {stage1_11[109]}
   );
   gpc1_1 gpc304 (
      {stage0_11[188]},
      {stage1_11[110]}
   );
   gpc2135_5 gpc305 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc306 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc307 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc308 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc309 (
      {stage1_0[20], stage1_0[21], stage1_0[22]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[4]},
      {stage1_3[8]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc310 (
      {stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[5]},
      {stage1_3[9]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc311 (
      {stage1_0[26], stage1_0[27], stage1_0[28]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[6]},
      {stage1_3[10]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc312 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage2_5[0],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc313 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage2_5[1],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc314 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage2_5[2],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc606_5 gpc315 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34]},
      {stage2_5[3],stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10]}
   );
   gpc606_5 gpc316 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40]},
      {stage2_5[4],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc317 (
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[5],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc606_5 gpc318 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[6],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc606_5 gpc319 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[7],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc606_5 gpc320 (
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[8],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc606_5 gpc321 (
      {stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[9],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc606_5 gpc322 (
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[10],stage2_4[17],stage2_3[17],stage2_2[17]}
   );
   gpc606_5 gpc323 (
      {stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[11],stage2_4[18],stage2_3[18],stage2_2[18]}
   );
   gpc615_5 gpc324 (
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_3[41]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[12],stage2_4[19],stage2_3[19],stage2_2[19]}
   );
   gpc615_5 gpc325 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58]},
      {stage1_3[42]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[13],stage2_4[20],stage2_3[20],stage2_2[20]}
   );
   gpc615_5 gpc326 (
      {stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage1_3[43]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[14],stage2_4[21],stage2_3[21],stage2_2[21]}
   );
   gpc615_5 gpc327 (
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68]},
      {stage1_3[44]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[15],stage2_4[22],stage2_3[22],stage2_2[22]}
   );
   gpc615_5 gpc328 (
      {stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73]},
      {stage1_3[45]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[16],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc329 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[72]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[12],stage2_5[17],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc330 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[73]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[13],stage2_5[18],stage2_4[25],stage2_3[25]}
   );
   gpc615_5 gpc331 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[74]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[14],stage2_5[19],stage2_4[26],stage2_3[26]}
   );
   gpc606_5 gpc332 (
      {stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[15],stage2_5[20],stage2_4[27]}
   );
   gpc606_5 gpc333 (
      {stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[16],stage2_5[21],stage2_4[28]}
   );
   gpc606_5 gpc334 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[17],stage2_5[22],stage2_4[29]}
   );
   gpc606_5 gpc335 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[3],stage2_7[6],stage2_6[18],stage2_5[23]}
   );
   gpc606_5 gpc336 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[4],stage2_7[7],stage2_6[19],stage2_5[24]}
   );
   gpc606_5 gpc337 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[5],stage2_7[8],stage2_6[20],stage2_5[25]}
   );
   gpc606_5 gpc338 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[6],stage2_7[9],stage2_6[21],stage2_5[26]}
   );
   gpc606_5 gpc339 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[7],stage2_7[10],stage2_6[22],stage2_5[27]}
   );
   gpc606_5 gpc340 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[8],stage2_7[11],stage2_6[23],stage2_5[28]}
   );
   gpc606_5 gpc341 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[9],stage2_7[12],stage2_6[24],stage2_5[29]}
   );
   gpc606_5 gpc342 (
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[10],stage2_7[13],stage2_6[25],stage2_5[30]}
   );
   gpc606_5 gpc343 (
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[11],stage2_7[14],stage2_6[26],stage2_5[31]}
   );
   gpc606_5 gpc344 (
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[12],stage2_7[15],stage2_6[27],stage2_5[32]}
   );
   gpc606_5 gpc345 (
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[13],stage2_7[16],stage2_6[28],stage2_5[33]}
   );
   gpc606_5 gpc346 (
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[11],stage2_8[14],stage2_7[17],stage2_6[29]}
   );
   gpc606_5 gpc347 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[12],stage2_8[15],stage2_7[18],stage2_6[30]}
   );
   gpc606_5 gpc348 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[13],stage2_8[16],stage2_7[19],stage2_6[31]}
   );
   gpc615_5 gpc349 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[66]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[14],stage2_8[17],stage2_7[20],stage2_6[32]}
   );
   gpc615_5 gpc350 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[67]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[15],stage2_8[18],stage2_7[21],stage2_6[33]}
   );
   gpc615_5 gpc351 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[68]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[16],stage2_8[19],stage2_7[22],stage2_6[34]}
   );
   gpc615_5 gpc352 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[69]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[17],stage2_8[20],stage2_7[23],stage2_6[35]}
   );
   gpc615_5 gpc353 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[70]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[18],stage2_8[21],stage2_7[24],stage2_6[36]}
   );
   gpc615_5 gpc354 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[71]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[19],stage2_8[22],stage2_7[25],stage2_6[37]}
   );
   gpc615_5 gpc355 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[72]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[20],stage2_8[23],stage2_7[26],stage2_6[38]}
   );
   gpc615_5 gpc356 (
      {stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage1_8[60]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[10],stage2_9[21],stage2_8[24],stage2_7[27]}
   );
   gpc606_5 gpc357 (
      {stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[11],stage2_9[22],stage2_8[25]}
   );
   gpc606_5 gpc358 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[12],stage2_9[23],stage2_8[26]}
   );
   gpc606_5 gpc359 (
      {stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[13],stage2_9[24],stage2_8[27]}
   );
   gpc606_5 gpc360 (
      {stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[4],stage2_10[14],stage2_9[25],stage2_8[28]}
   );
   gpc606_5 gpc361 (
      {stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89], stage1_8[90]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[5],stage2_10[15],stage2_9[26],stage2_8[29]}
   );
   gpc606_5 gpc362 (
      {stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95], stage1_8[96]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[6],stage2_10[16],stage2_9[27],stage2_8[30]}
   );
   gpc606_5 gpc363 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[6],stage2_11[7],stage2_10[17],stage2_9[28]}
   );
   gpc606_5 gpc364 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[7],stage2_11[8],stage2_10[18],stage2_9[29]}
   );
   gpc606_5 gpc365 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[8],stage2_11[9],stage2_10[19],stage2_9[30]}
   );
   gpc606_5 gpc366 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[9],stage2_11[10],stage2_10[20],stage2_9[31]}
   );
   gpc606_5 gpc367 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[10],stage2_11[11],stage2_10[21],stage2_9[32]}
   );
   gpc606_5 gpc368 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[11],stage2_11[12],stage2_10[22],stage2_9[33]}
   );
   gpc606_5 gpc369 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[12],stage2_11[13],stage2_10[23],stage2_9[34]}
   );
   gpc606_5 gpc370 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[13],stage2_11[14],stage2_10[24],stage2_9[35]}
   );
   gpc606_5 gpc371 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[14],stage2_11[15],stage2_10[25],stage2_9[36]}
   );
   gpc606_5 gpc372 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[15],stage2_11[16],stage2_10[26],stage2_9[37]}
   );
   gpc606_5 gpc373 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[16],stage2_11[17],stage2_10[27],stage2_9[38]}
   );
   gpc606_5 gpc374 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[17],stage2_11[18],stage2_10[28],stage2_9[39]}
   );
   gpc606_5 gpc375 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[18],stage2_11[19],stage2_10[29],stage2_9[40]}
   );
   gpc606_5 gpc376 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[19],stage2_11[20],stage2_10[30],stage2_9[41]}
   );
   gpc606_5 gpc377 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[14],stage2_12[20],stage2_11[21],stage2_10[31]}
   );
   gpc606_5 gpc378 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[15],stage2_12[21],stage2_11[22],stage2_10[32]}
   );
   gpc606_5 gpc379 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[16],stage2_12[22],stage2_11[23],stage2_10[33]}
   );
   gpc606_5 gpc380 (
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[17],stage2_12[23],stage2_11[24],stage2_10[34]}
   );
   gpc606_5 gpc381 (
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[18],stage2_12[24],stage2_11[25],stage2_10[35]}
   );
   gpc615_5 gpc382 (
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88]},
      {stage1_12[30]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[19],stage2_12[25],stage2_11[26]}
   );
   gpc1_1 gpc383 (
      {stage1_0[29]},
      {stage2_0[7]}
   );
   gpc1_1 gpc384 (
      {stage1_0[30]},
      {stage2_0[8]}
   );
   gpc1_1 gpc385 (
      {stage1_0[31]},
      {stage2_0[9]}
   );
   gpc1_1 gpc386 (
      {stage1_0[32]},
      {stage2_0[10]}
   );
   gpc1_1 gpc387 (
      {stage1_0[33]},
      {stage2_0[11]}
   );
   gpc1_1 gpc388 (
      {stage1_0[34]},
      {stage2_0[12]}
   );
   gpc1_1 gpc389 (
      {stage1_0[35]},
      {stage2_0[13]}
   );
   gpc1_1 gpc390 (
      {stage1_0[36]},
      {stage2_0[14]}
   );
   gpc1_1 gpc391 (
      {stage1_0[37]},
      {stage2_0[15]}
   );
   gpc1_1 gpc392 (
      {stage1_1[60]},
      {stage2_1[12]}
   );
   gpc1_1 gpc393 (
      {stage1_1[61]},
      {stage2_1[13]}
   );
   gpc1_1 gpc394 (
      {stage1_1[62]},
      {stage2_1[14]}
   );
   gpc1_1 gpc395 (
      {stage1_1[63]},
      {stage2_1[15]}
   );
   gpc1_1 gpc396 (
      {stage1_1[64]},
      {stage2_1[16]}
   );
   gpc1_1 gpc397 (
      {stage1_1[65]},
      {stage2_1[17]}
   );
   gpc1_1 gpc398 (
      {stage1_1[66]},
      {stage2_1[18]}
   );
   gpc1_1 gpc399 (
      {stage1_1[67]},
      {stage2_1[19]}
   );
   gpc1_1 gpc400 (
      {stage1_1[68]},
      {stage2_1[20]}
   );
   gpc1_1 gpc401 (
      {stage1_1[69]},
      {stage2_1[21]}
   );
   gpc1_1 gpc402 (
      {stage1_1[70]},
      {stage2_1[22]}
   );
   gpc1_1 gpc403 (
      {stage1_1[71]},
      {stage2_1[23]}
   );
   gpc1_1 gpc404 (
      {stage1_3[61]},
      {stage2_3[27]}
   );
   gpc1_1 gpc405 (
      {stage1_3[62]},
      {stage2_3[28]}
   );
   gpc1_1 gpc406 (
      {stage1_3[63]},
      {stage2_3[29]}
   );
   gpc1_1 gpc407 (
      {stage1_3[64]},
      {stage2_3[30]}
   );
   gpc1_1 gpc408 (
      {stage1_4[93]},
      {stage2_4[30]}
   );
   gpc1_1 gpc409 (
      {stage1_4[94]},
      {stage2_4[31]}
   );
   gpc1_1 gpc410 (
      {stage1_5[84]},
      {stage2_5[34]}
   );
   gpc1_1 gpc411 (
      {stage1_5[85]},
      {stage2_5[35]}
   );
   gpc1_1 gpc412 (
      {stage1_10[66]},
      {stage2_10[36]}
   );
   gpc1_1 gpc413 (
      {stage1_10[67]},
      {stage2_10[37]}
   );
   gpc1_1 gpc414 (
      {stage1_11[89]},
      {stage2_11[27]}
   );
   gpc1_1 gpc415 (
      {stage1_11[90]},
      {stage2_11[28]}
   );
   gpc1_1 gpc416 (
      {stage1_11[91]},
      {stage2_11[29]}
   );
   gpc1_1 gpc417 (
      {stage1_11[92]},
      {stage2_11[30]}
   );
   gpc1_1 gpc418 (
      {stage1_11[93]},
      {stage2_11[31]}
   );
   gpc1_1 gpc419 (
      {stage1_11[94]},
      {stage2_11[32]}
   );
   gpc1_1 gpc420 (
      {stage1_11[95]},
      {stage2_11[33]}
   );
   gpc1_1 gpc421 (
      {stage1_11[96]},
      {stage2_11[34]}
   );
   gpc1_1 gpc422 (
      {stage1_11[97]},
      {stage2_11[35]}
   );
   gpc1_1 gpc423 (
      {stage1_11[98]},
      {stage2_11[36]}
   );
   gpc1_1 gpc424 (
      {stage1_11[99]},
      {stage2_11[37]}
   );
   gpc1_1 gpc425 (
      {stage1_11[100]},
      {stage2_11[38]}
   );
   gpc1_1 gpc426 (
      {stage1_11[101]},
      {stage2_11[39]}
   );
   gpc1_1 gpc427 (
      {stage1_11[102]},
      {stage2_11[40]}
   );
   gpc1_1 gpc428 (
      {stage1_11[103]},
      {stage2_11[41]}
   );
   gpc1_1 gpc429 (
      {stage1_11[104]},
      {stage2_11[42]}
   );
   gpc1_1 gpc430 (
      {stage1_11[105]},
      {stage2_11[43]}
   );
   gpc1_1 gpc431 (
      {stage1_11[106]},
      {stage2_11[44]}
   );
   gpc1_1 gpc432 (
      {stage1_11[107]},
      {stage2_11[45]}
   );
   gpc1_1 gpc433 (
      {stage1_11[108]},
      {stage2_11[46]}
   );
   gpc1_1 gpc434 (
      {stage1_11[109]},
      {stage2_11[47]}
   );
   gpc1_1 gpc435 (
      {stage1_11[110]},
      {stage2_11[48]}
   );
   gpc1_1 gpc436 (
      {stage1_12[31]},
      {stage2_12[26]}
   );
   gpc1_1 gpc437 (
      {stage1_12[32]},
      {stage2_12[27]}
   );
   gpc1_1 gpc438 (
      {stage1_12[33]},
      {stage2_12[28]}
   );
   gpc1_1 gpc439 (
      {stage1_12[34]},
      {stage2_12[29]}
   );
   gpc1_1 gpc440 (
      {stage1_12[35]},
      {stage2_12[30]}
   );
   gpc1_1 gpc441 (
      {stage1_12[36]},
      {stage2_12[31]}
   );
   gpc1_1 gpc442 (
      {stage1_12[37]},
      {stage2_12[32]}
   );
   gpc1_1 gpc443 (
      {stage1_12[38]},
      {stage2_12[33]}
   );
   gpc1_1 gpc444 (
      {stage1_12[39]},
      {stage2_12[34]}
   );
   gpc1_1 gpc445 (
      {stage1_12[40]},
      {stage2_12[35]}
   );
   gpc1_1 gpc446 (
      {stage1_12[41]},
      {stage2_12[36]}
   );
   gpc1_1 gpc447 (
      {stage1_12[42]},
      {stage2_12[37]}
   );
   gpc1_1 gpc448 (
      {stage1_12[43]},
      {stage2_12[38]}
   );
   gpc1_1 gpc449 (
      {stage1_12[44]},
      {stage2_12[39]}
   );
   gpc1_1 gpc450 (
      {stage1_12[45]},
      {stage2_12[40]}
   );
   gpc1_1 gpc451 (
      {stage1_12[46]},
      {stage2_12[41]}
   );
   gpc1_1 gpc452 (
      {stage1_12[47]},
      {stage2_12[42]}
   );
   gpc1_1 gpc453 (
      {stage1_12[48]},
      {stage2_12[43]}
   );
   gpc1_1 gpc454 (
      {stage1_12[49]},
      {stage2_12[44]}
   );
   gpc1_1 gpc455 (
      {stage1_12[50]},
      {stage2_12[45]}
   );
   gpc1_1 gpc456 (
      {stage1_12[51]},
      {stage2_12[46]}
   );
   gpc1_1 gpc457 (
      {stage1_12[52]},
      {stage2_12[47]}
   );
   gpc1_1 gpc458 (
      {stage1_13[6]},
      {stage2_13[20]}
   );
   gpc1_1 gpc459 (
      {stage1_13[7]},
      {stage2_13[21]}
   );
   gpc1_1 gpc460 (
      {stage1_13[8]},
      {stage2_13[22]}
   );
   gpc1_1 gpc461 (
      {stage1_13[9]},
      {stage2_13[23]}
   );
   gpc1_1 gpc462 (
      {stage1_13[10]},
      {stage2_13[24]}
   );
   gpc1_1 gpc463 (
      {stage1_13[11]},
      {stage2_13[25]}
   );
   gpc1_1 gpc464 (
      {stage1_13[12]},
      {stage2_13[26]}
   );
   gpc1_1 gpc465 (
      {stage1_13[13]},
      {stage2_13[27]}
   );
   gpc1_1 gpc466 (
      {stage1_13[14]},
      {stage2_13[28]}
   );
   gpc1_1 gpc467 (
      {stage1_13[15]},
      {stage2_13[29]}
   );
   gpc1_1 gpc468 (
      {stage1_13[16]},
      {stage2_13[30]}
   );
   gpc1_1 gpc469 (
      {stage1_13[17]},
      {stage2_13[31]}
   );
   gpc1_1 gpc470 (
      {stage1_13[18]},
      {stage2_13[32]}
   );
   gpc1_1 gpc471 (
      {stage1_13[19]},
      {stage2_13[33]}
   );
   gpc1_1 gpc472 (
      {stage1_13[20]},
      {stage2_13[34]}
   );
   gpc1_1 gpc473 (
      {stage1_13[21]},
      {stage2_13[35]}
   );
   gpc1_1 gpc474 (
      {stage1_13[22]},
      {stage2_13[36]}
   );
   gpc606_5 gpc475 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc476 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_1[0]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc477 (
      {stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc478 (
      {stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11], stage2_1[12]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc479 (
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc606_5 gpc480 (
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[3],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc481 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc615_5 gpc482 (
      {stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21]},
      {stage2_4[13]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[3],stage3_5[5],stage3_4[7],stage3_3[7]}
   );
   gpc615_5 gpc483 (
      {stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26]},
      {stage2_4[14]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[4],stage3_5[6],stage3_4[8],stage3_3[8]}
   );
   gpc606_5 gpc484 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[5],stage3_5[7],stage3_4[9]}
   );
   gpc615_5 gpc485 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[18]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[6],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc486 (
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30]},
      {stage2_5[19]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[7],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc487 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[8]}
   );
   gpc615_5 gpc488 (
      {stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27]},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[9]}
   );
   gpc615_5 gpc489 (
      {stage2_6[28], stage2_6[29], stage2_6[30], stage2_6[31], stage2_6[32]},
      {stage2_7[2]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[2],stage3_8[5],stage3_7[8],stage3_6[10]}
   );
   gpc615_5 gpc490 (
      {stage2_6[33], stage2_6[34], stage2_6[35], stage2_6[36], stage2_6[37]},
      {stage2_7[3]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[3],stage3_8[6],stage3_7[9],stage3_6[11]}
   );
   gpc615_5 gpc491 (
      {stage2_7[4], stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8]},
      {stage2_8[24]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[4],stage3_9[4],stage3_8[7],stage3_7[10]}
   );
   gpc615_5 gpc492 (
      {stage2_7[9], stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage2_8[25]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[5],stage3_9[5],stage3_8[8],stage3_7[11]}
   );
   gpc615_5 gpc493 (
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_8[26]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[6],stage3_9[6],stage3_8[9],stage3_7[12]}
   );
   gpc615_5 gpc494 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[27]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[7],stage3_9[7],stage3_8[10],stage3_7[13]}
   );
   gpc1163_5 gpc495 (
      {stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_10[0]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[4],stage3_10[8],stage3_9[8],stage3_8[11]}
   );
   gpc606_5 gpc496 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage3_13[0],stage3_12[1],stage3_11[5],stage3_10[9],stage3_9[9]}
   );
   gpc606_5 gpc497 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage3_13[1],stage3_12[2],stage3_11[6],stage3_10[10],stage3_9[10]}
   );
   gpc606_5 gpc498 (
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[2],stage3_12[3],stage3_11[7],stage3_10[11]}
   );
   gpc606_5 gpc499 (
      {stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[3],stage3_12[4],stage3_11[8],stage3_10[12]}
   );
   gpc606_5 gpc500 (
      {stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[4],stage3_12[5],stage3_11[9],stage3_10[13]}
   );
   gpc606_5 gpc501 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[5],stage3_12[6],stage3_11[10],stage3_10[14]}
   );
   gpc606_5 gpc502 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[6],stage3_12[7],stage3_11[11],stage3_10[15]}
   );
   gpc606_5 gpc503 (
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[5],stage3_13[7],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc504 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[6],stage3_13[8],stage3_12[9],stage3_11[13]}
   );
   gpc606_5 gpc505 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[7],stage3_13[9],stage3_12[10],stage3_11[14]}
   );
   gpc606_5 gpc506 (
      {stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[8],stage3_13[10],stage3_12[11],stage3_11[15]}
   );
   gpc606_5 gpc507 (
      {stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[9],stage3_13[11],stage3_12[12],stage3_11[16]}
   );
   gpc606_5 gpc508 (
      {stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[10],stage3_13[12],stage3_12[13],stage3_11[17]}
   );
   gpc606_5 gpc509 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[6],stage3_14[11],stage3_13[13],stage3_12[14]}
   );
   gpc1_1 gpc510 (
      {stage2_0[11]},
      {stage3_0[2]}
   );
   gpc1_1 gpc511 (
      {stage2_0[12]},
      {stage3_0[3]}
   );
   gpc1_1 gpc512 (
      {stage2_0[13]},
      {stage3_0[4]}
   );
   gpc1_1 gpc513 (
      {stage2_0[14]},
      {stage3_0[5]}
   );
   gpc1_1 gpc514 (
      {stage2_0[15]},
      {stage3_0[6]}
   );
   gpc1_1 gpc515 (
      {stage2_1[13]},
      {stage3_1[4]}
   );
   gpc1_1 gpc516 (
      {stage2_1[14]},
      {stage3_1[5]}
   );
   gpc1_1 gpc517 (
      {stage2_1[15]},
      {stage3_1[6]}
   );
   gpc1_1 gpc518 (
      {stage2_1[16]},
      {stage3_1[7]}
   );
   gpc1_1 gpc519 (
      {stage2_1[17]},
      {stage3_1[8]}
   );
   gpc1_1 gpc520 (
      {stage2_1[18]},
      {stage3_1[9]}
   );
   gpc1_1 gpc521 (
      {stage2_1[19]},
      {stage3_1[10]}
   );
   gpc1_1 gpc522 (
      {stage2_1[20]},
      {stage3_1[11]}
   );
   gpc1_1 gpc523 (
      {stage2_1[21]},
      {stage3_1[12]}
   );
   gpc1_1 gpc524 (
      {stage2_1[22]},
      {stage3_1[13]}
   );
   gpc1_1 gpc525 (
      {stage2_1[23]},
      {stage3_1[14]}
   );
   gpc1_1 gpc526 (
      {stage2_3[27]},
      {stage3_3[9]}
   );
   gpc1_1 gpc527 (
      {stage2_3[28]},
      {stage3_3[10]}
   );
   gpc1_1 gpc528 (
      {stage2_3[29]},
      {stage3_3[11]}
   );
   gpc1_1 gpc529 (
      {stage2_3[30]},
      {stage3_3[12]}
   );
   gpc1_1 gpc530 (
      {stage2_4[31]},
      {stage3_4[12]}
   );
   gpc1_1 gpc531 (
      {stage2_5[20]},
      {stage3_5[10]}
   );
   gpc1_1 gpc532 (
      {stage2_5[21]},
      {stage3_5[11]}
   );
   gpc1_1 gpc533 (
      {stage2_5[22]},
      {stage3_5[12]}
   );
   gpc1_1 gpc534 (
      {stage2_5[23]},
      {stage3_5[13]}
   );
   gpc1_1 gpc535 (
      {stage2_5[24]},
      {stage3_5[14]}
   );
   gpc1_1 gpc536 (
      {stage2_5[25]},
      {stage3_5[15]}
   );
   gpc1_1 gpc537 (
      {stage2_5[26]},
      {stage3_5[16]}
   );
   gpc1_1 gpc538 (
      {stage2_5[27]},
      {stage3_5[17]}
   );
   gpc1_1 gpc539 (
      {stage2_5[28]},
      {stage3_5[18]}
   );
   gpc1_1 gpc540 (
      {stage2_5[29]},
      {stage3_5[19]}
   );
   gpc1_1 gpc541 (
      {stage2_5[30]},
      {stage3_5[20]}
   );
   gpc1_1 gpc542 (
      {stage2_5[31]},
      {stage3_5[21]}
   );
   gpc1_1 gpc543 (
      {stage2_5[32]},
      {stage3_5[22]}
   );
   gpc1_1 gpc544 (
      {stage2_5[33]},
      {stage3_5[23]}
   );
   gpc1_1 gpc545 (
      {stage2_5[34]},
      {stage3_5[24]}
   );
   gpc1_1 gpc546 (
      {stage2_5[35]},
      {stage3_5[25]}
   );
   gpc1_1 gpc547 (
      {stage2_6[38]},
      {stage3_6[12]}
   );
   gpc1_1 gpc548 (
      {stage2_7[24]},
      {stage3_7[14]}
   );
   gpc1_1 gpc549 (
      {stage2_7[25]},
      {stage3_7[15]}
   );
   gpc1_1 gpc550 (
      {stage2_7[26]},
      {stage3_7[16]}
   );
   gpc1_1 gpc551 (
      {stage2_7[27]},
      {stage3_7[17]}
   );
   gpc1_1 gpc552 (
      {stage2_10[31]},
      {stage3_10[16]}
   );
   gpc1_1 gpc553 (
      {stage2_10[32]},
      {stage3_10[17]}
   );
   gpc1_1 gpc554 (
      {stage2_10[33]},
      {stage3_10[18]}
   );
   gpc1_1 gpc555 (
      {stage2_10[34]},
      {stage3_10[19]}
   );
   gpc1_1 gpc556 (
      {stage2_10[35]},
      {stage3_10[20]}
   );
   gpc1_1 gpc557 (
      {stage2_10[36]},
      {stage3_10[21]}
   );
   gpc1_1 gpc558 (
      {stage2_10[37]},
      {stage3_10[22]}
   );
   gpc1_1 gpc559 (
      {stage2_12[36]},
      {stage3_12[15]}
   );
   gpc1_1 gpc560 (
      {stage2_12[37]},
      {stage3_12[16]}
   );
   gpc1_1 gpc561 (
      {stage2_12[38]},
      {stage3_12[17]}
   );
   gpc1_1 gpc562 (
      {stage2_12[39]},
      {stage3_12[18]}
   );
   gpc1_1 gpc563 (
      {stage2_12[40]},
      {stage3_12[19]}
   );
   gpc1_1 gpc564 (
      {stage2_12[41]},
      {stage3_12[20]}
   );
   gpc1_1 gpc565 (
      {stage2_12[42]},
      {stage3_12[21]}
   );
   gpc1_1 gpc566 (
      {stage2_12[43]},
      {stage3_12[22]}
   );
   gpc1_1 gpc567 (
      {stage2_12[44]},
      {stage3_12[23]}
   );
   gpc1_1 gpc568 (
      {stage2_12[45]},
      {stage3_12[24]}
   );
   gpc1_1 gpc569 (
      {stage2_12[46]},
      {stage3_12[25]}
   );
   gpc1_1 gpc570 (
      {stage2_12[47]},
      {stage3_12[26]}
   );
   gpc1_1 gpc571 (
      {stage2_13[36]},
      {stage3_13[14]}
   );
   gpc1_1 gpc572 (
      {stage2_15[0]},
      {stage3_15[7]}
   );
   gpc606_5 gpc573 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc574 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc575 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc576 (
      {stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc577 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc606_5 gpc578 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[2],stage4_7[3],stage4_6[3],stage4_5[4]}
   );
   gpc606_5 gpc579 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[3],stage4_7[4],stage4_6[4],stage4_5[5]}
   );
   gpc615_5 gpc580 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22]},
      {stage3_6[12]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[4],stage4_7[5],stage4_6[5],stage4_5[6]}
   );
   gpc606_5 gpc581 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[3],stage4_8[5]}
   );
   gpc606_5 gpc582 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[4],stage4_8[6]}
   );
   gpc615_5 gpc583 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[12]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[5]}
   );
   gpc615_5 gpc584 (
      {stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage3_11[6]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[1],stage4_12[3],stage4_11[3],stage4_10[3]}
   );
   gpc615_5 gpc585 (
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22]},
      {stage3_11[7]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[2],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc606_5 gpc586 (
      {stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12], stage3_11[13]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[2],stage4_13[3],stage4_12[5],stage4_11[5]}
   );
   gpc615_5 gpc587 (
      {stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17], 1'b0},
      {stage3_12[12]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[3],stage4_13[4],stage4_12[6],stage4_11[6]}
   );
   gpc606_5 gpc588 (
      {stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[4],stage4_13[5],stage4_12[7]}
   );
   gpc606_5 gpc589 (
      {stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23], stage3_12[24]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[5],stage4_13[6],stage4_12[8]}
   );
   gpc1_1 gpc590 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc591 (
      {stage3_1[6]},
      {stage4_1[2]}
   );
   gpc1_1 gpc592 (
      {stage3_1[7]},
      {stage4_1[3]}
   );
   gpc1_1 gpc593 (
      {stage3_1[8]},
      {stage4_1[4]}
   );
   gpc1_1 gpc594 (
      {stage3_1[9]},
      {stage4_1[5]}
   );
   gpc1_1 gpc595 (
      {stage3_1[10]},
      {stage4_1[6]}
   );
   gpc1_1 gpc596 (
      {stage3_1[11]},
      {stage4_1[7]}
   );
   gpc1_1 gpc597 (
      {stage3_1[12]},
      {stage4_1[8]}
   );
   gpc1_1 gpc598 (
      {stage3_1[13]},
      {stage4_1[9]}
   );
   gpc1_1 gpc599 (
      {stage3_1[14]},
      {stage4_1[10]}
   );
   gpc1_1 gpc600 (
      {stage3_3[11]},
      {stage4_3[3]}
   );
   gpc1_1 gpc601 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc602 (
      {stage3_5[23]},
      {stage4_5[7]}
   );
   gpc1_1 gpc603 (
      {stage3_5[24]},
      {stage4_5[8]}
   );
   gpc1_1 gpc604 (
      {stage3_5[25]},
      {stage4_5[9]}
   );
   gpc1_1 gpc605 (
      {stage3_9[5]},
      {stage4_9[6]}
   );
   gpc1_1 gpc606 (
      {stage3_9[6]},
      {stage4_9[7]}
   );
   gpc1_1 gpc607 (
      {stage3_9[7]},
      {stage4_9[8]}
   );
   gpc1_1 gpc608 (
      {stage3_9[8]},
      {stage4_9[9]}
   );
   gpc1_1 gpc609 (
      {stage3_9[9]},
      {stage4_9[10]}
   );
   gpc1_1 gpc610 (
      {stage3_9[10]},
      {stage4_9[11]}
   );
   gpc1_1 gpc611 (
      {stage3_12[25]},
      {stage4_12[9]}
   );
   gpc1_1 gpc612 (
      {stage3_12[26]},
      {stage4_12[10]}
   );
   gpc1_1 gpc613 (
      {stage3_13[12]},
      {stage4_13[7]}
   );
   gpc1_1 gpc614 (
      {stage3_13[13]},
      {stage4_13[8]}
   );
   gpc1_1 gpc615 (
      {stage3_13[14]},
      {stage4_13[9]}
   );
   gpc1_1 gpc616 (
      {stage3_15[0]},
      {stage4_15[4]}
   );
   gpc1_1 gpc617 (
      {stage3_15[1]},
      {stage4_15[5]}
   );
   gpc1_1 gpc618 (
      {stage3_15[2]},
      {stage4_15[6]}
   );
   gpc1_1 gpc619 (
      {stage3_15[3]},
      {stage4_15[7]}
   );
   gpc1_1 gpc620 (
      {stage3_15[4]},
      {stage4_15[8]}
   );
   gpc1_1 gpc621 (
      {stage3_15[5]},
      {stage4_15[9]}
   );
   gpc1_1 gpc622 (
      {stage3_15[6]},
      {stage4_15[10]}
   );
   gpc1_1 gpc623 (
      {stage3_15[7]},
      {stage4_15[11]}
   );
   gpc1_1 gpc624 (
      {stage3_16[0]},
      {stage4_16[2]}
   );
   gpc1415_5 gpc625 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc2116_5 gpc626 (
      {stage4_1[5], stage4_1[6], stage4_1[7], stage4_1[8], stage4_1[9], stage4_1[10]},
      {stage4_2[1]},
      {stage4_3[4]},
      {stage4_4[1], stage4_4[2]},
      {stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc627 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[2]}
   );
   gpc606_5 gpc628 (
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc2135_5 gpc629 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[2]}
   );
   gpc606_5 gpc630 (
      {stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10]},
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2],stage5_9[3]}
   );
   gpc606_5 gpc631 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[2],stage5_12[2]}
   );
   gpc606_5 gpc632 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1],stage5_13[3]}
   );
   gpc606_5 gpc633 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], 1'b0, 1'b0},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[2],stage5_15[2],stage5_14[2],stage5_13[4]}
   );
   gpc1_1 gpc634 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc635 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc636 (
      {stage4_4[3]},
      {stage5_4[2]}
   );
   gpc1_1 gpc637 (
      {stage4_4[4]},
      {stage5_4[3]}
   );
   gpc1_1 gpc638 (
      {stage4_5[6]},
      {stage5_5[3]}
   );
   gpc1_1 gpc639 (
      {stage4_5[7]},
      {stage5_5[4]}
   );
   gpc1_1 gpc640 (
      {stage4_5[8]},
      {stage5_5[5]}
   );
   gpc1_1 gpc641 (
      {stage4_5[9]},
      {stage5_5[6]}
   );
   gpc1_1 gpc642 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc643 (
      {stage4_9[11]},
      {stage5_9[4]}
   );
   gpc1_1 gpc644 (
      {stage4_10[3]},
      {stage5_10[3]}
   );
   gpc1_1 gpc645 (
      {stage4_10[4]},
      {stage5_10[4]}
   );
   gpc1_1 gpc646 (
      {stage4_12[8]},
      {stage5_12[3]}
   );
   gpc1_1 gpc647 (
      {stage4_12[9]},
      {stage5_12[4]}
   );
   gpc1_1 gpc648 (
      {stage4_12[10]},
      {stage5_12[5]}
   );
   gpc1_1 gpc649 (
      {stage4_16[0]},
      {stage5_16[3]}
   );
   gpc1_1 gpc650 (
      {stage4_16[1]},
      {stage5_16[4]}
   );
   gpc1_1 gpc651 (
      {stage4_16[2]},
      {stage5_16[5]}
   );
   gpc1163_5 gpc652 (
      {stage5_4[0], stage5_4[1], stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage5_6[0]},
      {stage5_7[0]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0]}
   );
   gpc1163_5 gpc653 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], 1'b0},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc615_5 gpc654 (
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], 1'b0},
      {stage5_11[1]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1],stage6_10[1]}
   );
   gpc135_4 gpc655 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4]},
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1163_5 gpc656 (
      {stage5_15[1], stage5_15[2], 1'b0},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[0]},
      {1'b0},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1]}
   );
   gpc1_1 gpc657 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc658 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc659 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc660 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc661 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc662 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc663 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc664 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc665 (
      {stage5_4[3]},
      {stage6_4[1]}
   );
   gpc1_1 gpc666 (
      {stage5_5[6]},
      {stage6_5[1]}
   );
   gpc1_1 gpc667 (
      {stage5_6[1]},
      {stage6_6[1]}
   );
   gpc1_1 gpc668 (
      {stage5_7[1]},
      {stage6_7[1]}
   );
   gpc1_1 gpc669 (
      {stage5_17[1]},
      {stage6_17[1]}
   );
endmodule
module rowadder2_1_20(input [19:0] src0, input [19:0] src1, output [20:0] dst0);
    wire [19:0] gene;
    wire [19:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    assign dst0 = {carryout[19], out[19:0]};
endmodule


module comp2_1test_189_12_189_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    reg [11:0] src128;
    reg [11:0] src129;
    reg [11:0] src130;
    reg [11:0] src131;
    reg [11:0] src132;
    reg [11:0] src133;
    reg [11:0] src134;
    reg [11:0] src135;
    reg [11:0] src136;
    reg [11:0] src137;
    reg [11:0] src138;
    reg [11:0] src139;
    reg [11:0] src140;
    reg [11:0] src141;
    reg [11:0] src142;
    reg [11:0] src143;
    reg [11:0] src144;
    reg [11:0] src145;
    reg [11:0] src146;
    reg [11:0] src147;
    reg [11:0] src148;
    reg [11:0] src149;
    reg [11:0] src150;
    reg [11:0] src151;
    reg [11:0] src152;
    reg [11:0] src153;
    reg [11:0] src154;
    reg [11:0] src155;
    reg [11:0] src156;
    reg [11:0] src157;
    reg [11:0] src158;
    reg [11:0] src159;
    reg [11:0] src160;
    reg [11:0] src161;
    reg [11:0] src162;
    reg [11:0] src163;
    reg [11:0] src164;
    reg [11:0] src165;
    reg [11:0] src166;
    reg [11:0] src167;
    reg [11:0] src168;
    reg [11:0] src169;
    reg [11:0] src170;
    reg [11:0] src171;
    reg [11:0] src172;
    reg [11:0] src173;
    reg [11:0] src174;
    reg [11:0] src175;
    reg [11:0] src176;
    reg [11:0] src177;
    reg [11:0] src178;
    reg [11:0] src179;
    reg [11:0] src180;
    reg [11:0] src181;
    reg [11:0] src182;
    reg [11:0] src183;
    reg [11:0] src184;
    reg [11:0] src185;
    reg [11:0] src186;
    reg [11:0] src187;
    reg [11:0] src188;
    reg [19:0] exp;
    wire [19:0] dst;
    assign test = dst == exp;
    compressor2_1_189_12 compressor2_1_189_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .src128(src128),
        .src129(src129),
        .src130(src130),
        .src131(src131),
        .src132(src132),
        .src133(src133),
        .src134(src134),
        .src135(src135),
        .src136(src136),
        .src137(src137),
        .src138(src138),
        .src139(src139),
        .src140(src140),
        .src141(src141),
        .src142(src142),
        .src143(src143),
        .src144(src144),
        .src145(src145),
        .src146(src146),
        .src147(src147),
        .src148(src148),
        .src149(src149),
        .src150(src150),
        .src151(src151),
        .src152(src152),
        .src153(src153),
        .src154(src154),
        .src155(src155),
        .src156(src156),
        .src157(src157),
        .src158(src158),
        .src159(src159),
        .src160(src160),
        .src161(src161),
        .src162(src162),
        .src163(src163),
        .src164(src164),
        .src165(src165),
        .src166(src166),
        .src167(src167),
        .src168(src168),
        .src169(src169),
        .src170(src170),
        .src171(src171),
        .src172(src172),
        .src173(src173),
        .src174(src174),
        .src175(src175),
        .src176(src176),
        .src177(src177),
        .src178(src178),
        .src179(src179),
        .src180(src180),
        .src181(src181),
        .src182(src182),
        .src183(src183),
        .src184(src184),
        .src185(src185),
        .src186(src186),
        .src187(src187),
        .src188(src188),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, src128, src129, src130, src131, src132, src133, src134, src135, src136, src137, src138, src139, src140, src141, src142, src143, src144, src145, src146, src147, src148, src149, src150, src151, src152, src153, src154, src155, src156, src157, src158, src159, src160, src161, src162, src163, src164, src165, src166, src167, src168, src169, src170, src171, src172, src173, src174, src175, src176, src177, src178, src179, src180, src181, src182, src183, src184, src185, src186, src187, src188, dst, exp, test);
        src0 <= 12'h589;
        src1 <= 12'h75c;
        src2 <= 12'h81c;
        src3 <= 12'hc59;
        src4 <= 12'hcbb;
        src5 <= 12'h302;
        src6 <= 12'h7db;
        src7 <= 12'hfe3;
        src8 <= 12'hfac;
        src9 <= 12'h1f5;
        src10 <= 12'hc78;
        src11 <= 12'haf0;
        src12 <= 12'h852;
        src13 <= 12'h3a8;
        src14 <= 12'h395;
        src15 <= 12'h354;
        src16 <= 12'hd0b;
        src17 <= 12'h1c5;
        src18 <= 12'hda9;
        src19 <= 12'hf34;
        src20 <= 12'h1c2;
        src21 <= 12'h186;
        src22 <= 12'h39c;
        src23 <= 12'h7f9;
        src24 <= 12'hd38;
        src25 <= 12'h8bc;
        src26 <= 12'hc54;
        src27 <= 12'h320;
        src28 <= 12'h674;
        src29 <= 12'had7;
        src30 <= 12'hdea;
        src31 <= 12'h59c;
        src32 <= 12'hc97;
        src33 <= 12'hdca;
        src34 <= 12'h2cd;
        src35 <= 12'hc45;
        src36 <= 12'hd2b;
        src37 <= 12'hc66;
        src38 <= 12'he25;
        src39 <= 12'h364;
        src40 <= 12'h4b3;
        src41 <= 12'h184;
        src42 <= 12'h129;
        src43 <= 12'h926;
        src44 <= 12'h7b9;
        src45 <= 12'h777;
        src46 <= 12'h392;
        src47 <= 12'hea;
        src48 <= 12'hf9;
        src49 <= 12'h135;
        src50 <= 12'h5ce;
        src51 <= 12'hd09;
        src52 <= 12'he3c;
        src53 <= 12'h869;
        src54 <= 12'h39a;
        src55 <= 12'h8ee;
        src56 <= 12'h9d2;
        src57 <= 12'hfd9;
        src58 <= 12'he3f;
        src59 <= 12'hded;
        src60 <= 12'hc9;
        src61 <= 12'hffa;
        src62 <= 12'hdfd;
        src63 <= 12'h3bb;
        src64 <= 12'h337;
        src65 <= 12'h928;
        src66 <= 12'hdb;
        src67 <= 12'h1a1;
        src68 <= 12'h925;
        src69 <= 12'hda7;
        src70 <= 12'h8f6;
        src71 <= 12'h494;
        src72 <= 12'h9cd;
        src73 <= 12'hc2d;
        src74 <= 12'h947;
        src75 <= 12'h4fe;
        src76 <= 12'h9fd;
        src77 <= 12'h7d;
        src78 <= 12'hee7;
        src79 <= 12'h9c8;
        src80 <= 12'hf5e;
        src81 <= 12'h3d2;
        src82 <= 12'h7e1;
        src83 <= 12'h270;
        src84 <= 12'h808;
        src85 <= 12'h5b0;
        src86 <= 12'ha5a;
        src87 <= 12'h157;
        src88 <= 12'h272;
        src89 <= 12'h78c;
        src90 <= 12'hc66;
        src91 <= 12'h811;
        src92 <= 12'h124;
        src93 <= 12'h17;
        src94 <= 12'h83c;
        src95 <= 12'hc9c;
        src96 <= 12'hb37;
        src97 <= 12'hcd;
        src98 <= 12'h1a;
        src99 <= 12'h65b;
        src100 <= 12'h875;
        src101 <= 12'h77c;
        src102 <= 12'h3eb;
        src103 <= 12'h649;
        src104 <= 12'h99c;
        src105 <= 12'h814;
        src106 <= 12'he84;
        src107 <= 12'h377;
        src108 <= 12'h8f6;
        src109 <= 12'h7a6;
        src110 <= 12'h851;
        src111 <= 12'h6c8;
        src112 <= 12'h459;
        src113 <= 12'h6d2;
        src114 <= 12'h282;
        src115 <= 12'h64a;
        src116 <= 12'h284;
        src117 <= 12'h391;
        src118 <= 12'h126;
        src119 <= 12'hb7f;
        src120 <= 12'h9ba;
        src121 <= 12'h335;
        src122 <= 12'hc07;
        src123 <= 12'hb1f;
        src124 <= 12'hf10;
        src125 <= 12'h34c;
        src126 <= 12'h91f;
        src127 <= 12'h459;
        src128 <= 12'h400;
        src129 <= 12'h85e;
        src130 <= 12'h672;
        src131 <= 12'h45a;
        src132 <= 12'h8cd;
        src133 <= 12'hefd;
        src134 <= 12'hd03;
        src135 <= 12'hb59;
        src136 <= 12'h2b6;
        src137 <= 12'h9fd;
        src138 <= 12'he21;
        src139 <= 12'hb42;
        src140 <= 12'h459;
        src141 <= 12'h27a;
        src142 <= 12'h437;
        src143 <= 12'h469;
        src144 <= 12'hed7;
        src145 <= 12'hd;
        src146 <= 12'h6cb;
        src147 <= 12'hd52;
        src148 <= 12'h9;
        src149 <= 12'h3ff;
        src150 <= 12'h35e;
        src151 <= 12'h340;
        src152 <= 12'h89;
        src153 <= 12'h741;
        src154 <= 12'hb1e;
        src155 <= 12'h517;
        src156 <= 12'h214;
        src157 <= 12'ha99;
        src158 <= 12'h303;
        src159 <= 12'hed7;
        src160 <= 12'ha1b;
        src161 <= 12'h25c;
        src162 <= 12'hfa9;
        src163 <= 12'hf95;
        src164 <= 12'h3b7;
        src165 <= 12'hcd7;
        src166 <= 12'h755;
        src167 <= 12'h67f;
        src168 <= 12'h1b5;
        src169 <= 12'h89c;
        src170 <= 12'hf26;
        src171 <= 12'hb05;
        src172 <= 12'ha5a;
        src173 <= 12'h481;
        src174 <= 12'ha44;
        src175 <= 12'h3e1;
        src176 <= 12'hb14;
        src177 <= 12'h47f;
        src178 <= 12'hc4d;
        src179 <= 12'h903;
        src180 <= 12'h4c9;
        src181 <= 12'h91e;
        src182 <= 12'h87c;
        src183 <= 12'hc98;
        src184 <= 12'h3df;
        src185 <= 12'hdf2;
        src186 <= 12'hf41;
        src187 <= 12'h313;
        src188 <= 12'hdff;
        exp <= 20'h5ba05;
        #1
        src0 <= 12'h25;
        src1 <= 12'h41a;
        src2 <= 12'hf7c;
        src3 <= 12'had4;
        src4 <= 12'h3d8;
        src5 <= 12'h95c;
        src6 <= 12'ha6;
        src7 <= 12'hfe3;
        src8 <= 12'hb86;
        src9 <= 12'hcb1;
        src10 <= 12'h63d;
        src11 <= 12'hafe;
        src12 <= 12'h3f4;
        src13 <= 12'h374;
        src14 <= 12'h5c0;
        src15 <= 12'ha7;
        src16 <= 12'h58e;
        src17 <= 12'h6d4;
        src18 <= 12'h23d;
        src19 <= 12'h138;
        src20 <= 12'haac;
        src21 <= 12'hb04;
        src22 <= 12'hf64;
        src23 <= 12'h756;
        src24 <= 12'h293;
        src25 <= 12'h991;
        src26 <= 12'h2d2;
        src27 <= 12'ha9c;
        src28 <= 12'h737;
        src29 <= 12'h1ec;
        src30 <= 12'h15d;
        src31 <= 12'h890;
        src32 <= 12'h8f7;
        src33 <= 12'h94a;
        src34 <= 12'h990;
        src35 <= 12'h499;
        src36 <= 12'hfef;
        src37 <= 12'h5e8;
        src38 <= 12'h104;
        src39 <= 12'h5c4;
        src40 <= 12'hfbb;
        src41 <= 12'he7a;
        src42 <= 12'he6b;
        src43 <= 12'h6dc;
        src44 <= 12'hb1d;
        src45 <= 12'hb18;
        src46 <= 12'h894;
        src47 <= 12'hdf2;
        src48 <= 12'ha6;
        src49 <= 12'hfb1;
        src50 <= 12'hf91;
        src51 <= 12'h9a8;
        src52 <= 12'hbe6;
        src53 <= 12'hb1f;
        src54 <= 12'h4e8;
        src55 <= 12'hc85;
        src56 <= 12'h45e;
        src57 <= 12'h33a;
        src58 <= 12'h594;
        src59 <= 12'h7d7;
        src60 <= 12'hcf4;
        src61 <= 12'h98a;
        src62 <= 12'h433;
        src63 <= 12'h69e;
        src64 <= 12'h81;
        src65 <= 12'h7c3;
        src66 <= 12'hb2e;
        src67 <= 12'h66;
        src68 <= 12'hb69;
        src69 <= 12'hc56;
        src70 <= 12'h905;
        src71 <= 12'haf1;
        src72 <= 12'hbc1;
        src73 <= 12'hd86;
        src74 <= 12'h923;
        src75 <= 12'hd63;
        src76 <= 12'h1c2;
        src77 <= 12'h61d;
        src78 <= 12'haff;
        src79 <= 12'h636;
        src80 <= 12'h653;
        src81 <= 12'h32b;
        src82 <= 12'h564;
        src83 <= 12'h663;
        src84 <= 12'he93;
        src85 <= 12'h46f;
        src86 <= 12'hfae;
        src87 <= 12'h8dd;
        src88 <= 12'hd4c;
        src89 <= 12'h25b;
        src90 <= 12'h694;
        src91 <= 12'h901;
        src92 <= 12'hd65;
        src93 <= 12'had9;
        src94 <= 12'hc82;
        src95 <= 12'h593;
        src96 <= 12'hd2f;
        src97 <= 12'hff8;
        src98 <= 12'h2e0;
        src99 <= 12'hb7f;
        src100 <= 12'h867;
        src101 <= 12'h74f;
        src102 <= 12'h58b;
        src103 <= 12'h245;
        src104 <= 12'had1;
        src105 <= 12'h93a;
        src106 <= 12'haa;
        src107 <= 12'he79;
        src108 <= 12'h80d;
        src109 <= 12'hc99;
        src110 <= 12'hbe1;
        src111 <= 12'h74d;
        src112 <= 12'hce2;
        src113 <= 12'h35b;
        src114 <= 12'he2f;
        src115 <= 12'hedb;
        src116 <= 12'haf2;
        src117 <= 12'h27c;
        src118 <= 12'h8ed;
        src119 <= 12'hac2;
        src120 <= 12'h70e;
        src121 <= 12'h28a;
        src122 <= 12'h1cb;
        src123 <= 12'h890;
        src124 <= 12'ha4;
        src125 <= 12'hb9a;
        src126 <= 12'h8ad;
        src127 <= 12'hd14;
        src128 <= 12'h2dd;
        src129 <= 12'ha06;
        src130 <= 12'h254;
        src131 <= 12'hce7;
        src132 <= 12'h931;
        src133 <= 12'he22;
        src134 <= 12'h64d;
        src135 <= 12'h975;
        src136 <= 12'hb04;
        src137 <= 12'hb1c;
        src138 <= 12'h258;
        src139 <= 12'h9f9;
        src140 <= 12'he94;
        src141 <= 12'h5a;
        src142 <= 12'h78a;
        src143 <= 12'hb9c;
        src144 <= 12'h4bd;
        src145 <= 12'h5b2;
        src146 <= 12'h869;
        src147 <= 12'h9de;
        src148 <= 12'hf87;
        src149 <= 12'h9b1;
        src150 <= 12'hcf9;
        src151 <= 12'h883;
        src152 <= 12'hdab;
        src153 <= 12'hbad;
        src154 <= 12'h49e;
        src155 <= 12'hc5f;
        src156 <= 12'h848;
        src157 <= 12'h40d;
        src158 <= 12'h6e8;
        src159 <= 12'h961;
        src160 <= 12'hddb;
        src161 <= 12'h167;
        src162 <= 12'h39c;
        src163 <= 12'he5a;
        src164 <= 12'hd;
        src165 <= 12'h59a;
        src166 <= 12'hcbd;
        src167 <= 12'h775;
        src168 <= 12'he76;
        src169 <= 12'hbee;
        src170 <= 12'h2e;
        src171 <= 12'h920;
        src172 <= 12'hee6;
        src173 <= 12'h276;
        src174 <= 12'hb9d;
        src175 <= 12'h12c;
        src176 <= 12'h9bd;
        src177 <= 12'hc26;
        src178 <= 12'hc47;
        src179 <= 12'hc78;
        src180 <= 12'h5f7;
        src181 <= 12'h374;
        src182 <= 12'h8b0;
        src183 <= 12'h85b;
        src184 <= 12'hdaf;
        src185 <= 12'hf50;
        src186 <= 12'hca;
        src187 <= 12'h718;
        src188 <= 12'h71b;
        exp <= 20'h63348;
        #1
        src0 <= 12'hf2e;
        src1 <= 12'h4fa;
        src2 <= 12'hb96;
        src3 <= 12'hafe;
        src4 <= 12'h369;
        src5 <= 12'h593;
        src6 <= 12'h63e;
        src7 <= 12'hae5;
        src8 <= 12'ha13;
        src9 <= 12'h103;
        src10 <= 12'h274;
        src11 <= 12'h345;
        src12 <= 12'h13d;
        src13 <= 12'hd50;
        src14 <= 12'hf20;
        src15 <= 12'hd59;
        src16 <= 12'hfea;
        src17 <= 12'hb36;
        src18 <= 12'hd89;
        src19 <= 12'h1c2;
        src20 <= 12'hecb;
        src21 <= 12'he25;
        src22 <= 12'hfcc;
        src23 <= 12'h91b;
        src24 <= 12'hb24;
        src25 <= 12'h950;
        src26 <= 12'h14c;
        src27 <= 12'hd86;
        src28 <= 12'h156;
        src29 <= 12'ha19;
        src30 <= 12'hc01;
        src31 <= 12'heda;
        src32 <= 12'h7cc;
        src33 <= 12'h12c;
        src34 <= 12'ha3c;
        src35 <= 12'haa8;
        src36 <= 12'h5eb;
        src37 <= 12'h696;
        src38 <= 12'h429;
        src39 <= 12'hf3e;
        src40 <= 12'he83;
        src41 <= 12'h3b8;
        src42 <= 12'hcb3;
        src43 <= 12'h532;
        src44 <= 12'hab;
        src45 <= 12'ha6f;
        src46 <= 12'h44e;
        src47 <= 12'h60d;
        src48 <= 12'h8c5;
        src49 <= 12'h3df;
        src50 <= 12'hde6;
        src51 <= 12'h7b4;
        src52 <= 12'ha2f;
        src53 <= 12'h49c;
        src54 <= 12'h8f8;
        src55 <= 12'h52a;
        src56 <= 12'h4a8;
        src57 <= 12'h7f2;
        src58 <= 12'h2a5;
        src59 <= 12'h707;
        src60 <= 12'hb86;
        src61 <= 12'hc;
        src62 <= 12'hf4b;
        src63 <= 12'hebd;
        src64 <= 12'h418;
        src65 <= 12'h340;
        src66 <= 12'hf9e;
        src67 <= 12'hf4e;
        src68 <= 12'he6c;
        src69 <= 12'haac;
        src70 <= 12'h2c4;
        src71 <= 12'h57d;
        src72 <= 12'h462;
        src73 <= 12'h27d;
        src74 <= 12'hf42;
        src75 <= 12'h171;
        src76 <= 12'h8e2;
        src77 <= 12'h6f8;
        src78 <= 12'h76;
        src79 <= 12'hfc9;
        src80 <= 12'h5ad;
        src81 <= 12'h313;
        src82 <= 12'hc60;
        src83 <= 12'h32a;
        src84 <= 12'h489;
        src85 <= 12'h742;
        src86 <= 12'he7f;
        src87 <= 12'h967;
        src88 <= 12'hb7c;
        src89 <= 12'hdcc;
        src90 <= 12'hf3b;
        src91 <= 12'h2f4;
        src92 <= 12'h35a;
        src93 <= 12'h4d0;
        src94 <= 12'he2a;
        src95 <= 12'h34a;
        src96 <= 12'he5b;
        src97 <= 12'ha34;
        src98 <= 12'h712;
        src99 <= 12'h2fe;
        src100 <= 12'h76c;
        src101 <= 12'hd63;
        src102 <= 12'h4fe;
        src103 <= 12'h7a0;
        src104 <= 12'h403;
        src105 <= 12'h869;
        src106 <= 12'heb;
        src107 <= 12'hf36;
        src108 <= 12'hd93;
        src109 <= 12'had4;
        src110 <= 12'hb0f;
        src111 <= 12'hae8;
        src112 <= 12'hf07;
        src113 <= 12'ha59;
        src114 <= 12'h5fd;
        src115 <= 12'h790;
        src116 <= 12'he87;
        src117 <= 12'hc5a;
        src118 <= 12'hc13;
        src119 <= 12'ha86;
        src120 <= 12'h355;
        src121 <= 12'h5d4;
        src122 <= 12'h9cc;
        src123 <= 12'h860;
        src124 <= 12'h448;
        src125 <= 12'ha19;
        src126 <= 12'hac2;
        src127 <= 12'hc2f;
        src128 <= 12'h4cf;
        src129 <= 12'hef9;
        src130 <= 12'h8d5;
        src131 <= 12'hce3;
        src132 <= 12'h25d;
        src133 <= 12'hc7e;
        src134 <= 12'h8b0;
        src135 <= 12'h516;
        src136 <= 12'h641;
        src137 <= 12'ha48;
        src138 <= 12'h9cb;
        src139 <= 12'hd31;
        src140 <= 12'hda6;
        src141 <= 12'h193;
        src142 <= 12'h507;
        src143 <= 12'hb7c;
        src144 <= 12'hac2;
        src145 <= 12'h302;
        src146 <= 12'h7ca;
        src147 <= 12'hfd2;
        src148 <= 12'h470;
        src149 <= 12'hb11;
        src150 <= 12'hbcf;
        src151 <= 12'h5af;
        src152 <= 12'h27c;
        src153 <= 12'hf86;
        src154 <= 12'h716;
        src155 <= 12'hfe7;
        src156 <= 12'h55a;
        src157 <= 12'h963;
        src158 <= 12'h930;
        src159 <= 12'h66b;
        src160 <= 12'hf8d;
        src161 <= 12'h61;
        src162 <= 12'h4db;
        src163 <= 12'ha41;
        src164 <= 12'he68;
        src165 <= 12'h709;
        src166 <= 12'h47;
        src167 <= 12'hfbe;
        src168 <= 12'hdca;
        src169 <= 12'h3f2;
        src170 <= 12'h6ce;
        src171 <= 12'h357;
        src172 <= 12'h947;
        src173 <= 12'hcb9;
        src174 <= 12'h43a;
        src175 <= 12'hc7e;
        src176 <= 12'ha9c;
        src177 <= 12'hfb3;
        src178 <= 12'hd0d;
        src179 <= 12'hfec;
        src180 <= 12'h596;
        src181 <= 12'h965;
        src182 <= 12'h42c;
        src183 <= 12'hf34;
        src184 <= 12'h1a6;
        src185 <= 12'hc26;
        src186 <= 12'hafd;
        src187 <= 12'hb2f;
        src188 <= 12'h83e;
        exp <= 20'h6714d;
        #1
        src0 <= 12'h841;
        src1 <= 12'hb55;
        src2 <= 12'he3;
        src3 <= 12'h2a;
        src4 <= 12'h906;
        src5 <= 12'hbaa;
        src6 <= 12'h8c0;
        src7 <= 12'hcee;
        src8 <= 12'h532;
        src9 <= 12'hf59;
        src10 <= 12'h835;
        src11 <= 12'hdcf;
        src12 <= 12'hf12;
        src13 <= 12'h9d6;
        src14 <= 12'h5b5;
        src15 <= 12'h5f0;
        src16 <= 12'hed6;
        src17 <= 12'h88c;
        src18 <= 12'h14c;
        src19 <= 12'hd1f;
        src20 <= 12'hdb4;
        src21 <= 12'heae;
        src22 <= 12'h31f;
        src23 <= 12'hab7;
        src24 <= 12'h74f;
        src25 <= 12'h2fa;
        src26 <= 12'ha83;
        src27 <= 12'h3b4;
        src28 <= 12'h935;
        src29 <= 12'h8c0;
        src30 <= 12'h386;
        src31 <= 12'h30;
        src32 <= 12'h816;
        src33 <= 12'h953;
        src34 <= 12'ha0;
        src35 <= 12'h901;
        src36 <= 12'h2cb;
        src37 <= 12'hb46;
        src38 <= 12'hfe2;
        src39 <= 12'h51b;
        src40 <= 12'h93;
        src41 <= 12'h57b;
        src42 <= 12'he7;
        src43 <= 12'h799;
        src44 <= 12'h796;
        src45 <= 12'h23a;
        src46 <= 12'hff2;
        src47 <= 12'h708;
        src48 <= 12'h54e;
        src49 <= 12'h130;
        src50 <= 12'h965;
        src51 <= 12'hd6;
        src52 <= 12'h412;
        src53 <= 12'h567;
        src54 <= 12'hc28;
        src55 <= 12'ha80;
        src56 <= 12'h784;
        src57 <= 12'h946;
        src58 <= 12'h8f5;
        src59 <= 12'h1ee;
        src60 <= 12'hf9b;
        src61 <= 12'h5dc;
        src62 <= 12'hdb2;
        src63 <= 12'h83d;
        src64 <= 12'h886;
        src65 <= 12'hf63;
        src66 <= 12'h936;
        src67 <= 12'hc73;
        src68 <= 12'h15c;
        src69 <= 12'h31b;
        src70 <= 12'h321;
        src71 <= 12'hf30;
        src72 <= 12'h263;
        src73 <= 12'h84b;
        src74 <= 12'h108;
        src75 <= 12'hefa;
        src76 <= 12'he9a;
        src77 <= 12'hd1e;
        src78 <= 12'hcc5;
        src79 <= 12'h8be;
        src80 <= 12'h1ae;
        src81 <= 12'h5d4;
        src82 <= 12'hd23;
        src83 <= 12'h1ef;
        src84 <= 12'ha4f;
        src85 <= 12'h9a8;
        src86 <= 12'h973;
        src87 <= 12'h718;
        src88 <= 12'h150;
        src89 <= 12'h61d;
        src90 <= 12'h890;
        src91 <= 12'hb65;
        src92 <= 12'hdca;
        src93 <= 12'haaf;
        src94 <= 12'h5f3;
        src95 <= 12'h21b;
        src96 <= 12'h2b6;
        src97 <= 12'h0;
        src98 <= 12'h4bc;
        src99 <= 12'hb7c;
        src100 <= 12'h918;
        src101 <= 12'hfbd;
        src102 <= 12'hdd7;
        src103 <= 12'h319;
        src104 <= 12'h368;
        src105 <= 12'hab9;
        src106 <= 12'hced;
        src107 <= 12'h498;
        src108 <= 12'h72c;
        src109 <= 12'h94;
        src110 <= 12'hef8;
        src111 <= 12'h54c;
        src112 <= 12'h152;
        src113 <= 12'h11a;
        src114 <= 12'h597;
        src115 <= 12'hd29;
        src116 <= 12'h1e9;
        src117 <= 12'h9f4;
        src118 <= 12'h7a1;
        src119 <= 12'h11a;
        src120 <= 12'h447;
        src121 <= 12'h3dd;
        src122 <= 12'h757;
        src123 <= 12'hbe5;
        src124 <= 12'he6f;
        src125 <= 12'h914;
        src126 <= 12'hdb4;
        src127 <= 12'h326;
        src128 <= 12'h976;
        src129 <= 12'h23;
        src130 <= 12'h1b5;
        src131 <= 12'h988;
        src132 <= 12'ha4a;
        src133 <= 12'he8e;
        src134 <= 12'h4ed;
        src135 <= 12'hff4;
        src136 <= 12'hb8b;
        src137 <= 12'haea;
        src138 <= 12'h539;
        src139 <= 12'hc68;
        src140 <= 12'h229;
        src141 <= 12'h745;
        src142 <= 12'hb72;
        src143 <= 12'h20d;
        src144 <= 12'h5dc;
        src145 <= 12'hdcd;
        src146 <= 12'ha7;
        src147 <= 12'hcc4;
        src148 <= 12'ha35;
        src149 <= 12'h4c6;
        src150 <= 12'h2fa;
        src151 <= 12'he29;
        src152 <= 12'h542;
        src153 <= 12'h2ef;
        src154 <= 12'h14c;
        src155 <= 12'he46;
        src156 <= 12'hb78;
        src157 <= 12'h3bd;
        src158 <= 12'h5e0;
        src159 <= 12'hd78;
        src160 <= 12'h1f4;
        src161 <= 12'h918;
        src162 <= 12'h697;
        src163 <= 12'h488;
        src164 <= 12'h290;
        src165 <= 12'h260;
        src166 <= 12'ha81;
        src167 <= 12'hefd;
        src168 <= 12'h8fe;
        src169 <= 12'hdbe;
        src170 <= 12'h917;
        src171 <= 12'h681;
        src172 <= 12'h823;
        src173 <= 12'ha79;
        src174 <= 12'hbd7;
        src175 <= 12'h28a;
        src176 <= 12'h165;
        src177 <= 12'h8ce;
        src178 <= 12'h701;
        src179 <= 12'hfc2;
        src180 <= 12'hf;
        src181 <= 12'h510;
        src182 <= 12'hf66;
        src183 <= 12'hbcf;
        src184 <= 12'h6b8;
        src185 <= 12'h671;
        src186 <= 12'h65e;
        src187 <= 12'h6e9;
        src188 <= 12'hcf1;
        exp <= 20'h5c075;
        #1
        src0 <= 12'h507;
        src1 <= 12'hd5f;
        src2 <= 12'ha52;
        src3 <= 12'h8d4;
        src4 <= 12'h3c6;
        src5 <= 12'h392;
        src6 <= 12'ha51;
        src7 <= 12'he18;
        src8 <= 12'h44c;
        src9 <= 12'h94e;
        src10 <= 12'h3c3;
        src11 <= 12'hff6;
        src12 <= 12'h499;
        src13 <= 12'h3ce;
        src14 <= 12'h2cd;
        src15 <= 12'h3d4;
        src16 <= 12'hebf;
        src17 <= 12'h978;
        src18 <= 12'h33b;
        src19 <= 12'h3b5;
        src20 <= 12'h4d8;
        src21 <= 12'h867;
        src22 <= 12'hd82;
        src23 <= 12'h567;
        src24 <= 12'h370;
        src25 <= 12'hfcb;
        src26 <= 12'h76b;
        src27 <= 12'h509;
        src28 <= 12'h901;
        src29 <= 12'h9d4;
        src30 <= 12'hcf5;
        src31 <= 12'h1d7;
        src32 <= 12'ha36;
        src33 <= 12'hb29;
        src34 <= 12'h299;
        src35 <= 12'h477;
        src36 <= 12'hc1c;
        src37 <= 12'hd4a;
        src38 <= 12'h5b0;
        src39 <= 12'h226;
        src40 <= 12'hee9;
        src41 <= 12'hd46;
        src42 <= 12'h396;
        src43 <= 12'hc7;
        src44 <= 12'heb0;
        src45 <= 12'hdd7;
        src46 <= 12'h4c9;
        src47 <= 12'haae;
        src48 <= 12'he92;
        src49 <= 12'h3b2;
        src50 <= 12'h18e;
        src51 <= 12'h1f8;
        src52 <= 12'hdac;
        src53 <= 12'hacf;
        src54 <= 12'h630;
        src55 <= 12'hae3;
        src56 <= 12'h969;
        src57 <= 12'hb52;
        src58 <= 12'h410;
        src59 <= 12'h70e;
        src60 <= 12'h2b2;
        src61 <= 12'he37;
        src62 <= 12'hc3d;
        src63 <= 12'he73;
        src64 <= 12'h26f;
        src65 <= 12'he21;
        src66 <= 12'hc0f;
        src67 <= 12'h11c;
        src68 <= 12'h34e;
        src69 <= 12'h3b5;
        src70 <= 12'ha92;
        src71 <= 12'h157;
        src72 <= 12'hc63;
        src73 <= 12'hc42;
        src74 <= 12'h6bc;
        src75 <= 12'hb6d;
        src76 <= 12'h6dd;
        src77 <= 12'hd2e;
        src78 <= 12'h838;
        src79 <= 12'hdaf;
        src80 <= 12'hcde;
        src81 <= 12'h53;
        src82 <= 12'hd33;
        src83 <= 12'hc70;
        src84 <= 12'h223;
        src85 <= 12'h267;
        src86 <= 12'h749;
        src87 <= 12'h230;
        src88 <= 12'h546;
        src89 <= 12'hb72;
        src90 <= 12'h28c;
        src91 <= 12'hf47;
        src92 <= 12'h4ee;
        src93 <= 12'h583;
        src94 <= 12'h119;
        src95 <= 12'hbf2;
        src96 <= 12'h889;
        src97 <= 12'h4e6;
        src98 <= 12'he45;
        src99 <= 12'h39d;
        src100 <= 12'h5ca;
        src101 <= 12'hfe9;
        src102 <= 12'haed;
        src103 <= 12'hba9;
        src104 <= 12'h3ea;
        src105 <= 12'hbcf;
        src106 <= 12'he64;
        src107 <= 12'hd35;
        src108 <= 12'had9;
        src109 <= 12'h9bd;
        src110 <= 12'h3e5;
        src111 <= 12'h3b2;
        src112 <= 12'h56b;
        src113 <= 12'ha4c;
        src114 <= 12'h115;
        src115 <= 12'h34d;
        src116 <= 12'hb57;
        src117 <= 12'h4dd;
        src118 <= 12'h683;
        src119 <= 12'hd80;
        src120 <= 12'hf46;
        src121 <= 12'h446;
        src122 <= 12'h345;
        src123 <= 12'hec0;
        src124 <= 12'h273;
        src125 <= 12'h6ea;
        src126 <= 12'h19b;
        src127 <= 12'h33b;
        src128 <= 12'h49f;
        src129 <= 12'hd2c;
        src130 <= 12'h6c;
        src131 <= 12'h5c2;
        src132 <= 12'h569;
        src133 <= 12'h19c;
        src134 <= 12'hb76;
        src135 <= 12'h47a;
        src136 <= 12'h692;
        src137 <= 12'h52f;
        src138 <= 12'h346;
        src139 <= 12'h129;
        src140 <= 12'hcf5;
        src141 <= 12'h76f;
        src142 <= 12'he4a;
        src143 <= 12'heb9;
        src144 <= 12'hb84;
        src145 <= 12'hf57;
        src146 <= 12'h159;
        src147 <= 12'hb49;
        src148 <= 12'h5a3;
        src149 <= 12'haa0;
        src150 <= 12'ha9d;
        src151 <= 12'h480;
        src152 <= 12'h2ad;
        src153 <= 12'h1a3;
        src154 <= 12'h9ed;
        src155 <= 12'h3ee;
        src156 <= 12'h801;
        src157 <= 12'h78f;
        src158 <= 12'h983;
        src159 <= 12'h445;
        src160 <= 12'h256;
        src161 <= 12'h9c3;
        src162 <= 12'h7ae;
        src163 <= 12'hf3b;
        src164 <= 12'h5b6;
        src165 <= 12'h3e3;
        src166 <= 12'hb93;
        src167 <= 12'hae3;
        src168 <= 12'h19f;
        src169 <= 12'h29b;
        src170 <= 12'h206;
        src171 <= 12'he73;
        src172 <= 12'h6e0;
        src173 <= 12'heb1;
        src174 <= 12'h3ce;
        src175 <= 12'h1d;
        src176 <= 12'h7c3;
        src177 <= 12'he5b;
        src178 <= 12'hddf;
        src179 <= 12'h9a1;
        src180 <= 12'hd7;
        src181 <= 12'heb9;
        src182 <= 12'h444;
        src183 <= 12'h529;
        src184 <= 12'h8c0;
        src185 <= 12'h9d5;
        src186 <= 12'h180;
        src187 <= 12'hf8d;
        src188 <= 12'h535;
        exp <= 20'h5c64f;
        #1
        src0 <= 12'h6b0;
        src1 <= 12'h613;
        src2 <= 12'ha4c;
        src3 <= 12'hf39;
        src4 <= 12'h9b2;
        src5 <= 12'h7de;
        src6 <= 12'h162;
        src7 <= 12'h891;
        src8 <= 12'h8a3;
        src9 <= 12'h4e;
        src10 <= 12'h2fc;
        src11 <= 12'hfec;
        src12 <= 12'he54;
        src13 <= 12'h6ef;
        src14 <= 12'hc37;
        src15 <= 12'ha05;
        src16 <= 12'hfc4;
        src17 <= 12'h8ce;
        src18 <= 12'h10e;
        src19 <= 12'h312;
        src20 <= 12'hdd9;
        src21 <= 12'h23e;
        src22 <= 12'h84e;
        src23 <= 12'h411;
        src24 <= 12'h497;
        src25 <= 12'h199;
        src26 <= 12'hc7c;
        src27 <= 12'h3d2;
        src28 <= 12'h641;
        src29 <= 12'h37c;
        src30 <= 12'hc4;
        src31 <= 12'h952;
        src32 <= 12'hdd2;
        src33 <= 12'h1f8;
        src34 <= 12'h59d;
        src35 <= 12'h282;
        src36 <= 12'hc7f;
        src37 <= 12'h94c;
        src38 <= 12'hec9;
        src39 <= 12'hc93;
        src40 <= 12'h476;
        src41 <= 12'hd5a;
        src42 <= 12'hc3;
        src43 <= 12'habf;
        src44 <= 12'h355;
        src45 <= 12'hc9e;
        src46 <= 12'h6ed;
        src47 <= 12'hc15;
        src48 <= 12'h9a4;
        src49 <= 12'h71f;
        src50 <= 12'h173;
        src51 <= 12'h4f7;
        src52 <= 12'hc86;
        src53 <= 12'hae1;
        src54 <= 12'h343;
        src55 <= 12'hdcc;
        src56 <= 12'hff4;
        src57 <= 12'h1cd;
        src58 <= 12'h35d;
        src59 <= 12'h781;
        src60 <= 12'h385;
        src61 <= 12'hdda;
        src62 <= 12'h21;
        src63 <= 12'h18e;
        src64 <= 12'h76f;
        src65 <= 12'h47f;
        src66 <= 12'heb2;
        src67 <= 12'hb76;
        src68 <= 12'hc9;
        src69 <= 12'he2b;
        src70 <= 12'h70a;
        src71 <= 12'h9c9;
        src72 <= 12'h30d;
        src73 <= 12'hc7;
        src74 <= 12'h383;
        src75 <= 12'h9a5;
        src76 <= 12'heb1;
        src77 <= 12'h6eb;
        src78 <= 12'ha86;
        src79 <= 12'h482;
        src80 <= 12'h816;
        src81 <= 12'h5fd;
        src82 <= 12'h7d9;
        src83 <= 12'hb10;
        src84 <= 12'h1fc;
        src85 <= 12'h985;
        src86 <= 12'h1ce;
        src87 <= 12'hd16;
        src88 <= 12'hfd7;
        src89 <= 12'h7d;
        src90 <= 12'h45a;
        src91 <= 12'h495;
        src92 <= 12'hf42;
        src93 <= 12'h9e2;
        src94 <= 12'h4e5;
        src95 <= 12'h815;
        src96 <= 12'h1ad;
        src97 <= 12'hc83;
        src98 <= 12'h636;
        src99 <= 12'hc5e;
        src100 <= 12'h692;
        src101 <= 12'h8b5;
        src102 <= 12'h7c7;
        src103 <= 12'h218;
        src104 <= 12'h294;
        src105 <= 12'h44;
        src106 <= 12'h2bd;
        src107 <= 12'hf0a;
        src108 <= 12'hab4;
        src109 <= 12'h228;
        src110 <= 12'hdfc;
        src111 <= 12'h258;
        src112 <= 12'ha90;
        src113 <= 12'h184;
        src114 <= 12'h402;
        src115 <= 12'h274;
        src116 <= 12'h484;
        src117 <= 12'h529;
        src118 <= 12'hb54;
        src119 <= 12'hfcd;
        src120 <= 12'h257;
        src121 <= 12'hab4;
        src122 <= 12'h5c7;
        src123 <= 12'hd1;
        src124 <= 12'hc33;
        src125 <= 12'hb82;
        src126 <= 12'h91f;
        src127 <= 12'ha07;
        src128 <= 12'h46c;
        src129 <= 12'h824;
        src130 <= 12'h9f3;
        src131 <= 12'hb07;
        src132 <= 12'h6b4;
        src133 <= 12'h9f9;
        src134 <= 12'h1cc;
        src135 <= 12'hc31;
        src136 <= 12'h911;
        src137 <= 12'hf01;
        src138 <= 12'h387;
        src139 <= 12'h627;
        src140 <= 12'hdc5;
        src141 <= 12'hb8a;
        src142 <= 12'hd77;
        src143 <= 12'hd50;
        src144 <= 12'h447;
        src145 <= 12'hf72;
        src146 <= 12'h174;
        src147 <= 12'ha8e;
        src148 <= 12'h4a1;
        src149 <= 12'hf24;
        src150 <= 12'h2fa;
        src151 <= 12'h8cd;
        src152 <= 12'h5bc;
        src153 <= 12'h58a;
        src154 <= 12'h1a9;
        src155 <= 12'h2b2;
        src156 <= 12'hd94;
        src157 <= 12'h2ae;
        src158 <= 12'h1e8;
        src159 <= 12'h488;
        src160 <= 12'h930;
        src161 <= 12'h9f1;
        src162 <= 12'hd1d;
        src163 <= 12'h8ce;
        src164 <= 12'h275;
        src165 <= 12'h3c3;
        src166 <= 12'h2b3;
        src167 <= 12'hfee;
        src168 <= 12'h208;
        src169 <= 12'h98c;
        src170 <= 12'h6b6;
        src171 <= 12'h30e;
        src172 <= 12'h218;
        src173 <= 12'h7f2;
        src174 <= 12'h195;
        src175 <= 12'h5e3;
        src176 <= 12'hd81;
        src177 <= 12'h15c;
        src178 <= 12'hb61;
        src179 <= 12'hf3b;
        src180 <= 12'h966;
        src181 <= 12'hbf3;
        src182 <= 12'h507;
        src183 <= 12'h630;
        src184 <= 12'h5da;
        src185 <= 12'hbe3;
        src186 <= 12'h766;
        src187 <= 12'hf5f;
        src188 <= 12'h735;
        exp <= 20'h59b34;
        #1
        src0 <= 12'hb1d;
        src1 <= 12'hafd;
        src2 <= 12'he7c;
        src3 <= 12'h57e;
        src4 <= 12'ha3f;
        src5 <= 12'h1bf;
        src6 <= 12'h73;
        src7 <= 12'h2c5;
        src8 <= 12'h130;
        src9 <= 12'h46f;
        src10 <= 12'haeb;
        src11 <= 12'h4e9;
        src12 <= 12'he66;
        src13 <= 12'hefd;
        src14 <= 12'hb68;
        src15 <= 12'h802;
        src16 <= 12'h698;
        src17 <= 12'hc79;
        src18 <= 12'h779;
        src19 <= 12'hc72;
        src20 <= 12'h25a;
        src21 <= 12'hcde;
        src22 <= 12'h329;
        src23 <= 12'h36e;
        src24 <= 12'h6b3;
        src25 <= 12'hc45;
        src26 <= 12'h743;
        src27 <= 12'h2a4;
        src28 <= 12'hf81;
        src29 <= 12'h95;
        src30 <= 12'h27c;
        src31 <= 12'h473;
        src32 <= 12'h360;
        src33 <= 12'hb88;
        src34 <= 12'h97f;
        src35 <= 12'h5b6;
        src36 <= 12'h554;
        src37 <= 12'hd9a;
        src38 <= 12'h5b9;
        src39 <= 12'hfc;
        src40 <= 12'hcb0;
        src41 <= 12'h61b;
        src42 <= 12'ha7;
        src43 <= 12'hce7;
        src44 <= 12'he4f;
        src45 <= 12'h825;
        src46 <= 12'h1b7;
        src47 <= 12'h25a;
        src48 <= 12'h52f;
        src49 <= 12'hfb6;
        src50 <= 12'h803;
        src51 <= 12'ha2f;
        src52 <= 12'ha11;
        src53 <= 12'h2d4;
        src54 <= 12'h1f;
        src55 <= 12'hf92;
        src56 <= 12'h1f3;
        src57 <= 12'h2f0;
        src58 <= 12'h4b7;
        src59 <= 12'hef2;
        src60 <= 12'h43a;
        src61 <= 12'h240;
        src62 <= 12'haa;
        src63 <= 12'h9c5;
        src64 <= 12'h55;
        src65 <= 12'heab;
        src66 <= 12'hf92;
        src67 <= 12'hdae;
        src68 <= 12'he4b;
        src69 <= 12'h896;
        src70 <= 12'h5f6;
        src71 <= 12'hdb9;
        src72 <= 12'h4d9;
        src73 <= 12'h3d8;
        src74 <= 12'h61b;
        src75 <= 12'h98b;
        src76 <= 12'hea6;
        src77 <= 12'h953;
        src78 <= 12'h6bb;
        src79 <= 12'h8cf;
        src80 <= 12'hca9;
        src81 <= 12'heec;
        src82 <= 12'hecc;
        src83 <= 12'hb7a;
        src84 <= 12'h6f6;
        src85 <= 12'hc0;
        src86 <= 12'heda;
        src87 <= 12'h93;
        src88 <= 12'ha72;
        src89 <= 12'h5fd;
        src90 <= 12'h44e;
        src91 <= 12'ha4;
        src92 <= 12'hdd5;
        src93 <= 12'h81f;
        src94 <= 12'hb60;
        src95 <= 12'h571;
        src96 <= 12'h7;
        src97 <= 12'hfcc;
        src98 <= 12'hd3d;
        src99 <= 12'h1df;
        src100 <= 12'hcf7;
        src101 <= 12'h963;
        src102 <= 12'h319;
        src103 <= 12'h167;
        src104 <= 12'hfdb;
        src105 <= 12'h7cf;
        src106 <= 12'h250;
        src107 <= 12'hde3;
        src108 <= 12'h712;
        src109 <= 12'h26b;
        src110 <= 12'h9af;
        src111 <= 12'hb0b;
        src112 <= 12'h2fb;
        src113 <= 12'hea0;
        src114 <= 12'h5a4;
        src115 <= 12'hd84;
        src116 <= 12'h8be;
        src117 <= 12'hf8e;
        src118 <= 12'ha7a;
        src119 <= 12'hfc;
        src120 <= 12'h6c8;
        src121 <= 12'h128;
        src122 <= 12'h330;
        src123 <= 12'h682;
        src124 <= 12'hf17;
        src125 <= 12'hb61;
        src126 <= 12'h49d;
        src127 <= 12'h75a;
        src128 <= 12'hc6b;
        src129 <= 12'hf57;
        src130 <= 12'hfce;
        src131 <= 12'h685;
        src132 <= 12'hd01;
        src133 <= 12'hdab;
        src134 <= 12'ha8e;
        src135 <= 12'h25;
        src136 <= 12'h34c;
        src137 <= 12'ha78;
        src138 <= 12'h1b5;
        src139 <= 12'h181;
        src140 <= 12'h568;
        src141 <= 12'h662;
        src142 <= 12'h13a;
        src143 <= 12'h75b;
        src144 <= 12'h760;
        src145 <= 12'h73;
        src146 <= 12'hc89;
        src147 <= 12'hed4;
        src148 <= 12'h5f5;
        src149 <= 12'heef;
        src150 <= 12'h3f3;
        src151 <= 12'h2;
        src152 <= 12'hdc2;
        src153 <= 12'h6e5;
        src154 <= 12'h59e;
        src155 <= 12'he39;
        src156 <= 12'haa6;
        src157 <= 12'hfb3;
        src158 <= 12'haf4;
        src159 <= 12'h4d;
        src160 <= 12'h25b;
        src161 <= 12'h9ce;
        src162 <= 12'h98b;
        src163 <= 12'hf99;
        src164 <= 12'h493;
        src165 <= 12'ha32;
        src166 <= 12'h2b1;
        src167 <= 12'hb36;
        src168 <= 12'hcd;
        src169 <= 12'he95;
        src170 <= 12'h6dc;
        src171 <= 12'h4b;
        src172 <= 12'hc9d;
        src173 <= 12'hb7e;
        src174 <= 12'h9cd;
        src175 <= 12'hc80;
        src176 <= 12'hf6e;
        src177 <= 12'h3c9;
        src178 <= 12'h92f;
        src179 <= 12'h4df;
        src180 <= 12'hf1a;
        src181 <= 12'hfe8;
        src182 <= 12'ha6c;
        src183 <= 12'hfa3;
        src184 <= 12'h3f4;
        src185 <= 12'hfc4;
        src186 <= 12'h37f;
        src187 <= 12'h25;
        src188 <= 12'h879;
        exp <= 20'h5f83d;
        #1
        src0 <= 12'hbc6;
        src1 <= 12'h939;
        src2 <= 12'hba8;
        src3 <= 12'h9ca;
        src4 <= 12'hde4;
        src5 <= 12'h559;
        src6 <= 12'hc41;
        src7 <= 12'hb52;
        src8 <= 12'ha8e;
        src9 <= 12'h2e5;
        src10 <= 12'hd7a;
        src11 <= 12'h896;
        src12 <= 12'hedb;
        src13 <= 12'hf46;
        src14 <= 12'h8b3;
        src15 <= 12'h3da;
        src16 <= 12'hb0c;
        src17 <= 12'hd91;
        src18 <= 12'h305;
        src19 <= 12'hd65;
        src20 <= 12'hd55;
        src21 <= 12'h9ee;
        src22 <= 12'h6fe;
        src23 <= 12'h382;
        src24 <= 12'hc55;
        src25 <= 12'hcb9;
        src26 <= 12'h8a2;
        src27 <= 12'hd79;
        src28 <= 12'h35b;
        src29 <= 12'h3ad;
        src30 <= 12'h51c;
        src31 <= 12'hd10;
        src32 <= 12'h487;
        src33 <= 12'hc46;
        src34 <= 12'h42e;
        src35 <= 12'h35c;
        src36 <= 12'h8b0;
        src37 <= 12'h3f;
        src38 <= 12'h337;
        src39 <= 12'ha50;
        src40 <= 12'h74;
        src41 <= 12'hcc1;
        src42 <= 12'ha5;
        src43 <= 12'h8c6;
        src44 <= 12'h76b;
        src45 <= 12'h722;
        src46 <= 12'hb58;
        src47 <= 12'hc6e;
        src48 <= 12'he83;
        src49 <= 12'h1dc;
        src50 <= 12'h4f0;
        src51 <= 12'h529;
        src52 <= 12'he1b;
        src53 <= 12'hfd1;
        src54 <= 12'h28e;
        src55 <= 12'h892;
        src56 <= 12'h235;
        src57 <= 12'h166;
        src58 <= 12'h56e;
        src59 <= 12'hfd7;
        src60 <= 12'h5b7;
        src61 <= 12'hba5;
        src62 <= 12'hdfe;
        src63 <= 12'h334;
        src64 <= 12'h5d;
        src65 <= 12'h887;
        src66 <= 12'hbd4;
        src67 <= 12'h31c;
        src68 <= 12'h6d8;
        src69 <= 12'hae1;
        src70 <= 12'h964;
        src71 <= 12'hd1d;
        src72 <= 12'hed2;
        src73 <= 12'h631;
        src74 <= 12'hdf;
        src75 <= 12'h49c;
        src76 <= 12'hed1;
        src77 <= 12'h8fa;
        src78 <= 12'h60;
        src79 <= 12'hba2;
        src80 <= 12'hbe0;
        src81 <= 12'heb6;
        src82 <= 12'h670;
        src83 <= 12'hde9;
        src84 <= 12'h562;
        src85 <= 12'hf6b;
        src86 <= 12'h1a;
        src87 <= 12'he0d;
        src88 <= 12'h8b2;
        src89 <= 12'hfb9;
        src90 <= 12'hafd;
        src91 <= 12'h329;
        src92 <= 12'ha8a;
        src93 <= 12'hb41;
        src94 <= 12'h4cc;
        src95 <= 12'hf87;
        src96 <= 12'hf0c;
        src97 <= 12'hb76;
        src98 <= 12'h7a0;
        src99 <= 12'heba;
        src100 <= 12'h46b;
        src101 <= 12'hcba;
        src102 <= 12'h95e;
        src103 <= 12'hbdb;
        src104 <= 12'h700;
        src105 <= 12'h431;
        src106 <= 12'h66a;
        src107 <= 12'h433;
        src108 <= 12'hce2;
        src109 <= 12'h1c4;
        src110 <= 12'h488;
        src111 <= 12'h539;
        src112 <= 12'h191;
        src113 <= 12'h71d;
        src114 <= 12'h98c;
        src115 <= 12'h1d7;
        src116 <= 12'h25d;
        src117 <= 12'ha22;
        src118 <= 12'hc25;
        src119 <= 12'h5f1;
        src120 <= 12'h95e;
        src121 <= 12'h630;
        src122 <= 12'hdb3;
        src123 <= 12'hf39;
        src124 <= 12'h745;
        src125 <= 12'haf7;
        src126 <= 12'h9e7;
        src127 <= 12'hce;
        src128 <= 12'h55d;
        src129 <= 12'h2bd;
        src130 <= 12'h37;
        src131 <= 12'h9e7;
        src132 <= 12'hdf9;
        src133 <= 12'h747;
        src134 <= 12'hc52;
        src135 <= 12'h132;
        src136 <= 12'h4db;
        src137 <= 12'hbbb;
        src138 <= 12'h623;
        src139 <= 12'ha68;
        src140 <= 12'h5df;
        src141 <= 12'h3f7;
        src142 <= 12'h5d8;
        src143 <= 12'h6a8;
        src144 <= 12'h21e;
        src145 <= 12'h7d2;
        src146 <= 12'h84b;
        src147 <= 12'h3b8;
        src148 <= 12'h13a;
        src149 <= 12'h79d;
        src150 <= 12'h306;
        src151 <= 12'hb6b;
        src152 <= 12'h11c;
        src153 <= 12'hc4b;
        src154 <= 12'h78a;
        src155 <= 12'h880;
        src156 <= 12'hb87;
        src157 <= 12'hf61;
        src158 <= 12'h9d9;
        src159 <= 12'h6;
        src160 <= 12'h40;
        src161 <= 12'h483;
        src162 <= 12'h16b;
        src163 <= 12'hb26;
        src164 <= 12'h112;
        src165 <= 12'hd4b;
        src166 <= 12'hfd4;
        src167 <= 12'h9e4;
        src168 <= 12'hbc5;
        src169 <= 12'h5db;
        src170 <= 12'h27d;
        src171 <= 12'hfea;
        src172 <= 12'hb2;
        src173 <= 12'h5b;
        src174 <= 12'hce2;
        src175 <= 12'h4db;
        src176 <= 12'he44;
        src177 <= 12'h273;
        src178 <= 12'h59b;
        src179 <= 12'h81;
        src180 <= 12'h2ec;
        src181 <= 12'h184;
        src182 <= 12'h80c;
        src183 <= 12'he21;
        src184 <= 12'h2c2;
        src185 <= 12'h258;
        src186 <= 12'h16d;
        src187 <= 12'h12a;
        src188 <= 12'hbca;
        exp <= 20'h5d4c1;
        #1
        src0 <= 12'h5da;
        src1 <= 12'h9c5;
        src2 <= 12'hb8d;
        src3 <= 12'ha90;
        src4 <= 12'h60e;
        src5 <= 12'hc36;
        src6 <= 12'h450;
        src7 <= 12'hada;
        src8 <= 12'h8f8;
        src9 <= 12'h4df;
        src10 <= 12'h71d;
        src11 <= 12'h19f;
        src12 <= 12'h5d4;
        src13 <= 12'ha6b;
        src14 <= 12'hd96;
        src15 <= 12'h825;
        src16 <= 12'h8c5;
        src17 <= 12'h3ab;
        src18 <= 12'h9b1;
        src19 <= 12'h4b9;
        src20 <= 12'h5a3;
        src21 <= 12'h953;
        src22 <= 12'h5d6;
        src23 <= 12'ha20;
        src24 <= 12'h774;
        src25 <= 12'h72c;
        src26 <= 12'h6eb;
        src27 <= 12'hb86;
        src28 <= 12'hfd8;
        src29 <= 12'hd70;
        src30 <= 12'hfd0;
        src31 <= 12'h37b;
        src32 <= 12'h43f;
        src33 <= 12'h670;
        src34 <= 12'h1f5;
        src35 <= 12'h1c1;
        src36 <= 12'h319;
        src37 <= 12'he99;
        src38 <= 12'h49b;
        src39 <= 12'he76;
        src40 <= 12'hc51;
        src41 <= 12'h3e3;
        src42 <= 12'hf49;
        src43 <= 12'h218;
        src44 <= 12'h2f8;
        src45 <= 12'h95f;
        src46 <= 12'h5c4;
        src47 <= 12'h215;
        src48 <= 12'hdff;
        src49 <= 12'hc40;
        src50 <= 12'hfef;
        src51 <= 12'h238;
        src52 <= 12'h809;
        src53 <= 12'he07;
        src54 <= 12'he66;
        src55 <= 12'h24d;
        src56 <= 12'h580;
        src57 <= 12'ha2;
        src58 <= 12'h57;
        src59 <= 12'hd27;
        src60 <= 12'hc88;
        src61 <= 12'h378;
        src62 <= 12'h3b3;
        src63 <= 12'hd6b;
        src64 <= 12'he23;
        src65 <= 12'hf7e;
        src66 <= 12'h189;
        src67 <= 12'h2c3;
        src68 <= 12'h416;
        src69 <= 12'h3a8;
        src70 <= 12'hc47;
        src71 <= 12'h997;
        src72 <= 12'haa0;
        src73 <= 12'h182;
        src74 <= 12'h8ca;
        src75 <= 12'he7e;
        src76 <= 12'h2d5;
        src77 <= 12'ha08;
        src78 <= 12'h538;
        src79 <= 12'h4bc;
        src80 <= 12'h9a;
        src81 <= 12'h6e0;
        src82 <= 12'h701;
        src83 <= 12'h30f;
        src84 <= 12'he3d;
        src85 <= 12'h94;
        src86 <= 12'h8c1;
        src87 <= 12'hbf4;
        src88 <= 12'h91;
        src89 <= 12'h76c;
        src90 <= 12'h8e3;
        src91 <= 12'haa8;
        src92 <= 12'hebf;
        src93 <= 12'h2ce;
        src94 <= 12'h534;
        src95 <= 12'hd1d;
        src96 <= 12'h1f5;
        src97 <= 12'h29a;
        src98 <= 12'h33c;
        src99 <= 12'heb3;
        src100 <= 12'h4de;
        src101 <= 12'h747;
        src102 <= 12'h2d4;
        src103 <= 12'hd90;
        src104 <= 12'hfd8;
        src105 <= 12'hdf5;
        src106 <= 12'h349;
        src107 <= 12'h218;
        src108 <= 12'hf12;
        src109 <= 12'h536;
        src110 <= 12'h485;
        src111 <= 12'had0;
        src112 <= 12'h845;
        src113 <= 12'h6dc;
        src114 <= 12'h56a;
        src115 <= 12'hce9;
        src116 <= 12'h252;
        src117 <= 12'ha15;
        src118 <= 12'hdc0;
        src119 <= 12'hb16;
        src120 <= 12'hef1;
        src121 <= 12'hc8a;
        src122 <= 12'h381;
        src123 <= 12'hdfb;
        src124 <= 12'hfc0;
        src125 <= 12'hac1;
        src126 <= 12'hf6;
        src127 <= 12'hdaf;
        src128 <= 12'ha10;
        src129 <= 12'hf19;
        src130 <= 12'hed;
        src131 <= 12'h404;
        src132 <= 12'h4ab;
        src133 <= 12'he2f;
        src134 <= 12'hb8;
        src135 <= 12'ha56;
        src136 <= 12'hacf;
        src137 <= 12'h4cb;
        src138 <= 12'h319;
        src139 <= 12'h2be;
        src140 <= 12'hb04;
        src141 <= 12'h3a1;
        src142 <= 12'ha34;
        src143 <= 12'ha2a;
        src144 <= 12'h563;
        src145 <= 12'hef8;
        src146 <= 12'h29e;
        src147 <= 12'he2e;
        src148 <= 12'hd8a;
        src149 <= 12'hc03;
        src150 <= 12'h10d;
        src151 <= 12'h1cc;
        src152 <= 12'h8f3;
        src153 <= 12'h24d;
        src154 <= 12'h12;
        src155 <= 12'h6e2;
        src156 <= 12'h7fc;
        src157 <= 12'hf58;
        src158 <= 12'he95;
        src159 <= 12'h341;
        src160 <= 12'h60;
        src161 <= 12'h4f1;
        src162 <= 12'h1f;
        src163 <= 12'h4b1;
        src164 <= 12'he6b;
        src165 <= 12'hb23;
        src166 <= 12'hf8e;
        src167 <= 12'h963;
        src168 <= 12'hbe7;
        src169 <= 12'h53b;
        src170 <= 12'hff5;
        src171 <= 12'h615;
        src172 <= 12'hdca;
        src173 <= 12'h74c;
        src174 <= 12'h125;
        src175 <= 12'h3a;
        src176 <= 12'h525;
        src177 <= 12'h210;
        src178 <= 12'h54d;
        src179 <= 12'hb29;
        src180 <= 12'h626;
        src181 <= 12'hbd9;
        src182 <= 12'hef1;
        src183 <= 12'h47b;
        src184 <= 12'h398;
        src185 <= 12'hefa;
        src186 <= 12'h566;
        src187 <= 12'hc22;
        src188 <= 12'hf54;
        exp <= 20'h5e0f5;
        #1
        src0 <= 12'h34;
        src1 <= 12'hfba;
        src2 <= 12'hbfc;
        src3 <= 12'h80a;
        src4 <= 12'h52d;
        src5 <= 12'h450;
        src6 <= 12'h2ae;
        src7 <= 12'h5ef;
        src8 <= 12'h88c;
        src9 <= 12'h9ce;
        src10 <= 12'h6d;
        src11 <= 12'hd4e;
        src12 <= 12'hd65;
        src13 <= 12'h802;
        src14 <= 12'h29;
        src15 <= 12'ha07;
        src16 <= 12'h40d;
        src17 <= 12'h4c0;
        src18 <= 12'h912;
        src19 <= 12'h8c6;
        src20 <= 12'hf1c;
        src21 <= 12'h196;
        src22 <= 12'ha14;
        src23 <= 12'hddd;
        src24 <= 12'h473;
        src25 <= 12'h8b2;
        src26 <= 12'h48f;
        src27 <= 12'h8e5;
        src28 <= 12'h697;
        src29 <= 12'hc26;
        src30 <= 12'h48d;
        src31 <= 12'hbac;
        src32 <= 12'h3c4;
        src33 <= 12'h27e;
        src34 <= 12'ha62;
        src35 <= 12'hc30;
        src36 <= 12'h422;
        src37 <= 12'hdc1;
        src38 <= 12'h1c7;
        src39 <= 12'h3f7;
        src40 <= 12'h3a;
        src41 <= 12'h14b;
        src42 <= 12'heee;
        src43 <= 12'hc96;
        src44 <= 12'heae;
        src45 <= 12'h504;
        src46 <= 12'h55f;
        src47 <= 12'h1;
        src48 <= 12'hd2b;
        src49 <= 12'he02;
        src50 <= 12'hf1b;
        src51 <= 12'hdb;
        src52 <= 12'hb6a;
        src53 <= 12'h8ca;
        src54 <= 12'h6c3;
        src55 <= 12'h4c4;
        src56 <= 12'h40f;
        src57 <= 12'h8b2;
        src58 <= 12'hfda;
        src59 <= 12'h488;
        src60 <= 12'haf0;
        src61 <= 12'hbbe;
        src62 <= 12'hdb7;
        src63 <= 12'h8a;
        src64 <= 12'ha37;
        src65 <= 12'h704;
        src66 <= 12'h2f8;
        src67 <= 12'hbe2;
        src68 <= 12'h391;
        src69 <= 12'h9c5;
        src70 <= 12'hd61;
        src71 <= 12'hb15;
        src72 <= 12'hb1;
        src73 <= 12'h4bd;
        src74 <= 12'hf68;
        src75 <= 12'hae0;
        src76 <= 12'h3ac;
        src77 <= 12'hcd3;
        src78 <= 12'h5a6;
        src79 <= 12'h9bb;
        src80 <= 12'h6cd;
        src81 <= 12'h283;
        src82 <= 12'h998;
        src83 <= 12'h93f;
        src84 <= 12'h247;
        src85 <= 12'heea;
        src86 <= 12'h125;
        src87 <= 12'hda8;
        src88 <= 12'h6da;
        src89 <= 12'h9d;
        src90 <= 12'h561;
        src91 <= 12'h583;
        src92 <= 12'h4d8;
        src93 <= 12'hd70;
        src94 <= 12'hd97;
        src95 <= 12'h867;
        src96 <= 12'hf67;
        src97 <= 12'h3c2;
        src98 <= 12'h9b2;
        src99 <= 12'hda7;
        src100 <= 12'hd85;
        src101 <= 12'h970;
        src102 <= 12'hca3;
        src103 <= 12'h1f6;
        src104 <= 12'hb08;
        src105 <= 12'he7b;
        src106 <= 12'hab1;
        src107 <= 12'h353;
        src108 <= 12'h8af;
        src109 <= 12'h276;
        src110 <= 12'h457;
        src111 <= 12'h849;
        src112 <= 12'hcc8;
        src113 <= 12'h877;
        src114 <= 12'h6f7;
        src115 <= 12'hc2c;
        src116 <= 12'hd6a;
        src117 <= 12'hdf3;
        src118 <= 12'h313;
        src119 <= 12'h6ab;
        src120 <= 12'hd58;
        src121 <= 12'h724;
        src122 <= 12'hdca;
        src123 <= 12'hc05;
        src124 <= 12'h186;
        src125 <= 12'hdfd;
        src126 <= 12'h6c5;
        src127 <= 12'h72e;
        src128 <= 12'he19;
        src129 <= 12'h24e;
        src130 <= 12'hf5f;
        src131 <= 12'ha98;
        src132 <= 12'heae;
        src133 <= 12'hc84;
        src134 <= 12'h998;
        src135 <= 12'h8e0;
        src136 <= 12'hb6;
        src137 <= 12'hfe5;
        src138 <= 12'hc52;
        src139 <= 12'h904;
        src140 <= 12'h646;
        src141 <= 12'h537;
        src142 <= 12'hf09;
        src143 <= 12'h947;
        src144 <= 12'hfc6;
        src145 <= 12'h859;
        src146 <= 12'h2fa;
        src147 <= 12'h4ed;
        src148 <= 12'h377;
        src149 <= 12'h4fd;
        src150 <= 12'h15;
        src151 <= 12'hc75;
        src152 <= 12'h78c;
        src153 <= 12'ha3f;
        src154 <= 12'hbee;
        src155 <= 12'h767;
        src156 <= 12'h112;
        src157 <= 12'hef9;
        src158 <= 12'h394;
        src159 <= 12'he69;
        src160 <= 12'h1fd;
        src161 <= 12'h9b2;
        src162 <= 12'h913;
        src163 <= 12'haa7;
        src164 <= 12'h4e0;
        src165 <= 12'h4e6;
        src166 <= 12'h6e8;
        src167 <= 12'h2f9;
        src168 <= 12'hc7c;
        src169 <= 12'h17b;
        src170 <= 12'hbb;
        src171 <= 12'h2ff;
        src172 <= 12'h3c9;
        src173 <= 12'h7e4;
        src174 <= 12'he64;
        src175 <= 12'h71b;
        src176 <= 12'he74;
        src177 <= 12'h1b5;
        src178 <= 12'h53b;
        src179 <= 12'haa4;
        src180 <= 12'h205;
        src181 <= 12'ha05;
        src182 <= 12'hfe6;
        src183 <= 12'hbc9;
        src184 <= 12'haf9;
        src185 <= 12'h340;
        src186 <= 12'h8bd;
        src187 <= 12'h4ae;
        src188 <= 12'ha21;
        exp <= 20'h6084d;
        #1
        src0 <= 12'h2c3;
        src1 <= 12'h208;
        src2 <= 12'h3bd;
        src3 <= 12'hdea;
        src4 <= 12'hd73;
        src5 <= 12'h1d7;
        src6 <= 12'h299;
        src7 <= 12'hbbe;
        src8 <= 12'h627;
        src9 <= 12'h866;
        src10 <= 12'h1b1;
        src11 <= 12'h7ab;
        src12 <= 12'he95;
        src13 <= 12'hb76;
        src14 <= 12'h95c;
        src15 <= 12'h940;
        src16 <= 12'hffd;
        src17 <= 12'h866;
        src18 <= 12'h293;
        src19 <= 12'h754;
        src20 <= 12'h6cb;
        src21 <= 12'hcc6;
        src22 <= 12'h257;
        src23 <= 12'hd47;
        src24 <= 12'he63;
        src25 <= 12'hdf9;
        src26 <= 12'hf76;
        src27 <= 12'h9b6;
        src28 <= 12'hb69;
        src29 <= 12'h172;
        src30 <= 12'h2c5;
        src31 <= 12'h24d;
        src32 <= 12'hd3d;
        src33 <= 12'hc06;
        src34 <= 12'h95b;
        src35 <= 12'h70c;
        src36 <= 12'h633;
        src37 <= 12'hc92;
        src38 <= 12'h9c2;
        src39 <= 12'he73;
        src40 <= 12'he3a;
        src41 <= 12'h2b;
        src42 <= 12'h7de;
        src43 <= 12'h705;
        src44 <= 12'h5cf;
        src45 <= 12'h4e0;
        src46 <= 12'h23e;
        src47 <= 12'h8bb;
        src48 <= 12'hfa7;
        src49 <= 12'h7fc;
        src50 <= 12'hdcf;
        src51 <= 12'h49a;
        src52 <= 12'h3ff;
        src53 <= 12'h9d4;
        src54 <= 12'hc76;
        src55 <= 12'hf70;
        src56 <= 12'h337;
        src57 <= 12'hfad;
        src58 <= 12'h8bd;
        src59 <= 12'hcc8;
        src60 <= 12'h63f;
        src61 <= 12'h86f;
        src62 <= 12'hd0;
        src63 <= 12'h495;
        src64 <= 12'h2e0;
        src65 <= 12'h73d;
        src66 <= 12'haf2;
        src67 <= 12'hb33;
        src68 <= 12'h9f3;
        src69 <= 12'hf1f;
        src70 <= 12'h4e2;
        src71 <= 12'hdff;
        src72 <= 12'h32d;
        src73 <= 12'h5dd;
        src74 <= 12'h54a;
        src75 <= 12'h217;
        src76 <= 12'hb7e;
        src77 <= 12'h6f4;
        src78 <= 12'h9a3;
        src79 <= 12'h1a9;
        src80 <= 12'h394;
        src81 <= 12'ha0f;
        src82 <= 12'h3b5;
        src83 <= 12'h442;
        src84 <= 12'ha87;
        src85 <= 12'hdc5;
        src86 <= 12'h44f;
        src87 <= 12'hab0;
        src88 <= 12'h16;
        src89 <= 12'h2eb;
        src90 <= 12'he1a;
        src91 <= 12'h5cc;
        src92 <= 12'hb34;
        src93 <= 12'h5a9;
        src94 <= 12'h400;
        src95 <= 12'hf5;
        src96 <= 12'h3c6;
        src97 <= 12'ha11;
        src98 <= 12'h9cb;
        src99 <= 12'h665;
        src100 <= 12'h1f;
        src101 <= 12'h701;
        src102 <= 12'h871;
        src103 <= 12'h56;
        src104 <= 12'hf98;
        src105 <= 12'ha25;
        src106 <= 12'hf4c;
        src107 <= 12'h8eb;
        src108 <= 12'h7ca;
        src109 <= 12'h127;
        src110 <= 12'h39c;
        src111 <= 12'h46b;
        src112 <= 12'hd6c;
        src113 <= 12'heed;
        src114 <= 12'heb4;
        src115 <= 12'h3ce;
        src116 <= 12'hfb1;
        src117 <= 12'h214;
        src118 <= 12'hcc2;
        src119 <= 12'h99b;
        src120 <= 12'hed;
        src121 <= 12'h7f9;
        src122 <= 12'h368;
        src123 <= 12'hcce;
        src124 <= 12'hff0;
        src125 <= 12'h71f;
        src126 <= 12'hd77;
        src127 <= 12'h13c;
        src128 <= 12'h167;
        src129 <= 12'hd6a;
        src130 <= 12'he8e;
        src131 <= 12'h3c7;
        src132 <= 12'h65f;
        src133 <= 12'h91f;
        src134 <= 12'h841;
        src135 <= 12'hf7b;
        src136 <= 12'hf57;
        src137 <= 12'hdf8;
        src138 <= 12'h6a7;
        src139 <= 12'hff0;
        src140 <= 12'h27e;
        src141 <= 12'h863;
        src142 <= 12'h1b7;
        src143 <= 12'h194;
        src144 <= 12'h1dc;
        src145 <= 12'h8d6;
        src146 <= 12'hf03;
        src147 <= 12'h710;
        src148 <= 12'h4ac;
        src149 <= 12'h668;
        src150 <= 12'hc30;
        src151 <= 12'h25;
        src152 <= 12'h31b;
        src153 <= 12'h26;
        src154 <= 12'h618;
        src155 <= 12'h7a8;
        src156 <= 12'h4b8;
        src157 <= 12'hcb1;
        src158 <= 12'hf92;
        src159 <= 12'h768;
        src160 <= 12'h510;
        src161 <= 12'h139;
        src162 <= 12'hd2f;
        src163 <= 12'h7a7;
        src164 <= 12'hda3;
        src165 <= 12'ha9d;
        src166 <= 12'hf4;
        src167 <= 12'hb3f;
        src168 <= 12'heb3;
        src169 <= 12'h81;
        src170 <= 12'hb2c;
        src171 <= 12'hf9f;
        src172 <= 12'hb76;
        src173 <= 12'h56;
        src174 <= 12'hd89;
        src175 <= 12'h204;
        src176 <= 12'hbe2;
        src177 <= 12'h8ce;
        src178 <= 12'ha3b;
        src179 <= 12'h944;
        src180 <= 12'heeb;
        src181 <= 12'h64a;
        src182 <= 12'h944;
        src183 <= 12'ha5c;
        src184 <= 12'hb0f;
        src185 <= 12'hc64;
        src186 <= 12'h796;
        src187 <= 12'h230;
        src188 <= 12'h23;
        exp <= 20'h5fb65;
        #1
        src0 <= 12'h305;
        src1 <= 12'h7c7;
        src2 <= 12'h24a;
        src3 <= 12'h445;
        src4 <= 12'he81;
        src5 <= 12'h295;
        src6 <= 12'hcbc;
        src7 <= 12'h16a;
        src8 <= 12'h46a;
        src9 <= 12'hdd6;
        src10 <= 12'hce9;
        src11 <= 12'hf50;
        src12 <= 12'h1ae;
        src13 <= 12'hcda;
        src14 <= 12'hb77;
        src15 <= 12'h896;
        src16 <= 12'h8d9;
        src17 <= 12'hc61;
        src18 <= 12'h6c2;
        src19 <= 12'h70d;
        src20 <= 12'h187;
        src21 <= 12'h4db;
        src22 <= 12'h404;
        src23 <= 12'hde4;
        src24 <= 12'h470;
        src25 <= 12'h37c;
        src26 <= 12'h47d;
        src27 <= 12'h1e8;
        src28 <= 12'h6fb;
        src29 <= 12'h62a;
        src30 <= 12'hd25;
        src31 <= 12'h9bd;
        src32 <= 12'h243;
        src33 <= 12'h128;
        src34 <= 12'h4da;
        src35 <= 12'hca7;
        src36 <= 12'h94d;
        src37 <= 12'h5ff;
        src38 <= 12'hbf6;
        src39 <= 12'h8fe;
        src40 <= 12'hae2;
        src41 <= 12'h9e6;
        src42 <= 12'hc7;
        src43 <= 12'hab3;
        src44 <= 12'h171;
        src45 <= 12'h5a8;
        src46 <= 12'h59a;
        src47 <= 12'h95c;
        src48 <= 12'hdf7;
        src49 <= 12'h3fc;
        src50 <= 12'h826;
        src51 <= 12'h5c7;
        src52 <= 12'h945;
        src53 <= 12'h84a;
        src54 <= 12'h72;
        src55 <= 12'hb5a;
        src56 <= 12'hc57;
        src57 <= 12'hb29;
        src58 <= 12'h3c5;
        src59 <= 12'h1b2;
        src60 <= 12'h9;
        src61 <= 12'h6a6;
        src62 <= 12'h238;
        src63 <= 12'hf89;
        src64 <= 12'hfc7;
        src65 <= 12'h794;
        src66 <= 12'h229;
        src67 <= 12'h469;
        src68 <= 12'h3a1;
        src69 <= 12'hd58;
        src70 <= 12'h3c3;
        src71 <= 12'h17d;
        src72 <= 12'h6f1;
        src73 <= 12'he31;
        src74 <= 12'hf1e;
        src75 <= 12'hf08;
        src76 <= 12'ha3b;
        src77 <= 12'hdf9;
        src78 <= 12'hb69;
        src79 <= 12'h968;
        src80 <= 12'hcf3;
        src81 <= 12'h4f2;
        src82 <= 12'hfe4;
        src83 <= 12'h5b2;
        src84 <= 12'ha97;
        src85 <= 12'h2f6;
        src86 <= 12'h6b9;
        src87 <= 12'ha1;
        src88 <= 12'hfcf;
        src89 <= 12'h6fe;
        src90 <= 12'h24f;
        src91 <= 12'h673;
        src92 <= 12'h69;
        src93 <= 12'he68;
        src94 <= 12'h5da;
        src95 <= 12'h5db;
        src96 <= 12'h5fb;
        src97 <= 12'h8b7;
        src98 <= 12'hded;
        src99 <= 12'h2d7;
        src100 <= 12'h82b;
        src101 <= 12'h964;
        src102 <= 12'hfc1;
        src103 <= 12'h8b9;
        src104 <= 12'h675;
        src105 <= 12'h6f8;
        src106 <= 12'h23e;
        src107 <= 12'h40c;
        src108 <= 12'h207;
        src109 <= 12'h58b;
        src110 <= 12'h80;
        src111 <= 12'hb5a;
        src112 <= 12'h19a;
        src113 <= 12'hd0b;
        src114 <= 12'h3c6;
        src115 <= 12'h716;
        src116 <= 12'h537;
        src117 <= 12'h891;
        src118 <= 12'h81d;
        src119 <= 12'h5f5;
        src120 <= 12'habc;
        src121 <= 12'hbc2;
        src122 <= 12'hcc;
        src123 <= 12'hf25;
        src124 <= 12'hfa2;
        src125 <= 12'h2fe;
        src126 <= 12'hca9;
        src127 <= 12'h7d0;
        src128 <= 12'h5fb;
        src129 <= 12'h569;
        src130 <= 12'h71c;
        src131 <= 12'hb82;
        src132 <= 12'ha2;
        src133 <= 12'h835;
        src134 <= 12'h541;
        src135 <= 12'h2ef;
        src136 <= 12'hd14;
        src137 <= 12'hfa6;
        src138 <= 12'h4c5;
        src139 <= 12'h48;
        src140 <= 12'h5ad;
        src141 <= 12'he4e;
        src142 <= 12'hd31;
        src143 <= 12'h6ea;
        src144 <= 12'h800;
        src145 <= 12'he0c;
        src146 <= 12'he21;
        src147 <= 12'h267;
        src148 <= 12'haea;
        src149 <= 12'haf;
        src150 <= 12'ha37;
        src151 <= 12'h884;
        src152 <= 12'he19;
        src153 <= 12'h138;
        src154 <= 12'h1e0;
        src155 <= 12'h76b;
        src156 <= 12'h7f5;
        src157 <= 12'h972;
        src158 <= 12'hb3a;
        src159 <= 12'h3f1;
        src160 <= 12'hebc;
        src161 <= 12'hdb8;
        src162 <= 12'h8bb;
        src163 <= 12'h87d;
        src164 <= 12'hea8;
        src165 <= 12'h84f;
        src166 <= 12'h64b;
        src167 <= 12'h5ae;
        src168 <= 12'h1cb;
        src169 <= 12'hcbd;
        src170 <= 12'h20c;
        src171 <= 12'ha7c;
        src172 <= 12'h319;
        src173 <= 12'he3f;
        src174 <= 12'hbc4;
        src175 <= 12'had2;
        src176 <= 12'hc4f;
        src177 <= 12'hbee;
        src178 <= 12'h11f;
        src179 <= 12'h627;
        src180 <= 12'h45;
        src181 <= 12'h515;
        src182 <= 12'heef;
        src183 <= 12'hc12;
        src184 <= 12'h74d;
        src185 <= 12'h948;
        src186 <= 12'hee1;
        src187 <= 12'h47e;
        src188 <= 12'hf92;
        exp <= 20'h5cdd8;
        #1
        src0 <= 12'hd0b;
        src1 <= 12'heec;
        src2 <= 12'h965;
        src3 <= 12'h996;
        src4 <= 12'h3f0;
        src5 <= 12'h8aa;
        src6 <= 12'h5e1;
        src7 <= 12'hbbf;
        src8 <= 12'hf8b;
        src9 <= 12'h519;
        src10 <= 12'ha1;
        src11 <= 12'h3e3;
        src12 <= 12'h81c;
        src13 <= 12'h993;
        src14 <= 12'he;
        src15 <= 12'he23;
        src16 <= 12'h7fd;
        src17 <= 12'hd8a;
        src18 <= 12'h7fb;
        src19 <= 12'he9f;
        src20 <= 12'he2c;
        src21 <= 12'h26e;
        src22 <= 12'he50;
        src23 <= 12'hc2d;
        src24 <= 12'h728;
        src25 <= 12'h484;
        src26 <= 12'hbff;
        src27 <= 12'h7bb;
        src28 <= 12'h48b;
        src29 <= 12'h593;
        src30 <= 12'ha7b;
        src31 <= 12'hc9e;
        src32 <= 12'hc7e;
        src33 <= 12'hb10;
        src34 <= 12'h879;
        src35 <= 12'hef4;
        src36 <= 12'hd98;
        src37 <= 12'h501;
        src38 <= 12'hd98;
        src39 <= 12'he31;
        src40 <= 12'h527;
        src41 <= 12'h33b;
        src42 <= 12'h61f;
        src43 <= 12'h620;
        src44 <= 12'hf41;
        src45 <= 12'hbbf;
        src46 <= 12'h827;
        src47 <= 12'hef5;
        src48 <= 12'h8c;
        src49 <= 12'hb0;
        src50 <= 12'hbad;
        src51 <= 12'h378;
        src52 <= 12'h78b;
        src53 <= 12'h2db;
        src54 <= 12'h66d;
        src55 <= 12'h954;
        src56 <= 12'h637;
        src57 <= 12'h530;
        src58 <= 12'he92;
        src59 <= 12'h338;
        src60 <= 12'h5fa;
        src61 <= 12'he52;
        src62 <= 12'h1c5;
        src63 <= 12'he01;
        src64 <= 12'h790;
        src65 <= 12'hea2;
        src66 <= 12'h86d;
        src67 <= 12'h2d5;
        src68 <= 12'he7f;
        src69 <= 12'h48b;
        src70 <= 12'hdf8;
        src71 <= 12'hbd8;
        src72 <= 12'hd1a;
        src73 <= 12'h172;
        src74 <= 12'h570;
        src75 <= 12'hd96;
        src76 <= 12'h872;
        src77 <= 12'h895;
        src78 <= 12'hed1;
        src79 <= 12'h8a2;
        src80 <= 12'hf22;
        src81 <= 12'ha93;
        src82 <= 12'h27c;
        src83 <= 12'h5cc;
        src84 <= 12'hcd;
        src85 <= 12'h8a8;
        src86 <= 12'hb1f;
        src87 <= 12'ha31;
        src88 <= 12'h2bc;
        src89 <= 12'hfe;
        src90 <= 12'hfe2;
        src91 <= 12'hd6b;
        src92 <= 12'hef;
        src93 <= 12'hcc5;
        src94 <= 12'h61d;
        src95 <= 12'h5bb;
        src96 <= 12'hfc4;
        src97 <= 12'h929;
        src98 <= 12'h510;
        src99 <= 12'h832;
        src100 <= 12'h303;
        src101 <= 12'h7dd;
        src102 <= 12'hab6;
        src103 <= 12'h57e;
        src104 <= 12'h1de;
        src105 <= 12'h37a;
        src106 <= 12'ha60;
        src107 <= 12'ha26;
        src108 <= 12'h51c;
        src109 <= 12'h215;
        src110 <= 12'h6ba;
        src111 <= 12'h10b;
        src112 <= 12'h5a2;
        src113 <= 12'h449;
        src114 <= 12'h5f8;
        src115 <= 12'h7f2;
        src116 <= 12'h33d;
        src117 <= 12'hc40;
        src118 <= 12'h7e4;
        src119 <= 12'h265;
        src120 <= 12'h2ff;
        src121 <= 12'hce;
        src122 <= 12'hd0;
        src123 <= 12'h581;
        src124 <= 12'h663;
        src125 <= 12'hddc;
        src126 <= 12'ha82;
        src127 <= 12'h90c;
        src128 <= 12'h5f5;
        src129 <= 12'ha38;
        src130 <= 12'h56f;
        src131 <= 12'h156;
        src132 <= 12'hc6b;
        src133 <= 12'h794;
        src134 <= 12'hc2c;
        src135 <= 12'h6b0;
        src136 <= 12'h3c7;
        src137 <= 12'hd71;
        src138 <= 12'hf33;
        src139 <= 12'h92a;
        src140 <= 12'h5f1;
        src141 <= 12'hd6c;
        src142 <= 12'hb09;
        src143 <= 12'h932;
        src144 <= 12'h6d8;
        src145 <= 12'h1dd;
        src146 <= 12'h7bc;
        src147 <= 12'hc9c;
        src148 <= 12'h5f3;
        src149 <= 12'h665;
        src150 <= 12'h910;
        src151 <= 12'he24;
        src152 <= 12'he99;
        src153 <= 12'h96b;
        src154 <= 12'h41e;
        src155 <= 12'h791;
        src156 <= 12'h76c;
        src157 <= 12'h91f;
        src158 <= 12'h5d7;
        src159 <= 12'h291;
        src160 <= 12'hd31;
        src161 <= 12'h870;
        src162 <= 12'hbac;
        src163 <= 12'hea2;
        src164 <= 12'h4d4;
        src165 <= 12'hf8;
        src166 <= 12'hcba;
        src167 <= 12'h275;
        src168 <= 12'h6d0;
        src169 <= 12'hb5;
        src170 <= 12'h742;
        src171 <= 12'hf46;
        src172 <= 12'h8e;
        src173 <= 12'he7c;
        src174 <= 12'hd94;
        src175 <= 12'hfac;
        src176 <= 12'h644;
        src177 <= 12'ha44;
        src178 <= 12'haee;
        src179 <= 12'h70b;
        src180 <= 12'h2ef;
        src181 <= 12'hdc7;
        src182 <= 12'hfcc;
        src183 <= 12'h32d;
        src184 <= 12'h2cc;
        src185 <= 12'h6ba;
        src186 <= 12'hea8;
        src187 <= 12'hd65;
        src188 <= 12'hc49;
        exp <= 20'h622c0;
        #1
        src0 <= 12'h597;
        src1 <= 12'h7b1;
        src2 <= 12'ha04;
        src3 <= 12'h3c0;
        src4 <= 12'h34e;
        src5 <= 12'h59f;
        src6 <= 12'h18a;
        src7 <= 12'h5d2;
        src8 <= 12'h378;
        src9 <= 12'hfbc;
        src10 <= 12'h860;
        src11 <= 12'h872;
        src12 <= 12'h58f;
        src13 <= 12'h9dc;
        src14 <= 12'h4bf;
        src15 <= 12'h92f;
        src16 <= 12'h867;
        src17 <= 12'hff4;
        src18 <= 12'ha51;
        src19 <= 12'hce;
        src20 <= 12'h892;
        src21 <= 12'ha82;
        src22 <= 12'hc38;
        src23 <= 12'h27c;
        src24 <= 12'h8da;
        src25 <= 12'he1e;
        src26 <= 12'hb56;
        src27 <= 12'h605;
        src28 <= 12'h3b1;
        src29 <= 12'hce7;
        src30 <= 12'hdca;
        src31 <= 12'h9a9;
        src32 <= 12'hae5;
        src33 <= 12'h334;
        src34 <= 12'h851;
        src35 <= 12'h4cf;
        src36 <= 12'hc68;
        src37 <= 12'h92b;
        src38 <= 12'h637;
        src39 <= 12'hef4;
        src40 <= 12'h974;
        src41 <= 12'ha72;
        src42 <= 12'h288;
        src43 <= 12'hc5f;
        src44 <= 12'h691;
        src45 <= 12'ha46;
        src46 <= 12'h87f;
        src47 <= 12'he8;
        src48 <= 12'hf79;
        src49 <= 12'h4d7;
        src50 <= 12'ha7b;
        src51 <= 12'h941;
        src52 <= 12'h147;
        src53 <= 12'hcdb;
        src54 <= 12'hb31;
        src55 <= 12'h62c;
        src56 <= 12'h447;
        src57 <= 12'hb3c;
        src58 <= 12'ha63;
        src59 <= 12'h985;
        src60 <= 12'h625;
        src61 <= 12'hb35;
        src62 <= 12'ha12;
        src63 <= 12'h340;
        src64 <= 12'hf3;
        src65 <= 12'hac4;
        src66 <= 12'hbae;
        src67 <= 12'h553;
        src68 <= 12'hf4;
        src69 <= 12'ha62;
        src70 <= 12'h57d;
        src71 <= 12'hd00;
        src72 <= 12'hb59;
        src73 <= 12'hcfe;
        src74 <= 12'hab1;
        src75 <= 12'h7c6;
        src76 <= 12'hf41;
        src77 <= 12'he06;
        src78 <= 12'h9aa;
        src79 <= 12'h7e4;
        src80 <= 12'hfff;
        src81 <= 12'h32f;
        src82 <= 12'h6a4;
        src83 <= 12'hc28;
        src84 <= 12'hd81;
        src85 <= 12'hd0;
        src86 <= 12'h2dc;
        src87 <= 12'h72b;
        src88 <= 12'h74e;
        src89 <= 12'h3a;
        src90 <= 12'hbc8;
        src91 <= 12'h61c;
        src92 <= 12'h8ce;
        src93 <= 12'h7a8;
        src94 <= 12'hd48;
        src95 <= 12'h711;
        src96 <= 12'he64;
        src97 <= 12'h1b6;
        src98 <= 12'h92a;
        src99 <= 12'h4a6;
        src100 <= 12'h52b;
        src101 <= 12'h285;
        src102 <= 12'he98;
        src103 <= 12'h5fa;
        src104 <= 12'h6b2;
        src105 <= 12'h9ea;
        src106 <= 12'haf0;
        src107 <= 12'hcf;
        src108 <= 12'hb8f;
        src109 <= 12'h481;
        src110 <= 12'h72a;
        src111 <= 12'hb98;
        src112 <= 12'h3be;
        src113 <= 12'h6f4;
        src114 <= 12'h390;
        src115 <= 12'h589;
        src116 <= 12'hc6f;
        src117 <= 12'h74a;
        src118 <= 12'hcb0;
        src119 <= 12'h6f0;
        src120 <= 12'h721;
        src121 <= 12'h18c;
        src122 <= 12'hc88;
        src123 <= 12'h454;
        src124 <= 12'h7cd;
        src125 <= 12'hac3;
        src126 <= 12'h20d;
        src127 <= 12'h87f;
        src128 <= 12'h33e;
        src129 <= 12'h449;
        src130 <= 12'h72c;
        src131 <= 12'h770;
        src132 <= 12'h1a7;
        src133 <= 12'hee;
        src134 <= 12'h73;
        src135 <= 12'h534;
        src136 <= 12'h53f;
        src137 <= 12'h7a3;
        src138 <= 12'h444;
        src139 <= 12'hb22;
        src140 <= 12'hbda;
        src141 <= 12'h121;
        src142 <= 12'hb73;
        src143 <= 12'h14b;
        src144 <= 12'hcaf;
        src145 <= 12'h89b;
        src146 <= 12'h59f;
        src147 <= 12'h9ec;
        src148 <= 12'h92d;
        src149 <= 12'h41e;
        src150 <= 12'h45e;
        src151 <= 12'h952;
        src152 <= 12'h44f;
        src153 <= 12'h593;
        src154 <= 12'h600;
        src155 <= 12'h665;
        src156 <= 12'h969;
        src157 <= 12'h5cd;
        src158 <= 12'h5b6;
        src159 <= 12'hc5b;
        src160 <= 12'h596;
        src161 <= 12'h160;
        src162 <= 12'h163;
        src163 <= 12'h74f;
        src164 <= 12'hd90;
        src165 <= 12'h993;
        src166 <= 12'haeb;
        src167 <= 12'h535;
        src168 <= 12'h627;
        src169 <= 12'h5a9;
        src170 <= 12'h6a6;
        src171 <= 12'hda5;
        src172 <= 12'hdca;
        src173 <= 12'haae;
        src174 <= 12'hd03;
        src175 <= 12'h420;
        src176 <= 12'h62f;
        src177 <= 12'h43b;
        src178 <= 12'hd41;
        src179 <= 12'h22a;
        src180 <= 12'h3cd;
        src181 <= 12'h3f9;
        src182 <= 12'h12f;
        src183 <= 12'h69a;
        src184 <= 12'h282;
        src185 <= 12'ha7;
        src186 <= 12'hf6a;
        src187 <= 12'h815;
        src188 <= 12'ha1;
        exp <= 20'h59be1;
        #1
        src0 <= 12'hbce;
        src1 <= 12'hf90;
        src2 <= 12'h2a5;
        src3 <= 12'hcc4;
        src4 <= 12'hdef;
        src5 <= 12'h8f6;
        src6 <= 12'h11;
        src7 <= 12'h2c9;
        src8 <= 12'h841;
        src9 <= 12'h414;
        src10 <= 12'hd21;
        src11 <= 12'h49a;
        src12 <= 12'hb9a;
        src13 <= 12'hd93;
        src14 <= 12'he8a;
        src15 <= 12'hda0;
        src16 <= 12'h3c4;
        src17 <= 12'h358;
        src18 <= 12'ha4d;
        src19 <= 12'ha7a;
        src20 <= 12'hd2e;
        src21 <= 12'h8c9;
        src22 <= 12'h5a5;
        src23 <= 12'h89;
        src24 <= 12'h90f;
        src25 <= 12'hed4;
        src26 <= 12'h3c1;
        src27 <= 12'hc11;
        src28 <= 12'h402;
        src29 <= 12'h6d4;
        src30 <= 12'hee6;
        src31 <= 12'h8ae;
        src32 <= 12'h85c;
        src33 <= 12'h480;
        src34 <= 12'hb60;
        src35 <= 12'h5bc;
        src36 <= 12'he83;
        src37 <= 12'haca;
        src38 <= 12'ha33;
        src39 <= 12'h8ab;
        src40 <= 12'h5a1;
        src41 <= 12'ha3c;
        src42 <= 12'h1e9;
        src43 <= 12'h51f;
        src44 <= 12'hf92;
        src45 <= 12'h74f;
        src46 <= 12'h4e0;
        src47 <= 12'h975;
        src48 <= 12'he32;
        src49 <= 12'h29c;
        src50 <= 12'h48;
        src51 <= 12'hb88;
        src52 <= 12'hf77;
        src53 <= 12'hd9f;
        src54 <= 12'hea7;
        src55 <= 12'h685;
        src56 <= 12'h26b;
        src57 <= 12'hf62;
        src58 <= 12'hceb;
        src59 <= 12'h514;
        src60 <= 12'h598;
        src61 <= 12'h65e;
        src62 <= 12'h77e;
        src63 <= 12'h8e1;
        src64 <= 12'hd8f;
        src65 <= 12'h36a;
        src66 <= 12'h397;
        src67 <= 12'h296;
        src68 <= 12'hd7a;
        src69 <= 12'hc75;
        src70 <= 12'h499;
        src71 <= 12'hd86;
        src72 <= 12'h3cf;
        src73 <= 12'he5e;
        src74 <= 12'hf61;
        src75 <= 12'h903;
        src76 <= 12'h6f4;
        src77 <= 12'h45;
        src78 <= 12'h36b;
        src79 <= 12'h971;
        src80 <= 12'he18;
        src81 <= 12'h2e6;
        src82 <= 12'hde;
        src83 <= 12'h5e9;
        src84 <= 12'h34c;
        src85 <= 12'h536;
        src86 <= 12'h31;
        src87 <= 12'hdd8;
        src88 <= 12'h865;
        src89 <= 12'h5e1;
        src90 <= 12'he86;
        src91 <= 12'ha54;
        src92 <= 12'h81c;
        src93 <= 12'h31c;
        src94 <= 12'he0d;
        src95 <= 12'h42e;
        src96 <= 12'h2;
        src97 <= 12'h6a5;
        src98 <= 12'h14f;
        src99 <= 12'h2b8;
        src100 <= 12'h11f;
        src101 <= 12'h8bd;
        src102 <= 12'h661;
        src103 <= 12'h219;
        src104 <= 12'hbe0;
        src105 <= 12'h3e7;
        src106 <= 12'hffb;
        src107 <= 12'h667;
        src108 <= 12'h369;
        src109 <= 12'hd7c;
        src110 <= 12'hc75;
        src111 <= 12'hed2;
        src112 <= 12'hb2f;
        src113 <= 12'hc15;
        src114 <= 12'h7fc;
        src115 <= 12'h6d0;
        src116 <= 12'hbfa;
        src117 <= 12'h36c;
        src118 <= 12'haf6;
        src119 <= 12'h7bf;
        src120 <= 12'hb0c;
        src121 <= 12'h443;
        src122 <= 12'h7b3;
        src123 <= 12'h7a8;
        src124 <= 12'h156;
        src125 <= 12'h2b0;
        src126 <= 12'h939;
        src127 <= 12'ha4a;
        src128 <= 12'hbd1;
        src129 <= 12'h1fd;
        src130 <= 12'h4ce;
        src131 <= 12'h130;
        src132 <= 12'h916;
        src133 <= 12'he6d;
        src134 <= 12'h2a1;
        src135 <= 12'h5ef;
        src136 <= 12'h828;
        src137 <= 12'h7aa;
        src138 <= 12'heba;
        src139 <= 12'h203;
        src140 <= 12'h981;
        src141 <= 12'he15;
        src142 <= 12'hc8d;
        src143 <= 12'h41d;
        src144 <= 12'h78a;
        src145 <= 12'h1f6;
        src146 <= 12'h6de;
        src147 <= 12'hf47;
        src148 <= 12'hfd4;
        src149 <= 12'h5b7;
        src150 <= 12'ha40;
        src151 <= 12'h9cb;
        src152 <= 12'h8bd;
        src153 <= 12'ha5a;
        src154 <= 12'h505;
        src155 <= 12'hec2;
        src156 <= 12'hc3d;
        src157 <= 12'ha68;
        src158 <= 12'h8a5;
        src159 <= 12'hbc6;
        src160 <= 12'h8ec;
        src161 <= 12'hf70;
        src162 <= 12'h9dc;
        src163 <= 12'hcf8;
        src164 <= 12'h79f;
        src165 <= 12'hecb;
        src166 <= 12'h96a;
        src167 <= 12'h7a7;
        src168 <= 12'hab9;
        src169 <= 12'h91f;
        src170 <= 12'h30e;
        src171 <= 12'h5d5;
        src172 <= 12'ha2a;
        src173 <= 12'h3a4;
        src174 <= 12'h30;
        src175 <= 12'h6bb;
        src176 <= 12'h2d8;
        src177 <= 12'h5a4;
        src178 <= 12'hcba;
        src179 <= 12'h475;
        src180 <= 12'h9bc;
        src181 <= 12'ha03;
        src182 <= 12'h68;
        src183 <= 12'heb;
        src184 <= 12'hde0;
        src185 <= 12'h9b6;
        src186 <= 12'hc84;
        src187 <= 12'h7a3;
        src188 <= 12'h38c;
        exp <= 20'h60fc3;
        #1
        src0 <= 12'hca9;
        src1 <= 12'h4e8;
        src2 <= 12'hd1c;
        src3 <= 12'h8ba;
        src4 <= 12'h1ec;
        src5 <= 12'h98e;
        src6 <= 12'hf63;
        src7 <= 12'h41b;
        src8 <= 12'h2e7;
        src9 <= 12'he8a;
        src10 <= 12'hb3f;
        src11 <= 12'he7c;
        src12 <= 12'h627;
        src13 <= 12'h8f;
        src14 <= 12'heb8;
        src15 <= 12'hae2;
        src16 <= 12'h8ae;
        src17 <= 12'h91a;
        src18 <= 12'h91f;
        src19 <= 12'hf1;
        src20 <= 12'h58;
        src21 <= 12'hf9d;
        src22 <= 12'h87a;
        src23 <= 12'he32;
        src24 <= 12'h4e1;
        src25 <= 12'h7f4;
        src26 <= 12'h45f;
        src27 <= 12'hf22;
        src28 <= 12'h54a;
        src29 <= 12'h3ad;
        src30 <= 12'he20;
        src31 <= 12'he38;
        src32 <= 12'h3fc;
        src33 <= 12'hced;
        src34 <= 12'h2c0;
        src35 <= 12'h838;
        src36 <= 12'h14a;
        src37 <= 12'hfd7;
        src38 <= 12'h94d;
        src39 <= 12'h601;
        src40 <= 12'h3c7;
        src41 <= 12'had5;
        src42 <= 12'h43d;
        src43 <= 12'ha5b;
        src44 <= 12'h5f8;
        src45 <= 12'h6c6;
        src46 <= 12'ha58;
        src47 <= 12'h715;
        src48 <= 12'h48d;
        src49 <= 12'h55;
        src50 <= 12'h26e;
        src51 <= 12'h4a8;
        src52 <= 12'h79b;
        src53 <= 12'h518;
        src54 <= 12'h7a6;
        src55 <= 12'h5cd;
        src56 <= 12'h3ff;
        src57 <= 12'hedb;
        src58 <= 12'h965;
        src59 <= 12'h337;
        src60 <= 12'hc55;
        src61 <= 12'h550;
        src62 <= 12'hdba;
        src63 <= 12'h489;
        src64 <= 12'h346;
        src65 <= 12'hdc9;
        src66 <= 12'h5f3;
        src67 <= 12'hc23;
        src68 <= 12'h646;
        src69 <= 12'he9d;
        src70 <= 12'h603;
        src71 <= 12'hfbd;
        src72 <= 12'he94;
        src73 <= 12'h5c7;
        src74 <= 12'h535;
        src75 <= 12'h777;
        src76 <= 12'hbf7;
        src77 <= 12'hd47;
        src78 <= 12'h78d;
        src79 <= 12'h1fb;
        src80 <= 12'hf5;
        src81 <= 12'hbdd;
        src82 <= 12'h3f8;
        src83 <= 12'hbdb;
        src84 <= 12'h7e0;
        src85 <= 12'hc9f;
        src86 <= 12'h1e0;
        src87 <= 12'h882;
        src88 <= 12'had5;
        src89 <= 12'hff3;
        src90 <= 12'hc21;
        src91 <= 12'hf17;
        src92 <= 12'h10e;
        src93 <= 12'h1e3;
        src94 <= 12'h90a;
        src95 <= 12'hc68;
        src96 <= 12'h79f;
        src97 <= 12'he3d;
        src98 <= 12'ha7c;
        src99 <= 12'he22;
        src100 <= 12'ha6f;
        src101 <= 12'hca0;
        src102 <= 12'h520;
        src103 <= 12'h10d;
        src104 <= 12'h23b;
        src105 <= 12'h86d;
        src106 <= 12'h285;
        src107 <= 12'haaa;
        src108 <= 12'h588;
        src109 <= 12'hd97;
        src110 <= 12'h69f;
        src111 <= 12'h777;
        src112 <= 12'hb72;
        src113 <= 12'h887;
        src114 <= 12'hf4b;
        src115 <= 12'h768;
        src116 <= 12'hef3;
        src117 <= 12'hd16;
        src118 <= 12'h20c;
        src119 <= 12'h5b1;
        src120 <= 12'hd25;
        src121 <= 12'hb88;
        src122 <= 12'h3ba;
        src123 <= 12'h9b8;
        src124 <= 12'h50;
        src125 <= 12'h92;
        src126 <= 12'h33d;
        src127 <= 12'h66c;
        src128 <= 12'hf2b;
        src129 <= 12'h925;
        src130 <= 12'h614;
        src131 <= 12'h1b7;
        src132 <= 12'hf45;
        src133 <= 12'h93c;
        src134 <= 12'h13f;
        src135 <= 12'hf1;
        src136 <= 12'h538;
        src137 <= 12'h80e;
        src138 <= 12'h252;
        src139 <= 12'hdd;
        src140 <= 12'h373;
        src141 <= 12'h121;
        src142 <= 12'h329;
        src143 <= 12'h3a4;
        src144 <= 12'h96c;
        src145 <= 12'h540;
        src146 <= 12'h4cc;
        src147 <= 12'ha6;
        src148 <= 12'ha49;
        src149 <= 12'h65e;
        src150 <= 12'h319;
        src151 <= 12'h1da;
        src152 <= 12'hf68;
        src153 <= 12'ha74;
        src154 <= 12'hf0c;
        src155 <= 12'h684;
        src156 <= 12'hfd;
        src157 <= 12'hdc4;
        src158 <= 12'h222;
        src159 <= 12'h2b3;
        src160 <= 12'h99a;
        src161 <= 12'hf2;
        src162 <= 12'hbb5;
        src163 <= 12'hc46;
        src164 <= 12'h4a8;
        src165 <= 12'h7ac;
        src166 <= 12'h622;
        src167 <= 12'h57a;
        src168 <= 12'hc7c;
        src169 <= 12'heee;
        src170 <= 12'h282;
        src171 <= 12'h383;
        src172 <= 12'h604;
        src173 <= 12'h855;
        src174 <= 12'h4d2;
        src175 <= 12'h4f;
        src176 <= 12'h79e;
        src177 <= 12'hc84;
        src178 <= 12'ha10;
        src179 <= 12'hf03;
        src180 <= 12'hdd0;
        src181 <= 12'he04;
        src182 <= 12'ha73;
        src183 <= 12'hdbc;
        src184 <= 12'h815;
        src185 <= 12'h727;
        src186 <= 12'h7ce;
        src187 <= 12'h83f;
        src188 <= 12'h169;
        exp <= 20'h5cf26;
        #1
        src0 <= 12'h21e;
        src1 <= 12'hf96;
        src2 <= 12'h39d;
        src3 <= 12'h36c;
        src4 <= 12'hcca;
        src5 <= 12'hc33;
        src6 <= 12'h30b;
        src7 <= 12'h5b3;
        src8 <= 12'h16a;
        src9 <= 12'h4d5;
        src10 <= 12'h4ca;
        src11 <= 12'h72e;
        src12 <= 12'h30d;
        src13 <= 12'hc3d;
        src14 <= 12'hca6;
        src15 <= 12'h3fb;
        src16 <= 12'h161;
        src17 <= 12'hc01;
        src18 <= 12'h1ea;
        src19 <= 12'hb18;
        src20 <= 12'h6c3;
        src21 <= 12'h81d;
        src22 <= 12'hc3f;
        src23 <= 12'he9a;
        src24 <= 12'h661;
        src25 <= 12'hb90;
        src26 <= 12'hc40;
        src27 <= 12'ha6d;
        src28 <= 12'hde7;
        src29 <= 12'h560;
        src30 <= 12'h7b2;
        src31 <= 12'h4c2;
        src32 <= 12'heae;
        src33 <= 12'h567;
        src34 <= 12'h84b;
        src35 <= 12'he55;
        src36 <= 12'h1fb;
        src37 <= 12'hf10;
        src38 <= 12'he8;
        src39 <= 12'h742;
        src40 <= 12'h1b9;
        src41 <= 12'hfde;
        src42 <= 12'hff3;
        src43 <= 12'hcbb;
        src44 <= 12'h923;
        src45 <= 12'hb98;
        src46 <= 12'hf7f;
        src47 <= 12'h5d3;
        src48 <= 12'h910;
        src49 <= 12'h406;
        src50 <= 12'hea9;
        src51 <= 12'h144;
        src52 <= 12'h416;
        src53 <= 12'haa4;
        src54 <= 12'hc55;
        src55 <= 12'h747;
        src56 <= 12'h529;
        src57 <= 12'hfab;
        src58 <= 12'h766;
        src59 <= 12'h646;
        src60 <= 12'hc95;
        src61 <= 12'he37;
        src62 <= 12'hb95;
        src63 <= 12'h245;
        src64 <= 12'h946;
        src65 <= 12'h626;
        src66 <= 12'h207;
        src67 <= 12'h90;
        src68 <= 12'hf11;
        src69 <= 12'h40d;
        src70 <= 12'hdb1;
        src71 <= 12'hd72;
        src72 <= 12'h37;
        src73 <= 12'hfe0;
        src74 <= 12'hfa3;
        src75 <= 12'h9f0;
        src76 <= 12'h64a;
        src77 <= 12'hecf;
        src78 <= 12'hd9c;
        src79 <= 12'ha44;
        src80 <= 12'h83f;
        src81 <= 12'h820;
        src82 <= 12'h6c1;
        src83 <= 12'h76a;
        src84 <= 12'ha38;
        src85 <= 12'h2d6;
        src86 <= 12'h243;
        src87 <= 12'h523;
        src88 <= 12'hb02;
        src89 <= 12'h8c4;
        src90 <= 12'h911;
        src91 <= 12'hf5a;
        src92 <= 12'h84;
        src93 <= 12'h9ab;
        src94 <= 12'ha7b;
        src95 <= 12'hcf4;
        src96 <= 12'h86d;
        src97 <= 12'h797;
        src98 <= 12'hc0b;
        src99 <= 12'h2af;
        src100 <= 12'h8a;
        src101 <= 12'hb29;
        src102 <= 12'hd25;
        src103 <= 12'h9bf;
        src104 <= 12'hb8b;
        src105 <= 12'h8ad;
        src106 <= 12'h4e8;
        src107 <= 12'hdc2;
        src108 <= 12'h57c;
        src109 <= 12'h7ad;
        src110 <= 12'hf13;
        src111 <= 12'hf57;
        src112 <= 12'ha3c;
        src113 <= 12'h21e;
        src114 <= 12'he01;
        src115 <= 12'h390;
        src116 <= 12'h393;
        src117 <= 12'hc60;
        src118 <= 12'hec;
        src119 <= 12'h946;
        src120 <= 12'h42d;
        src121 <= 12'hbf0;
        src122 <= 12'h21b;
        src123 <= 12'h2cc;
        src124 <= 12'h29b;
        src125 <= 12'h29f;
        src126 <= 12'hbd7;
        src127 <= 12'hf83;
        src128 <= 12'hfae;
        src129 <= 12'h1fc;
        src130 <= 12'hbbf;
        src131 <= 12'h5e8;
        src132 <= 12'hcc7;
        src133 <= 12'heb9;
        src134 <= 12'h8f5;
        src135 <= 12'h597;
        src136 <= 12'h86;
        src137 <= 12'h80;
        src138 <= 12'h619;
        src139 <= 12'hf42;
        src140 <= 12'h520;
        src141 <= 12'h33b;
        src142 <= 12'he3e;
        src143 <= 12'h8c5;
        src144 <= 12'haf9;
        src145 <= 12'heca;
        src146 <= 12'h995;
        src147 <= 12'h935;
        src148 <= 12'h32a;
        src149 <= 12'hd82;
        src150 <= 12'h261;
        src151 <= 12'h113;
        src152 <= 12'h848;
        src153 <= 12'h19b;
        src154 <= 12'h259;
        src155 <= 12'h45a;
        src156 <= 12'hd11;
        src157 <= 12'h28b;
        src158 <= 12'hd0d;
        src159 <= 12'h61f;
        src160 <= 12'h4a6;
        src161 <= 12'h788;
        src162 <= 12'ha40;
        src163 <= 12'hcdf;
        src164 <= 12'hed7;
        src165 <= 12'hf2;
        src166 <= 12'hc54;
        src167 <= 12'h654;
        src168 <= 12'hfbc;
        src169 <= 12'h2d;
        src170 <= 12'hb0f;
        src171 <= 12'h60a;
        src172 <= 12'h9fc;
        src173 <= 12'h4b5;
        src174 <= 12'h70;
        src175 <= 12'h138;
        src176 <= 12'h684;
        src177 <= 12'h167;
        src178 <= 12'h1cd;
        src179 <= 12'h234;
        src180 <= 12'hfec;
        src181 <= 12'he17;
        src182 <= 12'hae4;
        src183 <= 12'h5f2;
        src184 <= 12'h711;
        src185 <= 12'hc07;
        src186 <= 12'ha4a;
        src187 <= 12'h4af;
        src188 <= 12'h9b6;
        exp <= 20'h60dbd;
        #1
        src0 <= 12'hfc6;
        src1 <= 12'h139;
        src2 <= 12'h4a8;
        src3 <= 12'h91a;
        src4 <= 12'h49b;
        src5 <= 12'h1e4;
        src6 <= 12'hd6c;
        src7 <= 12'h974;
        src8 <= 12'hc32;
        src9 <= 12'h511;
        src10 <= 12'h61e;
        src11 <= 12'h3c6;
        src12 <= 12'hd6;
        src13 <= 12'h9e7;
        src14 <= 12'h24c;
        src15 <= 12'hf5b;
        src16 <= 12'ha53;
        src17 <= 12'h70c;
        src18 <= 12'h9b4;
        src19 <= 12'h664;
        src20 <= 12'h1de;
        src21 <= 12'h79e;
        src22 <= 12'h36f;
        src23 <= 12'h4f;
        src24 <= 12'hff2;
        src25 <= 12'h70;
        src26 <= 12'h277;
        src27 <= 12'h35c;
        src28 <= 12'hef5;
        src29 <= 12'hc71;
        src30 <= 12'hef9;
        src31 <= 12'h2b2;
        src32 <= 12'h9d6;
        src33 <= 12'h4b1;
        src34 <= 12'h5ea;
        src35 <= 12'hce8;
        src36 <= 12'h62f;
        src37 <= 12'h5d0;
        src38 <= 12'h8f3;
        src39 <= 12'h23b;
        src40 <= 12'h795;
        src41 <= 12'hce1;
        src42 <= 12'h59a;
        src43 <= 12'hd9c;
        src44 <= 12'h224;
        src45 <= 12'h6e2;
        src46 <= 12'h5b5;
        src47 <= 12'hff7;
        src48 <= 12'hcab;
        src49 <= 12'h782;
        src50 <= 12'h8c5;
        src51 <= 12'h60f;
        src52 <= 12'h6e6;
        src53 <= 12'ha4a;
        src54 <= 12'he03;
        src55 <= 12'hba3;
        src56 <= 12'he63;
        src57 <= 12'h940;
        src58 <= 12'h9;
        src59 <= 12'h129;
        src60 <= 12'h2e8;
        src61 <= 12'hb39;
        src62 <= 12'h17c;
        src63 <= 12'hcf3;
        src64 <= 12'h7a;
        src65 <= 12'h2b4;
        src66 <= 12'hca7;
        src67 <= 12'h45c;
        src68 <= 12'ha26;
        src69 <= 12'h331;
        src70 <= 12'h981;
        src71 <= 12'ha7;
        src72 <= 12'hc19;
        src73 <= 12'h9da;
        src74 <= 12'hec9;
        src75 <= 12'hd01;
        src76 <= 12'hd1e;
        src77 <= 12'hefb;
        src78 <= 12'hd8e;
        src79 <= 12'h4b;
        src80 <= 12'h828;
        src81 <= 12'h684;
        src82 <= 12'h7e9;
        src83 <= 12'h27;
        src84 <= 12'h907;
        src85 <= 12'h595;
        src86 <= 12'hdff;
        src87 <= 12'hd45;
        src88 <= 12'h38d;
        src89 <= 12'hcfb;
        src90 <= 12'had1;
        src91 <= 12'hfe5;
        src92 <= 12'hb0d;
        src93 <= 12'h2a4;
        src94 <= 12'h544;
        src95 <= 12'hcbc;
        src96 <= 12'h69e;
        src97 <= 12'hc5c;
        src98 <= 12'h6f7;
        src99 <= 12'h73;
        src100 <= 12'hfed;
        src101 <= 12'h97c;
        src102 <= 12'h990;
        src103 <= 12'h13d;
        src104 <= 12'h7b;
        src105 <= 12'ha85;
        src106 <= 12'h764;
        src107 <= 12'h7f8;
        src108 <= 12'h258;
        src109 <= 12'h376;
        src110 <= 12'hc46;
        src111 <= 12'h889;
        src112 <= 12'h917;
        src113 <= 12'h514;
        src114 <= 12'hb41;
        src115 <= 12'hee2;
        src116 <= 12'hca0;
        src117 <= 12'hb59;
        src118 <= 12'h7a7;
        src119 <= 12'h61d;
        src120 <= 12'h362;
        src121 <= 12'h3f8;
        src122 <= 12'h322;
        src123 <= 12'h8ce;
        src124 <= 12'hfb;
        src125 <= 12'h465;
        src126 <= 12'hfa8;
        src127 <= 12'hdb3;
        src128 <= 12'h3b0;
        src129 <= 12'h3cb;
        src130 <= 12'ha71;
        src131 <= 12'h8aa;
        src132 <= 12'ha81;
        src133 <= 12'h794;
        src134 <= 12'h74a;
        src135 <= 12'h4a3;
        src136 <= 12'hbd6;
        src137 <= 12'h897;
        src138 <= 12'hcbb;
        src139 <= 12'h8d0;
        src140 <= 12'h36;
        src141 <= 12'hb54;
        src142 <= 12'h669;
        src143 <= 12'he76;
        src144 <= 12'h16b;
        src145 <= 12'he4f;
        src146 <= 12'h22;
        src147 <= 12'h25c;
        src148 <= 12'h9;
        src149 <= 12'h273;
        src150 <= 12'hae8;
        src151 <= 12'hc3;
        src152 <= 12'he70;
        src153 <= 12'h36e;
        src154 <= 12'hb9c;
        src155 <= 12'h5ad;
        src156 <= 12'hce5;
        src157 <= 12'h8f2;
        src158 <= 12'h252;
        src159 <= 12'hf4f;
        src160 <= 12'hb3f;
        src161 <= 12'hea8;
        src162 <= 12'ha75;
        src163 <= 12'hfa1;
        src164 <= 12'hb9a;
        src165 <= 12'hac4;
        src166 <= 12'hec6;
        src167 <= 12'hf93;
        src168 <= 12'h255;
        src169 <= 12'h9f5;
        src170 <= 12'h37e;
        src171 <= 12'h305;
        src172 <= 12'ha0b;
        src173 <= 12'ha87;
        src174 <= 12'hd44;
        src175 <= 12'hd1;
        src176 <= 12'h706;
        src177 <= 12'h9b3;
        src178 <= 12'hc6d;
        src179 <= 12'h95a;
        src180 <= 12'he47;
        src181 <= 12'h1b2;
        src182 <= 12'h8f8;
        src183 <= 12'ha69;
        src184 <= 12'h1c1;
        src185 <= 12'h535;
        src186 <= 12'h44e;
        src187 <= 12'h652;
        src188 <= 12'h26e;
        exp <= 20'h5dc4c;
        #1
        src0 <= 12'h342;
        src1 <= 12'h855;
        src2 <= 12'h61d;
        src3 <= 12'h183;
        src4 <= 12'h8e1;
        src5 <= 12'hdd6;
        src6 <= 12'h58c;
        src7 <= 12'h16c;
        src8 <= 12'h3a9;
        src9 <= 12'h472;
        src10 <= 12'hf4f;
        src11 <= 12'h62c;
        src12 <= 12'h835;
        src13 <= 12'hc2;
        src14 <= 12'he7e;
        src15 <= 12'hec1;
        src16 <= 12'h6b1;
        src17 <= 12'heb7;
        src18 <= 12'h376;
        src19 <= 12'hc88;
        src20 <= 12'h942;
        src21 <= 12'hbb;
        src22 <= 12'h981;
        src23 <= 12'h8d0;
        src24 <= 12'ha58;
        src25 <= 12'h453;
        src26 <= 12'h7fe;
        src27 <= 12'ha1;
        src28 <= 12'ha61;
        src29 <= 12'h7e7;
        src30 <= 12'he95;
        src31 <= 12'h6cb;
        src32 <= 12'h207;
        src33 <= 12'h185;
        src34 <= 12'h593;
        src35 <= 12'hc40;
        src36 <= 12'h698;
        src37 <= 12'hc8d;
        src38 <= 12'h995;
        src39 <= 12'h27;
        src40 <= 12'h944;
        src41 <= 12'h5f9;
        src42 <= 12'h754;
        src43 <= 12'h35a;
        src44 <= 12'h7f;
        src45 <= 12'hbfe;
        src46 <= 12'hded;
        src47 <= 12'hf0a;
        src48 <= 12'h80;
        src49 <= 12'hf1c;
        src50 <= 12'h55e;
        src51 <= 12'h7ed;
        src52 <= 12'h11f;
        src53 <= 12'ha13;
        src54 <= 12'he54;
        src55 <= 12'h46a;
        src56 <= 12'h5a0;
        src57 <= 12'h8b9;
        src58 <= 12'h339;
        src59 <= 12'h752;
        src60 <= 12'hc42;
        src61 <= 12'h2d5;
        src62 <= 12'h641;
        src63 <= 12'h197;
        src64 <= 12'h3;
        src65 <= 12'h324;
        src66 <= 12'he73;
        src67 <= 12'h161;
        src68 <= 12'habf;
        src69 <= 12'h8a8;
        src70 <= 12'h3a4;
        src71 <= 12'h89a;
        src72 <= 12'hc46;
        src73 <= 12'hd5d;
        src74 <= 12'h58;
        src75 <= 12'hff0;
        src76 <= 12'h2b2;
        src77 <= 12'hc32;
        src78 <= 12'h2ec;
        src79 <= 12'ha50;
        src80 <= 12'h2ff;
        src81 <= 12'h39d;
        src82 <= 12'h5bf;
        src83 <= 12'h63b;
        src84 <= 12'hef7;
        src85 <= 12'habf;
        src86 <= 12'hbdc;
        src87 <= 12'h1b5;
        src88 <= 12'hfd2;
        src89 <= 12'h774;
        src90 <= 12'h37b;
        src91 <= 12'h946;
        src92 <= 12'h2b8;
        src93 <= 12'hb8e;
        src94 <= 12'hb12;
        src95 <= 12'h901;
        src96 <= 12'h30e;
        src97 <= 12'h7a2;
        src98 <= 12'h5f1;
        src99 <= 12'h9b;
        src100 <= 12'hb1a;
        src101 <= 12'h1a0;
        src102 <= 12'h62;
        src103 <= 12'hc82;
        src104 <= 12'h334;
        src105 <= 12'hee2;
        src106 <= 12'h5dd;
        src107 <= 12'h831;
        src108 <= 12'h869;
        src109 <= 12'hd3f;
        src110 <= 12'hcf3;
        src111 <= 12'hd8;
        src112 <= 12'h28;
        src113 <= 12'h67b;
        src114 <= 12'h2a4;
        src115 <= 12'h9d3;
        src116 <= 12'h2c7;
        src117 <= 12'h42b;
        src118 <= 12'h674;
        src119 <= 12'h63e;
        src120 <= 12'h974;
        src121 <= 12'h68d;
        src122 <= 12'he5c;
        src123 <= 12'h1f2;
        src124 <= 12'h44a;
        src125 <= 12'ha94;
        src126 <= 12'hc9a;
        src127 <= 12'hfe9;
        src128 <= 12'h939;
        src129 <= 12'h92e;
        src130 <= 12'hcd7;
        src131 <= 12'hc01;
        src132 <= 12'h5db;
        src133 <= 12'hf2;
        src134 <= 12'hd22;
        src135 <= 12'h295;
        src136 <= 12'haa8;
        src137 <= 12'hc2b;
        src138 <= 12'h419;
        src139 <= 12'h871;
        src140 <= 12'h3c7;
        src141 <= 12'hf0b;
        src142 <= 12'h43a;
        src143 <= 12'h3c1;
        src144 <= 12'h8b5;
        src145 <= 12'hbb4;
        src146 <= 12'ha6e;
        src147 <= 12'h40f;
        src148 <= 12'ha2d;
        src149 <= 12'h174;
        src150 <= 12'h264;
        src151 <= 12'h54d;
        src152 <= 12'h5c9;
        src153 <= 12'h5d3;
        src154 <= 12'h5a9;
        src155 <= 12'h3c3;
        src156 <= 12'h4a1;
        src157 <= 12'hcfe;
        src158 <= 12'h141;
        src159 <= 12'h6b;
        src160 <= 12'h7d7;
        src161 <= 12'h836;
        src162 <= 12'h6cc;
        src163 <= 12'h414;
        src164 <= 12'h433;
        src165 <= 12'h4e3;
        src166 <= 12'haf4;
        src167 <= 12'h637;
        src168 <= 12'hab8;
        src169 <= 12'h996;
        src170 <= 12'h563;
        src171 <= 12'h980;
        src172 <= 12'h702;
        src173 <= 12'h8ff;
        src174 <= 12'hf27;
        src175 <= 12'h622;
        src176 <= 12'he45;
        src177 <= 12'h46a;
        src178 <= 12'hbc0;
        src179 <= 12'h666;
        src180 <= 12'hb95;
        src181 <= 12'ha6d;
        src182 <= 12'h723;
        src183 <= 12'h3a5;
        src184 <= 12'h462;
        src185 <= 12'hd50;
        src186 <= 12'hfae;
        src187 <= 12'h79f;
        src188 <= 12'h518;
        exp <= 20'h57f3f;
        #1
        src0 <= 12'hfd6;
        src1 <= 12'hdaa;
        src2 <= 12'h9ec;
        src3 <= 12'hc57;
        src4 <= 12'h85e;
        src5 <= 12'ha09;
        src6 <= 12'hf0a;
        src7 <= 12'h543;
        src8 <= 12'h1b4;
        src9 <= 12'h63b;
        src10 <= 12'h9a3;
        src11 <= 12'hd3b;
        src12 <= 12'h6ea;
        src13 <= 12'h295;
        src14 <= 12'hdfa;
        src15 <= 12'h723;
        src16 <= 12'h161;
        src17 <= 12'h65b;
        src18 <= 12'h4eb;
        src19 <= 12'h523;
        src20 <= 12'h943;
        src21 <= 12'h58a;
        src22 <= 12'hfe0;
        src23 <= 12'h212;
        src24 <= 12'hec0;
        src25 <= 12'hee1;
        src26 <= 12'h3f5;
        src27 <= 12'h311;
        src28 <= 12'h987;
        src29 <= 12'h4dc;
        src30 <= 12'he7a;
        src31 <= 12'h4c0;
        src32 <= 12'h251;
        src33 <= 12'hb89;
        src34 <= 12'had7;
        src35 <= 12'h833;
        src36 <= 12'hb39;
        src37 <= 12'hac4;
        src38 <= 12'hb40;
        src39 <= 12'hee9;
        src40 <= 12'h1dc;
        src41 <= 12'h546;
        src42 <= 12'hfbf;
        src43 <= 12'hfd;
        src44 <= 12'h3c4;
        src45 <= 12'h786;
        src46 <= 12'h8f6;
        src47 <= 12'h7d6;
        src48 <= 12'h199;
        src49 <= 12'h5bc;
        src50 <= 12'he2;
        src51 <= 12'h543;
        src52 <= 12'h6dd;
        src53 <= 12'h496;
        src54 <= 12'h34a;
        src55 <= 12'haaf;
        src56 <= 12'h308;
        src57 <= 12'hc86;
        src58 <= 12'h581;
        src59 <= 12'hd24;
        src60 <= 12'hceb;
        src61 <= 12'h8f9;
        src62 <= 12'h64c;
        src63 <= 12'he67;
        src64 <= 12'hdc;
        src65 <= 12'h3cc;
        src66 <= 12'ha14;
        src67 <= 12'ha66;
        src68 <= 12'h6e7;
        src69 <= 12'h6cf;
        src70 <= 12'h38d;
        src71 <= 12'hf0a;
        src72 <= 12'h117;
        src73 <= 12'h1fc;
        src74 <= 12'h4d;
        src75 <= 12'h2bd;
        src76 <= 12'h6b7;
        src77 <= 12'hd32;
        src78 <= 12'hb9;
        src79 <= 12'hcd6;
        src80 <= 12'h4b8;
        src81 <= 12'h157;
        src82 <= 12'h651;
        src83 <= 12'heb3;
        src84 <= 12'h40b;
        src85 <= 12'hd01;
        src86 <= 12'h392;
        src87 <= 12'h78e;
        src88 <= 12'h885;
        src89 <= 12'h15a;
        src90 <= 12'hc25;
        src91 <= 12'h903;
        src92 <= 12'he68;
        src93 <= 12'h721;
        src94 <= 12'h2ad;
        src95 <= 12'hcfc;
        src96 <= 12'hbb8;
        src97 <= 12'hb77;
        src98 <= 12'h270;
        src99 <= 12'h3ff;
        src100 <= 12'hd8;
        src101 <= 12'hb4a;
        src102 <= 12'hef7;
        src103 <= 12'h15f;
        src104 <= 12'hd4c;
        src105 <= 12'hddd;
        src106 <= 12'h688;
        src107 <= 12'h487;
        src108 <= 12'hf0e;
        src109 <= 12'h6f;
        src110 <= 12'h2c9;
        src111 <= 12'h14f;
        src112 <= 12'hf08;
        src113 <= 12'h1f3;
        src114 <= 12'h4b1;
        src115 <= 12'h43a;
        src116 <= 12'h3a7;
        src117 <= 12'h89b;
        src118 <= 12'ha3e;
        src119 <= 12'h1cc;
        src120 <= 12'h8c3;
        src121 <= 12'hded;
        src122 <= 12'h694;
        src123 <= 12'h809;
        src124 <= 12'h8e1;
        src125 <= 12'h4a8;
        src126 <= 12'h4e8;
        src127 <= 12'hb22;
        src128 <= 12'h201;
        src129 <= 12'hb4f;
        src130 <= 12'h8f6;
        src131 <= 12'h46b;
        src132 <= 12'h8e3;
        src133 <= 12'hd1c;
        src134 <= 12'h21b;
        src135 <= 12'h6e7;
        src136 <= 12'hc35;
        src137 <= 12'hf23;
        src138 <= 12'h37d;
        src139 <= 12'h175;
        src140 <= 12'h45b;
        src141 <= 12'hec6;
        src142 <= 12'h330;
        src143 <= 12'h545;
        src144 <= 12'h615;
        src145 <= 12'he36;
        src146 <= 12'h4d8;
        src147 <= 12'ha3d;
        src148 <= 12'h5ff;
        src149 <= 12'h306;
        src150 <= 12'haf;
        src151 <= 12'hc8e;
        src152 <= 12'hb89;
        src153 <= 12'h7a1;
        src154 <= 12'he7a;
        src155 <= 12'h5fa;
        src156 <= 12'hb59;
        src157 <= 12'h581;
        src158 <= 12'h83f;
        src159 <= 12'h91e;
        src160 <= 12'h1fa;
        src161 <= 12'h653;
        src162 <= 12'hb8f;
        src163 <= 12'h6dd;
        src164 <= 12'hf60;
        src165 <= 12'h888;
        src166 <= 12'h59c;
        src167 <= 12'h5b6;
        src168 <= 12'h151;
        src169 <= 12'h191;
        src170 <= 12'h158;
        src171 <= 12'hd91;
        src172 <= 12'h479;
        src173 <= 12'h3f5;
        src174 <= 12'hc3f;
        src175 <= 12'h3cb;
        src176 <= 12'hcb4;
        src177 <= 12'hbb;
        src178 <= 12'ha90;
        src179 <= 12'he6;
        src180 <= 12'h987;
        src181 <= 12'h2a2;
        src182 <= 12'h35a;
        src183 <= 12'h4a5;
        src184 <= 12'hbf4;
        src185 <= 12'h445;
        src186 <= 12'h717;
        src187 <= 12'hf12;
        src188 <= 12'hbf7;
        exp <= 20'h58f71;
        #1
        src0 <= 12'ha1b;
        src1 <= 12'h8f8;
        src2 <= 12'he32;
        src3 <= 12'h2cf;
        src4 <= 12'hbc4;
        src5 <= 12'h71c;
        src6 <= 12'hc4a;
        src7 <= 12'h113;
        src8 <= 12'hcea;
        src9 <= 12'hf74;
        src10 <= 12'h1a;
        src11 <= 12'h6af;
        src12 <= 12'h730;
        src13 <= 12'hab0;
        src14 <= 12'ha41;
        src15 <= 12'hba0;
        src16 <= 12'h2e8;
        src17 <= 12'hee6;
        src18 <= 12'h422;
        src19 <= 12'h6c3;
        src20 <= 12'h1e0;
        src21 <= 12'h8b3;
        src22 <= 12'h558;
        src23 <= 12'h336;
        src24 <= 12'hed1;
        src25 <= 12'h515;
        src26 <= 12'h83f;
        src27 <= 12'h3e3;
        src28 <= 12'h496;
        src29 <= 12'hd5d;
        src30 <= 12'hbd8;
        src31 <= 12'hb44;
        src32 <= 12'ha67;
        src33 <= 12'h97d;
        src34 <= 12'h84f;
        src35 <= 12'hf2b;
        src36 <= 12'ha09;
        src37 <= 12'h865;
        src38 <= 12'he88;
        src39 <= 12'h9cb;
        src40 <= 12'ha72;
        src41 <= 12'h558;
        src42 <= 12'h21b;
        src43 <= 12'hf37;
        src44 <= 12'h880;
        src45 <= 12'hdf9;
        src46 <= 12'h316;
        src47 <= 12'h9cf;
        src48 <= 12'heef;
        src49 <= 12'h376;
        src50 <= 12'h9dc;
        src51 <= 12'h33;
        src52 <= 12'hdb2;
        src53 <= 12'h7c6;
        src54 <= 12'he3a;
        src55 <= 12'hba5;
        src56 <= 12'heaf;
        src57 <= 12'hbd6;
        src58 <= 12'hca0;
        src59 <= 12'h2ce;
        src60 <= 12'h50b;
        src61 <= 12'hdf9;
        src62 <= 12'h9a1;
        src63 <= 12'h11a;
        src64 <= 12'ha35;
        src65 <= 12'hb68;
        src66 <= 12'h2d6;
        src67 <= 12'h301;
        src68 <= 12'hea3;
        src69 <= 12'he2f;
        src70 <= 12'h393;
        src71 <= 12'hed2;
        src72 <= 12'h1e3;
        src73 <= 12'h713;
        src74 <= 12'he6;
        src75 <= 12'he25;
        src76 <= 12'ha1e;
        src77 <= 12'hdf3;
        src78 <= 12'h839;
        src79 <= 12'h42f;
        src80 <= 12'h2e7;
        src81 <= 12'hf61;
        src82 <= 12'hf85;
        src83 <= 12'hb73;
        src84 <= 12'h8d4;
        src85 <= 12'h4fe;
        src86 <= 12'h86a;
        src87 <= 12'hcac;
        src88 <= 12'h16e;
        src89 <= 12'h85a;
        src90 <= 12'h462;
        src91 <= 12'he25;
        src92 <= 12'hcb9;
        src93 <= 12'ha29;
        src94 <= 12'h220;
        src95 <= 12'h70d;
        src96 <= 12'h405;
        src97 <= 12'h99d;
        src98 <= 12'hc95;
        src99 <= 12'hf4a;
        src100 <= 12'h125;
        src101 <= 12'h18a;
        src102 <= 12'h612;
        src103 <= 12'h46b;
        src104 <= 12'he6f;
        src105 <= 12'h536;
        src106 <= 12'haba;
        src107 <= 12'h446;
        src108 <= 12'h67f;
        src109 <= 12'hfb9;
        src110 <= 12'h76a;
        src111 <= 12'hf52;
        src112 <= 12'he67;
        src113 <= 12'hb52;
        src114 <= 12'hcfc;
        src115 <= 12'h557;
        src116 <= 12'h3c9;
        src117 <= 12'hb1e;
        src118 <= 12'hbb8;
        src119 <= 12'hd16;
        src120 <= 12'hf75;
        src121 <= 12'h757;
        src122 <= 12'h6b7;
        src123 <= 12'h679;
        src124 <= 12'hf06;
        src125 <= 12'hbb4;
        src126 <= 12'hec;
        src127 <= 12'h13b;
        src128 <= 12'he31;
        src129 <= 12'h911;
        src130 <= 12'h6cf;
        src131 <= 12'h2c5;
        src132 <= 12'h5ae;
        src133 <= 12'hc3c;
        src134 <= 12'haf0;
        src135 <= 12'h3e5;
        src136 <= 12'hfa1;
        src137 <= 12'hba0;
        src138 <= 12'hebd;
        src139 <= 12'hb17;
        src140 <= 12'hc26;
        src141 <= 12'h474;
        src142 <= 12'h81b;
        src143 <= 12'h1dc;
        src144 <= 12'he8d;
        src145 <= 12'h88c;
        src146 <= 12'hce8;
        src147 <= 12'h842;
        src148 <= 12'h63b;
        src149 <= 12'h567;
        src150 <= 12'hcb7;
        src151 <= 12'ha91;
        src152 <= 12'ha93;
        src153 <= 12'h4d9;
        src154 <= 12'hfab;
        src155 <= 12'hf1d;
        src156 <= 12'h84a;
        src157 <= 12'h2a3;
        src158 <= 12'h271;
        src159 <= 12'ha52;
        src160 <= 12'h8c1;
        src161 <= 12'h250;
        src162 <= 12'hb3;
        src163 <= 12'h909;
        src164 <= 12'h4b1;
        src165 <= 12'h469;
        src166 <= 12'hacd;
        src167 <= 12'h262;
        src168 <= 12'h74;
        src169 <= 12'hae9;
        src170 <= 12'ha91;
        src171 <= 12'h936;
        src172 <= 12'hbcb;
        src173 <= 12'h8e;
        src174 <= 12'ha6;
        src175 <= 12'h3e3;
        src176 <= 12'h737;
        src177 <= 12'he63;
        src178 <= 12'h9f;
        src179 <= 12'hd90;
        src180 <= 12'h18f;
        src181 <= 12'h815;
        src182 <= 12'hbe9;
        src183 <= 12'h5a6;
        src184 <= 12'h8e9;
        src185 <= 12'hbc7;
        src186 <= 12'h545;
        src187 <= 12'ha59;
        src188 <= 12'hfa3;
        exp <= 20'h6591e;
        #1
        src0 <= 12'hab3;
        src1 <= 12'h854;
        src2 <= 12'h3d3;
        src3 <= 12'h633;
        src4 <= 12'h389;
        src5 <= 12'h25a;
        src6 <= 12'h87d;
        src7 <= 12'h63c;
        src8 <= 12'hd85;
        src9 <= 12'h63;
        src10 <= 12'h5bf;
        src11 <= 12'h25;
        src12 <= 12'hf64;
        src13 <= 12'h8a6;
        src14 <= 12'h625;
        src15 <= 12'h173;
        src16 <= 12'h1a6;
        src17 <= 12'hac5;
        src18 <= 12'hdd1;
        src19 <= 12'h7d6;
        src20 <= 12'h5f4;
        src21 <= 12'hdd8;
        src22 <= 12'hc20;
        src23 <= 12'h4c7;
        src24 <= 12'h8f4;
        src25 <= 12'h7f8;
        src26 <= 12'h88f;
        src27 <= 12'ha33;
        src28 <= 12'ha0d;
        src29 <= 12'hb20;
        src30 <= 12'h34d;
        src31 <= 12'h2a0;
        src32 <= 12'h48e;
        src33 <= 12'hd7b;
        src34 <= 12'he98;
        src35 <= 12'h679;
        src36 <= 12'hfaf;
        src37 <= 12'h6ff;
        src38 <= 12'hdb4;
        src39 <= 12'h243;
        src40 <= 12'h3d8;
        src41 <= 12'h390;
        src42 <= 12'h64e;
        src43 <= 12'h580;
        src44 <= 12'h12;
        src45 <= 12'hb0f;
        src46 <= 12'hc1c;
        src47 <= 12'hcd5;
        src48 <= 12'hdd8;
        src49 <= 12'h9af;
        src50 <= 12'h4ac;
        src51 <= 12'hd64;
        src52 <= 12'h4e;
        src53 <= 12'hbb4;
        src54 <= 12'h4fe;
        src55 <= 12'hba9;
        src56 <= 12'hca7;
        src57 <= 12'h1b7;
        src58 <= 12'h280;
        src59 <= 12'hc8b;
        src60 <= 12'ha9a;
        src61 <= 12'h8e3;
        src62 <= 12'he88;
        src63 <= 12'h16;
        src64 <= 12'hef4;
        src65 <= 12'h81c;
        src66 <= 12'hc55;
        src67 <= 12'hf0b;
        src68 <= 12'h298;
        src69 <= 12'h3ff;
        src70 <= 12'h83d;
        src71 <= 12'h703;
        src72 <= 12'h172;
        src73 <= 12'h1e5;
        src74 <= 12'h441;
        src75 <= 12'hcbb;
        src76 <= 12'h806;
        src77 <= 12'hec3;
        src78 <= 12'ha9b;
        src79 <= 12'h22f;
        src80 <= 12'h804;
        src81 <= 12'h985;
        src82 <= 12'hce0;
        src83 <= 12'h914;
        src84 <= 12'he8c;
        src85 <= 12'h62b;
        src86 <= 12'h531;
        src87 <= 12'h4b8;
        src88 <= 12'hf3d;
        src89 <= 12'hea2;
        src90 <= 12'h84f;
        src91 <= 12'hf6e;
        src92 <= 12'h95e;
        src93 <= 12'h279;
        src94 <= 12'hf9e;
        src95 <= 12'h297;
        src96 <= 12'h7e9;
        src97 <= 12'hf32;
        src98 <= 12'h2bb;
        src99 <= 12'h4e5;
        src100 <= 12'hf2f;
        src101 <= 12'h4a5;
        src102 <= 12'h6da;
        src103 <= 12'h38a;
        src104 <= 12'h58;
        src105 <= 12'h4a7;
        src106 <= 12'h7ed;
        src107 <= 12'h8da;
        src108 <= 12'h513;
        src109 <= 12'h750;
        src110 <= 12'h339;
        src111 <= 12'hafd;
        src112 <= 12'h6b1;
        src113 <= 12'he37;
        src114 <= 12'h160;
        src115 <= 12'haca;
        src116 <= 12'h693;
        src117 <= 12'hc23;
        src118 <= 12'hb34;
        src119 <= 12'h941;
        src120 <= 12'hc04;
        src121 <= 12'hea6;
        src122 <= 12'h2cf;
        src123 <= 12'hdd4;
        src124 <= 12'hd55;
        src125 <= 12'h8c5;
        src126 <= 12'ha50;
        src127 <= 12'hb8a;
        src128 <= 12'h437;
        src129 <= 12'hc25;
        src130 <= 12'h2d8;
        src131 <= 12'hfe1;
        src132 <= 12'h852;
        src133 <= 12'hb75;
        src134 <= 12'h8ff;
        src135 <= 12'heb5;
        src136 <= 12'h5ce;
        src137 <= 12'h6f6;
        src138 <= 12'hf49;
        src139 <= 12'h8a2;
        src140 <= 12'hc81;
        src141 <= 12'hb2f;
        src142 <= 12'h7da;
        src143 <= 12'h849;
        src144 <= 12'h5e6;
        src145 <= 12'ha8e;
        src146 <= 12'h553;
        src147 <= 12'he0f;
        src148 <= 12'hcbe;
        src149 <= 12'hcbe;
        src150 <= 12'h8e5;
        src151 <= 12'h630;
        src152 <= 12'hf10;
        src153 <= 12'ha3e;
        src154 <= 12'h9e4;
        src155 <= 12'he4d;
        src156 <= 12'hd3e;
        src157 <= 12'h3e2;
        src158 <= 12'hf0;
        src159 <= 12'h57f;
        src160 <= 12'h95a;
        src161 <= 12'haa4;
        src162 <= 12'hd07;
        src163 <= 12'ha9c;
        src164 <= 12'h3a9;
        src165 <= 12'hebe;
        src166 <= 12'h893;
        src167 <= 12'ha6b;
        src168 <= 12'h4d7;
        src169 <= 12'h751;
        src170 <= 12'he0c;
        src171 <= 12'ha7a;
        src172 <= 12'hcd;
        src173 <= 12'h4d3;
        src174 <= 12'hfc4;
        src175 <= 12'h23;
        src176 <= 12'hda4;
        src177 <= 12'h555;
        src178 <= 12'hce1;
        src179 <= 12'hace;
        src180 <= 12'h2a3;
        src181 <= 12'hf8c;
        src182 <= 12'haac;
        src183 <= 12'h29b;
        src184 <= 12'h7ee;
        src185 <= 12'h395;
        src186 <= 12'hc12;
        src187 <= 12'hfbf;
        src188 <= 12'hd00;
        exp <= 20'h65665;
        #1
        src0 <= 12'h834;
        src1 <= 12'h17;
        src2 <= 12'h8b7;
        src3 <= 12'hb3b;
        src4 <= 12'hf9c;
        src5 <= 12'hf7b;
        src6 <= 12'h150;
        src7 <= 12'h436;
        src8 <= 12'h383;
        src9 <= 12'h584;
        src10 <= 12'h8e;
        src11 <= 12'h3d1;
        src12 <= 12'hf6a;
        src13 <= 12'h7ea;
        src14 <= 12'h85;
        src15 <= 12'h6c2;
        src16 <= 12'h5c4;
        src17 <= 12'h454;
        src18 <= 12'h5ce;
        src19 <= 12'h869;
        src20 <= 12'h60a;
        src21 <= 12'h244;
        src22 <= 12'h72;
        src23 <= 12'hb5;
        src24 <= 12'h342;
        src25 <= 12'h882;
        src26 <= 12'h847;
        src27 <= 12'hdc;
        src28 <= 12'hd61;
        src29 <= 12'hd80;
        src30 <= 12'hd16;
        src31 <= 12'hc43;
        src32 <= 12'h758;
        src33 <= 12'h613;
        src34 <= 12'h2d;
        src35 <= 12'h1f2;
        src36 <= 12'h8fa;
        src37 <= 12'h370;
        src38 <= 12'hde8;
        src39 <= 12'h8b5;
        src40 <= 12'h5ea;
        src41 <= 12'h62e;
        src42 <= 12'h78d;
        src43 <= 12'h43;
        src44 <= 12'h998;
        src45 <= 12'h551;
        src46 <= 12'h793;
        src47 <= 12'he9c;
        src48 <= 12'h7b4;
        src49 <= 12'hb4c;
        src50 <= 12'hd7b;
        src51 <= 12'hc5e;
        src52 <= 12'h6d1;
        src53 <= 12'h56;
        src54 <= 12'h99e;
        src55 <= 12'h748;
        src56 <= 12'h56c;
        src57 <= 12'h50b;
        src58 <= 12'h174;
        src59 <= 12'h821;
        src60 <= 12'h272;
        src61 <= 12'h367;
        src62 <= 12'h717;
        src63 <= 12'h665;
        src64 <= 12'h33f;
        src65 <= 12'hb1c;
        src66 <= 12'h4c9;
        src67 <= 12'h613;
        src68 <= 12'he55;
        src69 <= 12'h39c;
        src70 <= 12'h4c;
        src71 <= 12'h107;
        src72 <= 12'h1dd;
        src73 <= 12'h9e0;
        src74 <= 12'h721;
        src75 <= 12'hcb0;
        src76 <= 12'h76;
        src77 <= 12'hc2c;
        src78 <= 12'hd28;
        src79 <= 12'h391;
        src80 <= 12'he69;
        src81 <= 12'hd6;
        src82 <= 12'h1de;
        src83 <= 12'hc;
        src84 <= 12'hacc;
        src85 <= 12'hc23;
        src86 <= 12'hee8;
        src87 <= 12'h54c;
        src88 <= 12'h4a9;
        src89 <= 12'h981;
        src90 <= 12'h180;
        src91 <= 12'h91;
        src92 <= 12'hacd;
        src93 <= 12'he52;
        src94 <= 12'h2fc;
        src95 <= 12'hfc1;
        src96 <= 12'heb;
        src97 <= 12'h703;
        src98 <= 12'ha4a;
        src99 <= 12'h5f2;
        src100 <= 12'hfb9;
        src101 <= 12'h7c;
        src102 <= 12'h27a;
        src103 <= 12'had9;
        src104 <= 12'ha64;
        src105 <= 12'h99c;
        src106 <= 12'hd2d;
        src107 <= 12'hb95;
        src108 <= 12'hb1e;
        src109 <= 12'h393;
        src110 <= 12'hf19;
        src111 <= 12'hb82;
        src112 <= 12'hc62;
        src113 <= 12'hdc5;
        src114 <= 12'h889;
        src115 <= 12'h66b;
        src116 <= 12'h32a;
        src117 <= 12'h886;
        src118 <= 12'h15c;
        src119 <= 12'h535;
        src120 <= 12'ha43;
        src121 <= 12'hdf2;
        src122 <= 12'h879;
        src123 <= 12'h44a;
        src124 <= 12'h1c;
        src125 <= 12'hc20;
        src126 <= 12'h3c8;
        src127 <= 12'h5be;
        src128 <= 12'h96f;
        src129 <= 12'h7d7;
        src130 <= 12'hb20;
        src131 <= 12'h212;
        src132 <= 12'h586;
        src133 <= 12'h30f;
        src134 <= 12'hc6e;
        src135 <= 12'hedf;
        src136 <= 12'ha6d;
        src137 <= 12'h6e0;
        src138 <= 12'hd52;
        src139 <= 12'h375;
        src140 <= 12'h9e2;
        src141 <= 12'h9a9;
        src142 <= 12'hc20;
        src143 <= 12'h208;
        src144 <= 12'h75a;
        src145 <= 12'h267;
        src146 <= 12'he5b;
        src147 <= 12'hc54;
        src148 <= 12'h49c;
        src149 <= 12'hff3;
        src150 <= 12'hd44;
        src151 <= 12'hd11;
        src152 <= 12'hc3d;
        src153 <= 12'h744;
        src154 <= 12'h9a1;
        src155 <= 12'h7da;
        src156 <= 12'h51a;
        src157 <= 12'ha4e;
        src158 <= 12'hd78;
        src159 <= 12'hf6d;
        src160 <= 12'hb02;
        src161 <= 12'h713;
        src162 <= 12'hf02;
        src163 <= 12'h95;
        src164 <= 12'h92b;
        src165 <= 12'hdb9;
        src166 <= 12'h7c5;
        src167 <= 12'hb95;
        src168 <= 12'h978;
        src169 <= 12'h855;
        src170 <= 12'hb0b;
        src171 <= 12'h80;
        src172 <= 12'h21c;
        src173 <= 12'h1d;
        src174 <= 12'h3c4;
        src175 <= 12'h130;
        src176 <= 12'hbb1;
        src177 <= 12'h2aa;
        src178 <= 12'h539;
        src179 <= 12'h9d0;
        src180 <= 12'hc07;
        src181 <= 12'hefb;
        src182 <= 12'hf67;
        src183 <= 12'h82c;
        src184 <= 12'h49f;
        src185 <= 12'ha18;
        src186 <= 12'hd3e;
        src187 <= 12'hed1;
        src188 <= 12'h6ba;
        exp <= 20'h5afdb;
        #1
        src0 <= 12'h5c9;
        src1 <= 12'hc3e;
        src2 <= 12'haa9;
        src3 <= 12'h55e;
        src4 <= 12'hfd2;
        src5 <= 12'h321;
        src6 <= 12'h54b;
        src7 <= 12'hc59;
        src8 <= 12'h66d;
        src9 <= 12'h2e2;
        src10 <= 12'h20f;
        src11 <= 12'h439;
        src12 <= 12'hcbf;
        src13 <= 12'h8bb;
        src14 <= 12'h7f3;
        src15 <= 12'h546;
        src16 <= 12'h94a;
        src17 <= 12'h407;
        src18 <= 12'hff8;
        src19 <= 12'h790;
        src20 <= 12'hbc;
        src21 <= 12'he13;
        src22 <= 12'hfb6;
        src23 <= 12'hfa;
        src24 <= 12'h10f;
        src25 <= 12'h784;
        src26 <= 12'hf2c;
        src27 <= 12'hf62;
        src28 <= 12'h572;
        src29 <= 12'h870;
        src30 <= 12'hf6;
        src31 <= 12'h75d;
        src32 <= 12'hcd7;
        src33 <= 12'hf1e;
        src34 <= 12'h7a6;
        src35 <= 12'hb50;
        src36 <= 12'h341;
        src37 <= 12'h362;
        src38 <= 12'h239;
        src39 <= 12'h7c7;
        src40 <= 12'hde9;
        src41 <= 12'hf83;
        src42 <= 12'hfba;
        src43 <= 12'h974;
        src44 <= 12'h71d;
        src45 <= 12'h596;
        src46 <= 12'hc6d;
        src47 <= 12'h136;
        src48 <= 12'hc88;
        src49 <= 12'h833;
        src50 <= 12'h34d;
        src51 <= 12'h4c;
        src52 <= 12'h7e3;
        src53 <= 12'hec3;
        src54 <= 12'h33a;
        src55 <= 12'ha58;
        src56 <= 12'hae4;
        src57 <= 12'h9c3;
        src58 <= 12'h332;
        src59 <= 12'had8;
        src60 <= 12'h2ba;
        src61 <= 12'hf63;
        src62 <= 12'h267;
        src63 <= 12'h140;
        src64 <= 12'h3d5;
        src65 <= 12'h670;
        src66 <= 12'hdc2;
        src67 <= 12'hbe8;
        src68 <= 12'hcd1;
        src69 <= 12'h553;
        src70 <= 12'h212;
        src71 <= 12'h316;
        src72 <= 12'he3a;
        src73 <= 12'haa2;
        src74 <= 12'h5fc;
        src75 <= 12'h45b;
        src76 <= 12'h47;
        src77 <= 12'h85f;
        src78 <= 12'h2eb;
        src79 <= 12'h1d1;
        src80 <= 12'h50e;
        src81 <= 12'h1a3;
        src82 <= 12'h27e;
        src83 <= 12'h4c0;
        src84 <= 12'h495;
        src85 <= 12'hc81;
        src86 <= 12'h52c;
        src87 <= 12'h3c2;
        src88 <= 12'h5ae;
        src89 <= 12'ha7a;
        src90 <= 12'he96;
        src91 <= 12'h49e;
        src92 <= 12'h346;
        src93 <= 12'h86b;
        src94 <= 12'ha4c;
        src95 <= 12'head;
        src96 <= 12'he91;
        src97 <= 12'h709;
        src98 <= 12'h984;
        src99 <= 12'ha71;
        src100 <= 12'hab3;
        src101 <= 12'h88a;
        src102 <= 12'hd2b;
        src103 <= 12'h7ad;
        src104 <= 12'hee6;
        src105 <= 12'h842;
        src106 <= 12'hea4;
        src107 <= 12'hae6;
        src108 <= 12'hea3;
        src109 <= 12'h537;
        src110 <= 12'ha8f;
        src111 <= 12'haab;
        src112 <= 12'ha5d;
        src113 <= 12'h78a;
        src114 <= 12'h1d2;
        src115 <= 12'h6e3;
        src116 <= 12'he8b;
        src117 <= 12'h75a;
        src118 <= 12'h36b;
        src119 <= 12'h90a;
        src120 <= 12'hf09;
        src121 <= 12'hb8b;
        src122 <= 12'hfbb;
        src123 <= 12'haf8;
        src124 <= 12'h2c7;
        src125 <= 12'h42d;
        src126 <= 12'h314;
        src127 <= 12'h647;
        src128 <= 12'h8f4;
        src129 <= 12'hba6;
        src130 <= 12'h813;
        src131 <= 12'h424;
        src132 <= 12'h7a2;
        src133 <= 12'h49e;
        src134 <= 12'h42;
        src135 <= 12'h270;
        src136 <= 12'h799;
        src137 <= 12'hc3b;
        src138 <= 12'hc1a;
        src139 <= 12'h5da;
        src140 <= 12'h541;
        src141 <= 12'h22e;
        src142 <= 12'h1e4;
        src143 <= 12'h1a;
        src144 <= 12'h6a8;
        src145 <= 12'haa9;
        src146 <= 12'h947;
        src147 <= 12'h61d;
        src148 <= 12'h8de;
        src149 <= 12'hf8c;
        src150 <= 12'h3f2;
        src151 <= 12'h36c;
        src152 <= 12'h627;
        src153 <= 12'hf1f;
        src154 <= 12'hcbf;
        src155 <= 12'h999;
        src156 <= 12'h85b;
        src157 <= 12'hb7a;
        src158 <= 12'h472;
        src159 <= 12'hdfb;
        src160 <= 12'h36d;
        src161 <= 12'hb68;
        src162 <= 12'h243;
        src163 <= 12'he15;
        src164 <= 12'h487;
        src165 <= 12'hb1f;
        src166 <= 12'h25;
        src167 <= 12'he2b;
        src168 <= 12'h6b2;
        src169 <= 12'h25e;
        src170 <= 12'hff8;
        src171 <= 12'h5b7;
        src172 <= 12'h9ce;
        src173 <= 12'hfba;
        src174 <= 12'h34b;
        src175 <= 12'h4a3;
        src176 <= 12'h2e0;
        src177 <= 12'h2eb;
        src178 <= 12'hc74;
        src179 <= 12'h8;
        src180 <= 12'hb13;
        src181 <= 12'hc56;
        src182 <= 12'hcd6;
        src183 <= 12'hdeb;
        src184 <= 12'h9a8;
        src185 <= 12'h756;
        src186 <= 12'hd3e;
        src187 <= 12'h664;
        src188 <= 12'h85d;
        exp <= 20'h5e9f6;
        #1
        src0 <= 12'h1e1;
        src1 <= 12'h56f;
        src2 <= 12'h57c;
        src3 <= 12'hf3c;
        src4 <= 12'h4f7;
        src5 <= 12'hab7;
        src6 <= 12'h791;
        src7 <= 12'hdc4;
        src8 <= 12'h131;
        src9 <= 12'h84b;
        src10 <= 12'h826;
        src11 <= 12'h5fe;
        src12 <= 12'h5b7;
        src13 <= 12'h36d;
        src14 <= 12'ha2d;
        src15 <= 12'h462;
        src16 <= 12'h32c;
        src17 <= 12'h3f3;
        src18 <= 12'h38c;
        src19 <= 12'h11f;
        src20 <= 12'h375;
        src21 <= 12'he44;
        src22 <= 12'h3f3;
        src23 <= 12'h8ee;
        src24 <= 12'h5ef;
        src25 <= 12'h284;
        src26 <= 12'h937;
        src27 <= 12'h671;
        src28 <= 12'h306;
        src29 <= 12'h8d5;
        src30 <= 12'hdc0;
        src31 <= 12'h886;
        src32 <= 12'h30f;
        src33 <= 12'h6ac;
        src34 <= 12'h898;
        src35 <= 12'hf2;
        src36 <= 12'h767;
        src37 <= 12'hefb;
        src38 <= 12'hf65;
        src39 <= 12'hef4;
        src40 <= 12'haac;
        src41 <= 12'h2f;
        src42 <= 12'hf85;
        src43 <= 12'hd1b;
        src44 <= 12'h415;
        src45 <= 12'hfde;
        src46 <= 12'h6a9;
        src47 <= 12'h399;
        src48 <= 12'hcbc;
        src49 <= 12'h6b5;
        src50 <= 12'hf38;
        src51 <= 12'haec;
        src52 <= 12'h3c;
        src53 <= 12'had2;
        src54 <= 12'h421;
        src55 <= 12'h86f;
        src56 <= 12'hbe1;
        src57 <= 12'h88;
        src58 <= 12'h162;
        src59 <= 12'hc7d;
        src60 <= 12'h5dd;
        src61 <= 12'h55d;
        src62 <= 12'hc8d;
        src63 <= 12'hec;
        src64 <= 12'he99;
        src65 <= 12'h4d7;
        src66 <= 12'hbc9;
        src67 <= 12'h739;
        src68 <= 12'hfe0;
        src69 <= 12'hd8d;
        src70 <= 12'h8f4;
        src71 <= 12'h360;
        src72 <= 12'h3dc;
        src73 <= 12'hb64;
        src74 <= 12'h692;
        src75 <= 12'h497;
        src76 <= 12'h86d;
        src77 <= 12'h7c9;
        src78 <= 12'h4e9;
        src79 <= 12'h63e;
        src80 <= 12'h887;
        src81 <= 12'h3a4;
        src82 <= 12'h604;
        src83 <= 12'h1ff;
        src84 <= 12'ha1f;
        src85 <= 12'h15a;
        src86 <= 12'ha69;
        src87 <= 12'he50;
        src88 <= 12'h140;
        src89 <= 12'hd67;
        src90 <= 12'h667;
        src91 <= 12'h7da;
        src92 <= 12'h25e;
        src93 <= 12'h55;
        src94 <= 12'h621;
        src95 <= 12'hb1a;
        src96 <= 12'h715;
        src97 <= 12'h719;
        src98 <= 12'h51a;
        src99 <= 12'h22f;
        src100 <= 12'h68b;
        src101 <= 12'h73d;
        src102 <= 12'h144;
        src103 <= 12'hfeb;
        src104 <= 12'hccf;
        src105 <= 12'hff7;
        src106 <= 12'hd05;
        src107 <= 12'ha6c;
        src108 <= 12'h1a1;
        src109 <= 12'h8d4;
        src110 <= 12'h4b;
        src111 <= 12'hc2e;
        src112 <= 12'hf9d;
        src113 <= 12'hdc8;
        src114 <= 12'h808;
        src115 <= 12'h631;
        src116 <= 12'h1ea;
        src117 <= 12'hd5f;
        src118 <= 12'h122;
        src119 <= 12'h515;
        src120 <= 12'h3dd;
        src121 <= 12'ha1d;
        src122 <= 12'hea4;
        src123 <= 12'h562;
        src124 <= 12'h444;
        src125 <= 12'h5aa;
        src126 <= 12'h598;
        src127 <= 12'h20f;
        src128 <= 12'h5a3;
        src129 <= 12'h7c7;
        src130 <= 12'hc0c;
        src131 <= 12'h479;
        src132 <= 12'hbee;
        src133 <= 12'haa8;
        src134 <= 12'h567;
        src135 <= 12'hf4d;
        src136 <= 12'h81f;
        src137 <= 12'hc54;
        src138 <= 12'h508;
        src139 <= 12'h3b6;
        src140 <= 12'h650;
        src141 <= 12'h7cb;
        src142 <= 12'h6b7;
        src143 <= 12'haff;
        src144 <= 12'haba;
        src145 <= 12'h879;
        src146 <= 12'h7eb;
        src147 <= 12'h946;
        src148 <= 12'h6a3;
        src149 <= 12'h9f2;
        src150 <= 12'h166;
        src151 <= 12'ha90;
        src152 <= 12'h168;
        src153 <= 12'ha02;
        src154 <= 12'h45;
        src155 <= 12'h591;
        src156 <= 12'haf2;
        src157 <= 12'hd6c;
        src158 <= 12'h643;
        src159 <= 12'hec1;
        src160 <= 12'hc4d;
        src161 <= 12'h2f;
        src162 <= 12'h5c7;
        src163 <= 12'h307;
        src164 <= 12'h835;
        src165 <= 12'h5e3;
        src166 <= 12'h396;
        src167 <= 12'h932;
        src168 <= 12'hb90;
        src169 <= 12'hece;
        src170 <= 12'hce6;
        src171 <= 12'h4a1;
        src172 <= 12'h18f;
        src173 <= 12'hd38;
        src174 <= 12'ha28;
        src175 <= 12'h3a3;
        src176 <= 12'h202;
        src177 <= 12'hfce;
        src178 <= 12'hf6f;
        src179 <= 12'he29;
        src180 <= 12'hef4;
        src181 <= 12'h2d2;
        src182 <= 12'h71e;
        src183 <= 12'hc37;
        src184 <= 12'h96d;
        src185 <= 12'h753;
        src186 <= 12'hb2f;
        src187 <= 12'h7b9;
        src188 <= 12'hcd3;
        exp <= 20'h5c1bc;
        #1
        src0 <= 12'h73f;
        src1 <= 12'h53c;
        src2 <= 12'h92b;
        src3 <= 12'h5ad;
        src4 <= 12'h660;
        src5 <= 12'hade;
        src6 <= 12'he44;
        src7 <= 12'h755;
        src8 <= 12'h6d9;
        src9 <= 12'h99;
        src10 <= 12'ha11;
        src11 <= 12'hdc5;
        src12 <= 12'he8c;
        src13 <= 12'he1b;
        src14 <= 12'hfb4;
        src15 <= 12'h155;
        src16 <= 12'hf65;
        src17 <= 12'h826;
        src18 <= 12'hfaf;
        src19 <= 12'h797;
        src20 <= 12'h9f9;
        src21 <= 12'h9d0;
        src22 <= 12'h611;
        src23 <= 12'h5e0;
        src24 <= 12'h281;
        src25 <= 12'ha92;
        src26 <= 12'ha7c;
        src27 <= 12'h475;
        src28 <= 12'h357;
        src29 <= 12'h608;
        src30 <= 12'h33a;
        src31 <= 12'h1fb;
        src32 <= 12'hb42;
        src33 <= 12'h4bd;
        src34 <= 12'h21a;
        src35 <= 12'h55f;
        src36 <= 12'hf4a;
        src37 <= 12'hdb3;
        src38 <= 12'h541;
        src39 <= 12'hc7c;
        src40 <= 12'h425;
        src41 <= 12'hfb0;
        src42 <= 12'he57;
        src43 <= 12'h676;
        src44 <= 12'hbe5;
        src45 <= 12'hda6;
        src46 <= 12'h298;
        src47 <= 12'h83a;
        src48 <= 12'h194;
        src49 <= 12'hee7;
        src50 <= 12'h244;
        src51 <= 12'h1cf;
        src52 <= 12'h16a;
        src53 <= 12'h5d1;
        src54 <= 12'hefb;
        src55 <= 12'h8d3;
        src56 <= 12'h7ee;
        src57 <= 12'hac8;
        src58 <= 12'h380;
        src59 <= 12'h906;
        src60 <= 12'h74a;
        src61 <= 12'h639;
        src62 <= 12'haa;
        src63 <= 12'hfcb;
        src64 <= 12'hcbe;
        src65 <= 12'hb7a;
        src66 <= 12'h17e;
        src67 <= 12'hdad;
        src68 <= 12'h3d6;
        src69 <= 12'he46;
        src70 <= 12'h477;
        src71 <= 12'h794;
        src72 <= 12'hb60;
        src73 <= 12'ha28;
        src74 <= 12'h937;
        src75 <= 12'h4d1;
        src76 <= 12'hd27;
        src77 <= 12'haaa;
        src78 <= 12'he67;
        src79 <= 12'h990;
        src80 <= 12'h406;
        src81 <= 12'hecd;
        src82 <= 12'he89;
        src83 <= 12'h881;
        src84 <= 12'h3ad;
        src85 <= 12'h22d;
        src86 <= 12'hccc;
        src87 <= 12'h3e;
        src88 <= 12'he36;
        src89 <= 12'he29;
        src90 <= 12'h384;
        src91 <= 12'h85a;
        src92 <= 12'h5df;
        src93 <= 12'hb1c;
        src94 <= 12'h126;
        src95 <= 12'h803;
        src96 <= 12'h440;
        src97 <= 12'h48c;
        src98 <= 12'hae7;
        src99 <= 12'he19;
        src100 <= 12'h59;
        src101 <= 12'h649;
        src102 <= 12'h2a0;
        src103 <= 12'hbf9;
        src104 <= 12'he51;
        src105 <= 12'hb30;
        src106 <= 12'h130;
        src107 <= 12'h85a;
        src108 <= 12'h247;
        src109 <= 12'h9b7;
        src110 <= 12'haba;
        src111 <= 12'h9f;
        src112 <= 12'he3f;
        src113 <= 12'h2d0;
        src114 <= 12'h596;
        src115 <= 12'h3b;
        src116 <= 12'had3;
        src117 <= 12'h20e;
        src118 <= 12'h291;
        src119 <= 12'hd31;
        src120 <= 12'h945;
        src121 <= 12'h6ce;
        src122 <= 12'h493;
        src123 <= 12'he79;
        src124 <= 12'hfbf;
        src125 <= 12'hef3;
        src126 <= 12'h32e;
        src127 <= 12'h6ed;
        src128 <= 12'h94c;
        src129 <= 12'h7d0;
        src130 <= 12'hc2a;
        src131 <= 12'h970;
        src132 <= 12'h734;
        src133 <= 12'h8f5;
        src134 <= 12'h779;
        src135 <= 12'h8e1;
        src136 <= 12'h3a2;
        src137 <= 12'h596;
        src138 <= 12'h89;
        src139 <= 12'hcf2;
        src140 <= 12'h799;
        src141 <= 12'h5d2;
        src142 <= 12'h111;
        src143 <= 12'he37;
        src144 <= 12'h8cd;
        src145 <= 12'h6c1;
        src146 <= 12'hc6d;
        src147 <= 12'h2dd;
        src148 <= 12'hd10;
        src149 <= 12'he5b;
        src150 <= 12'h14f;
        src151 <= 12'h388;
        src152 <= 12'hb43;
        src153 <= 12'h7d6;
        src154 <= 12'h2f0;
        src155 <= 12'h200;
        src156 <= 12'ha9b;
        src157 <= 12'hd79;
        src158 <= 12'h916;
        src159 <= 12'h76e;
        src160 <= 12'h631;
        src161 <= 12'h971;
        src162 <= 12'h5ff;
        src163 <= 12'h2dd;
        src164 <= 12'hecf;
        src165 <= 12'h90a;
        src166 <= 12'h3b2;
        src167 <= 12'h2ef;
        src168 <= 12'h33a;
        src169 <= 12'hf55;
        src170 <= 12'h51f;
        src171 <= 12'hf71;
        src172 <= 12'h678;
        src173 <= 12'hdce;
        src174 <= 12'h817;
        src175 <= 12'h8ee;
        src176 <= 12'h6fc;
        src177 <= 12'he79;
        src178 <= 12'hbe7;
        src179 <= 12'ha09;
        src180 <= 12'h6a8;
        src181 <= 12'h552;
        src182 <= 12'h469;
        src183 <= 12'h968;
        src184 <= 12'h65f;
        src185 <= 12'h299;
        src186 <= 12'h168;
        src187 <= 12'h663;
        src188 <= 12'h4c3;
        exp <= 20'h5ed8f;
        #1
        src0 <= 12'h90d;
        src1 <= 12'h882;
        src2 <= 12'h37c;
        src3 <= 12'hd65;
        src4 <= 12'hc10;
        src5 <= 12'hae8;
        src6 <= 12'h312;
        src7 <= 12'h3cc;
        src8 <= 12'h97d;
        src9 <= 12'ha55;
        src10 <= 12'hd04;
        src11 <= 12'hbf;
        src12 <= 12'h56e;
        src13 <= 12'hc88;
        src14 <= 12'hc17;
        src15 <= 12'he8b;
        src16 <= 12'ha9e;
        src17 <= 12'h9d7;
        src18 <= 12'h9cb;
        src19 <= 12'heca;
        src20 <= 12'hb43;
        src21 <= 12'hcf2;
        src22 <= 12'hc78;
        src23 <= 12'ha59;
        src24 <= 12'h9d3;
        src25 <= 12'h303;
        src26 <= 12'h415;
        src27 <= 12'h846;
        src28 <= 12'h6cd;
        src29 <= 12'hb0f;
        src30 <= 12'hcd5;
        src31 <= 12'h181;
        src32 <= 12'he77;
        src33 <= 12'h4b4;
        src34 <= 12'h270;
        src35 <= 12'hcfc;
        src36 <= 12'h754;
        src37 <= 12'h994;
        src38 <= 12'hd80;
        src39 <= 12'h9b2;
        src40 <= 12'hb53;
        src41 <= 12'hde1;
        src42 <= 12'h7a4;
        src43 <= 12'h7be;
        src44 <= 12'h9f8;
        src45 <= 12'h410;
        src46 <= 12'hddb;
        src47 <= 12'ha1;
        src48 <= 12'hce;
        src49 <= 12'h560;
        src50 <= 12'hc48;
        src51 <= 12'hb7c;
        src52 <= 12'h8a0;
        src53 <= 12'h7eb;
        src54 <= 12'hd55;
        src55 <= 12'he70;
        src56 <= 12'hc7;
        src57 <= 12'h152;
        src58 <= 12'h796;
        src59 <= 12'haee;
        src60 <= 12'h654;
        src61 <= 12'hc18;
        src62 <= 12'h386;
        src63 <= 12'h6d7;
        src64 <= 12'h6f6;
        src65 <= 12'h342;
        src66 <= 12'ha8a;
        src67 <= 12'h38c;
        src68 <= 12'hf28;
        src69 <= 12'hfba;
        src70 <= 12'h17f;
        src71 <= 12'hd4e;
        src72 <= 12'hd85;
        src73 <= 12'h4bf;
        src74 <= 12'hc18;
        src75 <= 12'hbde;
        src76 <= 12'h614;
        src77 <= 12'h9fe;
        src78 <= 12'h1f3;
        src79 <= 12'h9d5;
        src80 <= 12'h7b2;
        src81 <= 12'hec3;
        src82 <= 12'h600;
        src83 <= 12'h617;
        src84 <= 12'hd8f;
        src85 <= 12'ha7;
        src86 <= 12'h1b8;
        src87 <= 12'h2fd;
        src88 <= 12'hec0;
        src89 <= 12'h51e;
        src90 <= 12'h62a;
        src91 <= 12'h684;
        src92 <= 12'h2f4;
        src93 <= 12'hcd1;
        src94 <= 12'he8b;
        src95 <= 12'hb6a;
        src96 <= 12'h6b0;
        src97 <= 12'h2db;
        src98 <= 12'h803;
        src99 <= 12'h3d3;
        src100 <= 12'hbd8;
        src101 <= 12'hf27;
        src102 <= 12'h1a;
        src103 <= 12'hd14;
        src104 <= 12'h4c7;
        src105 <= 12'hb1b;
        src106 <= 12'he50;
        src107 <= 12'h3cc;
        src108 <= 12'he99;
        src109 <= 12'h5eb;
        src110 <= 12'h604;
        src111 <= 12'he68;
        src112 <= 12'he7f;
        src113 <= 12'h508;
        src114 <= 12'h559;
        src115 <= 12'h1;
        src116 <= 12'h9e1;
        src117 <= 12'h315;
        src118 <= 12'h88b;
        src119 <= 12'h8d1;
        src120 <= 12'h413;
        src121 <= 12'h90b;
        src122 <= 12'h5bd;
        src123 <= 12'hd38;
        src124 <= 12'h538;
        src125 <= 12'h962;
        src126 <= 12'he2b;
        src127 <= 12'hfdc;
        src128 <= 12'ha67;
        src129 <= 12'h422;
        src130 <= 12'h3f1;
        src131 <= 12'h1fa;
        src132 <= 12'h140;
        src133 <= 12'h273;
        src134 <= 12'hd1e;
        src135 <= 12'hb72;
        src136 <= 12'h810;
        src137 <= 12'h5ea;
        src138 <= 12'ha9a;
        src139 <= 12'hfd0;
        src140 <= 12'hc02;
        src141 <= 12'h66c;
        src142 <= 12'hfdb;
        src143 <= 12'h62;
        src144 <= 12'h7;
        src145 <= 12'h472;
        src146 <= 12'h99f;
        src147 <= 12'h107;
        src148 <= 12'hb3d;
        src149 <= 12'hca;
        src150 <= 12'h576;
        src151 <= 12'hf4a;
        src152 <= 12'h968;
        src153 <= 12'h7f7;
        src154 <= 12'he93;
        src155 <= 12'he48;
        src156 <= 12'hafe;
        src157 <= 12'hd72;
        src158 <= 12'h57f;
        src159 <= 12'heba;
        src160 <= 12'h62f;
        src161 <= 12'hb79;
        src162 <= 12'h402;
        src163 <= 12'h57a;
        src164 <= 12'h638;
        src165 <= 12'h7a0;
        src166 <= 12'h78f;
        src167 <= 12'haf9;
        src168 <= 12'he6;
        src169 <= 12'he7f;
        src170 <= 12'h140;
        src171 <= 12'h82d;
        src172 <= 12'h5eb;
        src173 <= 12'hc5c;
        src174 <= 12'hc1c;
        src175 <= 12'h94d;
        src176 <= 12'h432;
        src177 <= 12'h27d;
        src178 <= 12'ha78;
        src179 <= 12'hd11;
        src180 <= 12'hf2f;
        src181 <= 12'hd;
        src182 <= 12'h87c;
        src183 <= 12'hc3c;
        src184 <= 12'h27b;
        src185 <= 12'hff7;
        src186 <= 12'h430;
        src187 <= 12'h4ec;
        src188 <= 12'hf34;
        exp <= 20'h6370d;
        #1
        src0 <= 12'hae4;
        src1 <= 12'hdc6;
        src2 <= 12'hb0d;
        src3 <= 12'h9c6;
        src4 <= 12'h84f;
        src5 <= 12'h379;
        src6 <= 12'h91c;
        src7 <= 12'h843;
        src8 <= 12'h7ef;
        src9 <= 12'h894;
        src10 <= 12'ha98;
        src11 <= 12'hfdc;
        src12 <= 12'h2b9;
        src13 <= 12'h259;
        src14 <= 12'h37e;
        src15 <= 12'h68f;
        src16 <= 12'h4f3;
        src17 <= 12'h91c;
        src18 <= 12'hbf;
        src19 <= 12'h4a4;
        src20 <= 12'h3c3;
        src21 <= 12'h729;
        src22 <= 12'hda4;
        src23 <= 12'h4b1;
        src24 <= 12'he58;
        src25 <= 12'hff7;
        src26 <= 12'hc;
        src27 <= 12'h379;
        src28 <= 12'hdc2;
        src29 <= 12'h20a;
        src30 <= 12'hf17;
        src31 <= 12'h34e;
        src32 <= 12'h47e;
        src33 <= 12'h4e9;
        src34 <= 12'h22;
        src35 <= 12'hf32;
        src36 <= 12'hb3e;
        src37 <= 12'h34f;
        src38 <= 12'h3d7;
        src39 <= 12'h781;
        src40 <= 12'h87f;
        src41 <= 12'h4d8;
        src42 <= 12'hb90;
        src43 <= 12'h372;
        src44 <= 12'hdc2;
        src45 <= 12'hd0a;
        src46 <= 12'h6b6;
        src47 <= 12'h4e1;
        src48 <= 12'h176;
        src49 <= 12'hd8e;
        src50 <= 12'h298;
        src51 <= 12'h54b;
        src52 <= 12'haf2;
        src53 <= 12'h52d;
        src54 <= 12'h548;
        src55 <= 12'h36d;
        src56 <= 12'hec6;
        src57 <= 12'h8e;
        src58 <= 12'hb67;
        src59 <= 12'haf2;
        src60 <= 12'hfbc;
        src61 <= 12'h56c;
        src62 <= 12'hf3f;
        src63 <= 12'h29b;
        src64 <= 12'h701;
        src65 <= 12'h1d2;
        src66 <= 12'h47f;
        src67 <= 12'h4ed;
        src68 <= 12'hac3;
        src69 <= 12'he97;
        src70 <= 12'h95b;
        src71 <= 12'h10f;
        src72 <= 12'hacb;
        src73 <= 12'hed9;
        src74 <= 12'h6c8;
        src75 <= 12'hb4d;
        src76 <= 12'h4a3;
        src77 <= 12'hdf0;
        src78 <= 12'h176;
        src79 <= 12'h606;
        src80 <= 12'h74f;
        src81 <= 12'h7c5;
        src82 <= 12'hc1f;
        src83 <= 12'ha0e;
        src84 <= 12'h14f;
        src85 <= 12'h72a;
        src86 <= 12'h7f9;
        src87 <= 12'h7d4;
        src88 <= 12'h9cd;
        src89 <= 12'h3e;
        src90 <= 12'hbde;
        src91 <= 12'he2a;
        src92 <= 12'hbf7;
        src93 <= 12'h226;
        src94 <= 12'h9c7;
        src95 <= 12'hfb7;
        src96 <= 12'hd9b;
        src97 <= 12'h46f;
        src98 <= 12'h24b;
        src99 <= 12'h205;
        src100 <= 12'he2e;
        src101 <= 12'h890;
        src102 <= 12'h244;
        src103 <= 12'he51;
        src104 <= 12'h5cc;
        src105 <= 12'h2dc;
        src106 <= 12'h523;
        src107 <= 12'hda;
        src108 <= 12'ha1e;
        src109 <= 12'h74a;
        src110 <= 12'hd1b;
        src111 <= 12'h6ed;
        src112 <= 12'h87f;
        src113 <= 12'hbd4;
        src114 <= 12'h3df;
        src115 <= 12'h43e;
        src116 <= 12'hf61;
        src117 <= 12'he8;
        src118 <= 12'ha5e;
        src119 <= 12'h2e9;
        src120 <= 12'h59a;
        src121 <= 12'h6c0;
        src122 <= 12'h274;
        src123 <= 12'he47;
        src124 <= 12'h33b;
        src125 <= 12'h67;
        src126 <= 12'h7e4;
        src127 <= 12'haac;
        src128 <= 12'h279;
        src129 <= 12'hc29;
        src130 <= 12'hba7;
        src131 <= 12'h3b9;
        src132 <= 12'hccb;
        src133 <= 12'ha5b;
        src134 <= 12'h39b;
        src135 <= 12'h6dc;
        src136 <= 12'hae7;
        src137 <= 12'h4bb;
        src138 <= 12'hcd4;
        src139 <= 12'h94;
        src140 <= 12'h41a;
        src141 <= 12'h7d8;
        src142 <= 12'ha6d;
        src143 <= 12'h6c6;
        src144 <= 12'h8a4;
        src145 <= 12'h86d;
        src146 <= 12'hbb1;
        src147 <= 12'ha04;
        src148 <= 12'ha8f;
        src149 <= 12'hb56;
        src150 <= 12'h445;
        src151 <= 12'hb36;
        src152 <= 12'hfd4;
        src153 <= 12'h448;
        src154 <= 12'h34f;
        src155 <= 12'h242;
        src156 <= 12'h663;
        src157 <= 12'h86c;
        src158 <= 12'h87;
        src159 <= 12'h584;
        src160 <= 12'hc7f;
        src161 <= 12'h14c;
        src162 <= 12'h381;
        src163 <= 12'h688;
        src164 <= 12'h1f4;
        src165 <= 12'h95b;
        src166 <= 12'hbe5;
        src167 <= 12'h6b7;
        src168 <= 12'hd6f;
        src169 <= 12'h14;
        src170 <= 12'h673;
        src171 <= 12'he9d;
        src172 <= 12'h94c;
        src173 <= 12'h80c;
        src174 <= 12'h49e;
        src175 <= 12'h7f5;
        src176 <= 12'he84;
        src177 <= 12'hdd7;
        src178 <= 12'hc81;
        src179 <= 12'h42a;
        src180 <= 12'hc92;
        src181 <= 12'h679;
        src182 <= 12'h33;
        src183 <= 12'h653;
        src184 <= 12'h1dc;
        src185 <= 12'h1e3;
        src186 <= 12'h189;
        src187 <= 12'h123;
        src188 <= 12'h538;
        exp <= 20'h58c33;
        #1
        src0 <= 12'h6ea;
        src1 <= 12'h8a9;
        src2 <= 12'h96a;
        src3 <= 12'h162;
        src4 <= 12'h91b;
        src5 <= 12'hb9e;
        src6 <= 12'h499;
        src7 <= 12'had3;
        src8 <= 12'hf19;
        src9 <= 12'hecc;
        src10 <= 12'h472;
        src11 <= 12'h587;
        src12 <= 12'h4bb;
        src13 <= 12'h4f9;
        src14 <= 12'h87c;
        src15 <= 12'h96b;
        src16 <= 12'h443;
        src17 <= 12'h395;
        src18 <= 12'h5de;
        src19 <= 12'h1ed;
        src20 <= 12'hf37;
        src21 <= 12'h56;
        src22 <= 12'hdd0;
        src23 <= 12'h9ab;
        src24 <= 12'hd9c;
        src25 <= 12'hd12;
        src26 <= 12'h70;
        src27 <= 12'h187;
        src28 <= 12'hafa;
        src29 <= 12'hb4;
        src30 <= 12'hb61;
        src31 <= 12'h3bc;
        src32 <= 12'h653;
        src33 <= 12'h7e;
        src34 <= 12'he3a;
        src35 <= 12'ha7a;
        src36 <= 12'h1f6;
        src37 <= 12'hbee;
        src38 <= 12'h917;
        src39 <= 12'h514;
        src40 <= 12'h79b;
        src41 <= 12'h256;
        src42 <= 12'ha6e;
        src43 <= 12'h851;
        src44 <= 12'h4d1;
        src45 <= 12'h292;
        src46 <= 12'hba6;
        src47 <= 12'h91c;
        src48 <= 12'he4d;
        src49 <= 12'hdb0;
        src50 <= 12'hfe0;
        src51 <= 12'h656;
        src52 <= 12'ha5b;
        src53 <= 12'hb69;
        src54 <= 12'h12e;
        src55 <= 12'h3ff;
        src56 <= 12'h997;
        src57 <= 12'h982;
        src58 <= 12'h17a;
        src59 <= 12'h8ff;
        src60 <= 12'h553;
        src61 <= 12'h628;
        src62 <= 12'hcd5;
        src63 <= 12'h65d;
        src64 <= 12'h4ae;
        src65 <= 12'h3a3;
        src66 <= 12'he22;
        src67 <= 12'h170;
        src68 <= 12'hafc;
        src69 <= 12'h859;
        src70 <= 12'h2de;
        src71 <= 12'h790;
        src72 <= 12'h680;
        src73 <= 12'h126;
        src74 <= 12'h5ba;
        src75 <= 12'he67;
        src76 <= 12'h159;
        src77 <= 12'h7c7;
        src78 <= 12'h67;
        src79 <= 12'he45;
        src80 <= 12'h276;
        src81 <= 12'h4ea;
        src82 <= 12'h4b7;
        src83 <= 12'he2;
        src84 <= 12'h765;
        src85 <= 12'ha4d;
        src86 <= 12'h566;
        src87 <= 12'hd57;
        src88 <= 12'h96f;
        src89 <= 12'hd2f;
        src90 <= 12'h1b2;
        src91 <= 12'he7e;
        src92 <= 12'h5dd;
        src93 <= 12'h773;
        src94 <= 12'hd13;
        src95 <= 12'h5cc;
        src96 <= 12'h5b4;
        src97 <= 12'hd91;
        src98 <= 12'h267;
        src99 <= 12'hd55;
        src100 <= 12'h985;
        src101 <= 12'hd53;
        src102 <= 12'hd0b;
        src103 <= 12'h84a;
        src104 <= 12'h0;
        src105 <= 12'h9bc;
        src106 <= 12'hfcc;
        src107 <= 12'h395;
        src108 <= 12'hba6;
        src109 <= 12'h78;
        src110 <= 12'h892;
        src111 <= 12'h77b;
        src112 <= 12'h964;
        src113 <= 12'h126;
        src114 <= 12'h451;
        src115 <= 12'h77a;
        src116 <= 12'h5b6;
        src117 <= 12'h6e2;
        src118 <= 12'h4be;
        src119 <= 12'h786;
        src120 <= 12'he00;
        src121 <= 12'h48e;
        src122 <= 12'h805;
        src123 <= 12'h64a;
        src124 <= 12'hba9;
        src125 <= 12'h7e0;
        src126 <= 12'h49a;
        src127 <= 12'he20;
        src128 <= 12'h433;
        src129 <= 12'he7;
        src130 <= 12'hd35;
        src131 <= 12'h28b;
        src132 <= 12'h69f;
        src133 <= 12'h1be;
        src134 <= 12'h9c6;
        src135 <= 12'h7eb;
        src136 <= 12'ha2d;
        src137 <= 12'h184;
        src138 <= 12'h569;
        src139 <= 12'h43f;
        src140 <= 12'hbe0;
        src141 <= 12'ha4;
        src142 <= 12'hb40;
        src143 <= 12'hf7b;
        src144 <= 12'h8ff;
        src145 <= 12'h611;
        src146 <= 12'h16e;
        src147 <= 12'h291;
        src148 <= 12'hdbc;
        src149 <= 12'h6df;
        src150 <= 12'h79b;
        src151 <= 12'h12d;
        src152 <= 12'ha0b;
        src153 <= 12'h3b4;
        src154 <= 12'hcd1;
        src155 <= 12'hc7c;
        src156 <= 12'h7a7;
        src157 <= 12'h9ab;
        src158 <= 12'hf1;
        src159 <= 12'hd87;
        src160 <= 12'h135;
        src161 <= 12'hbf1;
        src162 <= 12'h371;
        src163 <= 12'h53e;
        src164 <= 12'h53f;
        src165 <= 12'h9db;
        src166 <= 12'hed5;
        src167 <= 12'h65f;
        src168 <= 12'h42c;
        src169 <= 12'h1dc;
        src170 <= 12'hd9c;
        src171 <= 12'h317;
        src172 <= 12'hb55;
        src173 <= 12'h7b3;
        src174 <= 12'h23d;
        src175 <= 12'h620;
        src176 <= 12'h71c;
        src177 <= 12'h888;
        src178 <= 12'hef3;
        src179 <= 12'hbb;
        src180 <= 12'hc58;
        src181 <= 12'h627;
        src182 <= 12'h20d;
        src183 <= 12'h8ca;
        src184 <= 12'hf0b;
        src185 <= 12'hf7c;
        src186 <= 12'ha6a;
        src187 <= 12'h209;
        src188 <= 12'hf43;
        exp <= 20'h59439;
        #1
        src0 <= 12'h7a0;
        src1 <= 12'h95a;
        src2 <= 12'hfac;
        src3 <= 12'h397;
        src4 <= 12'h469;
        src5 <= 12'h2e2;
        src6 <= 12'h859;
        src7 <= 12'h401;
        src8 <= 12'h15e;
        src9 <= 12'h254;
        src10 <= 12'h217;
        src11 <= 12'h979;
        src12 <= 12'ha1a;
        src13 <= 12'hf11;
        src14 <= 12'h131;
        src15 <= 12'hf89;
        src16 <= 12'h396;
        src17 <= 12'hd40;
        src18 <= 12'he16;
        src19 <= 12'had3;
        src20 <= 12'hfc2;
        src21 <= 12'he69;
        src22 <= 12'hc4b;
        src23 <= 12'hb1e;
        src24 <= 12'h2c3;
        src25 <= 12'h1ad;
        src26 <= 12'h96d;
        src27 <= 12'hc87;
        src28 <= 12'h455;
        src29 <= 12'hc21;
        src30 <= 12'haa;
        src31 <= 12'h9a3;
        src32 <= 12'h87a;
        src33 <= 12'hdab;
        src34 <= 12'he29;
        src35 <= 12'h97b;
        src36 <= 12'h4b0;
        src37 <= 12'h9e9;
        src38 <= 12'hc58;
        src39 <= 12'h1e7;
        src40 <= 12'h6e6;
        src41 <= 12'h4a9;
        src42 <= 12'hfd3;
        src43 <= 12'h109;
        src44 <= 12'hb38;
        src45 <= 12'h60d;
        src46 <= 12'h2eb;
        src47 <= 12'h7e1;
        src48 <= 12'hffb;
        src49 <= 12'h3e4;
        src50 <= 12'h8d5;
        src51 <= 12'h589;
        src52 <= 12'he64;
        src53 <= 12'h61b;
        src54 <= 12'hf14;
        src55 <= 12'h641;
        src56 <= 12'hbbc;
        src57 <= 12'hb73;
        src58 <= 12'h9a4;
        src59 <= 12'haf5;
        src60 <= 12'h903;
        src61 <= 12'hb43;
        src62 <= 12'h1e9;
        src63 <= 12'h74e;
        src64 <= 12'h841;
        src65 <= 12'h8a8;
        src66 <= 12'h991;
        src67 <= 12'h810;
        src68 <= 12'h382;
        src69 <= 12'h102;
        src70 <= 12'h8ae;
        src71 <= 12'h565;
        src72 <= 12'h7c5;
        src73 <= 12'h3cf;
        src74 <= 12'h5c1;
        src75 <= 12'hbc4;
        src76 <= 12'h7f5;
        src77 <= 12'h9de;
        src78 <= 12'h6f6;
        src79 <= 12'h77b;
        src80 <= 12'hf32;
        src81 <= 12'h828;
        src82 <= 12'h3bf;
        src83 <= 12'h358;
        src84 <= 12'hc0e;
        src85 <= 12'h81e;
        src86 <= 12'h361;
        src87 <= 12'h659;
        src88 <= 12'ha73;
        src89 <= 12'h1f8;
        src90 <= 12'h62f;
        src91 <= 12'h352;
        src92 <= 12'h373;
        src93 <= 12'ha07;
        src94 <= 12'h431;
        src95 <= 12'h155;
        src96 <= 12'hf6f;
        src97 <= 12'h368;
        src98 <= 12'hca0;
        src99 <= 12'h5cb;
        src100 <= 12'hefa;
        src101 <= 12'h711;
        src102 <= 12'h4ed;
        src103 <= 12'h624;
        src104 <= 12'h4e1;
        src105 <= 12'hc01;
        src106 <= 12'h9f7;
        src107 <= 12'ha13;
        src108 <= 12'h7cc;
        src109 <= 12'hab5;
        src110 <= 12'ha51;
        src111 <= 12'hfad;
        src112 <= 12'h31c;
        src113 <= 12'h55a;
        src114 <= 12'h87c;
        src115 <= 12'hbfc;
        src116 <= 12'h8d0;
        src117 <= 12'hd31;
        src118 <= 12'h349;
        src119 <= 12'h418;
        src120 <= 12'h213;
        src121 <= 12'h903;
        src122 <= 12'h282;
        src123 <= 12'h954;
        src124 <= 12'h57a;
        src125 <= 12'h9f0;
        src126 <= 12'h71e;
        src127 <= 12'h831;
        src128 <= 12'h5c2;
        src129 <= 12'hf19;
        src130 <= 12'h912;
        src131 <= 12'haae;
        src132 <= 12'h726;
        src133 <= 12'h66b;
        src134 <= 12'h2f3;
        src135 <= 12'h761;
        src136 <= 12'h2c3;
        src137 <= 12'hb52;
        src138 <= 12'hd00;
        src139 <= 12'hcbf;
        src140 <= 12'ha81;
        src141 <= 12'hd15;
        src142 <= 12'haf6;
        src143 <= 12'h72a;
        src144 <= 12'h19a;
        src145 <= 12'h839;
        src146 <= 12'h93d;
        src147 <= 12'h1a0;
        src148 <= 12'h1d;
        src149 <= 12'h3aa;
        src150 <= 12'h62f;
        src151 <= 12'h88a;
        src152 <= 12'hb82;
        src153 <= 12'h703;
        src154 <= 12'h86c;
        src155 <= 12'h9c0;
        src156 <= 12'hced;
        src157 <= 12'h2dc;
        src158 <= 12'h9d9;
        src159 <= 12'he19;
        src160 <= 12'hd0a;
        src161 <= 12'hacb;
        src162 <= 12'h310;
        src163 <= 12'h407;
        src164 <= 12'h73f;
        src165 <= 12'h2f9;
        src166 <= 12'hdf7;
        src167 <= 12'heb9;
        src168 <= 12'hfea;
        src169 <= 12'ha97;
        src170 <= 12'h9ad;
        src171 <= 12'hd93;
        src172 <= 12'h56b;
        src173 <= 12'hf1d;
        src174 <= 12'h728;
        src175 <= 12'h324;
        src176 <= 12'h4c3;
        src177 <= 12'hd75;
        src178 <= 12'h3ee;
        src179 <= 12'hdc7;
        src180 <= 12'hccf;
        src181 <= 12'h2fb;
        src182 <= 12'h761;
        src183 <= 12'h54d;
        src184 <= 12'h473;
        src185 <= 12'h5df;
        src186 <= 12'hec8;
        src187 <= 12'hc4d;
        src188 <= 12'h2d2;
        exp <= 20'h60222;
        #1
        src0 <= 12'h1f9;
        src1 <= 12'hfe8;
        src2 <= 12'h314;
        src3 <= 12'hf2e;
        src4 <= 12'h558;
        src5 <= 12'h9f2;
        src6 <= 12'h6e9;
        src7 <= 12'h4e5;
        src8 <= 12'h793;
        src9 <= 12'ha9;
        src10 <= 12'hc4;
        src11 <= 12'he26;
        src12 <= 12'h749;
        src13 <= 12'he7f;
        src14 <= 12'h1d9;
        src15 <= 12'h146;
        src16 <= 12'hf3d;
        src17 <= 12'h26;
        src18 <= 12'h9eb;
        src19 <= 12'hb70;
        src20 <= 12'h5f9;
        src21 <= 12'hec4;
        src22 <= 12'h2ef;
        src23 <= 12'h992;
        src24 <= 12'h5b;
        src25 <= 12'hbc4;
        src26 <= 12'hc16;
        src27 <= 12'h3ce;
        src28 <= 12'hf84;
        src29 <= 12'hb3f;
        src30 <= 12'h1e1;
        src31 <= 12'h670;
        src32 <= 12'h219;
        src33 <= 12'he03;
        src34 <= 12'h20c;
        src35 <= 12'h298;
        src36 <= 12'h6cd;
        src37 <= 12'hb7d;
        src38 <= 12'h9b4;
        src39 <= 12'h56;
        src40 <= 12'h33f;
        src41 <= 12'he58;
        src42 <= 12'he17;
        src43 <= 12'hb42;
        src44 <= 12'h968;
        src45 <= 12'h296;
        src46 <= 12'hd7c;
        src47 <= 12'h354;
        src48 <= 12'h8cd;
        src49 <= 12'h69f;
        src50 <= 12'he2d;
        src51 <= 12'hddc;
        src52 <= 12'h749;
        src53 <= 12'h432;
        src54 <= 12'h8b9;
        src55 <= 12'hbf7;
        src56 <= 12'he9c;
        src57 <= 12'h935;
        src58 <= 12'hf75;
        src59 <= 12'hf55;
        src60 <= 12'h776;
        src61 <= 12'h669;
        src62 <= 12'h5ae;
        src63 <= 12'hb5a;
        src64 <= 12'ha7a;
        src65 <= 12'h163;
        src66 <= 12'h5a0;
        src67 <= 12'h7a7;
        src68 <= 12'h597;
        src69 <= 12'h3ef;
        src70 <= 12'hd8d;
        src71 <= 12'hb4f;
        src72 <= 12'h9fe;
        src73 <= 12'h93d;
        src74 <= 12'he1a;
        src75 <= 12'hb1b;
        src76 <= 12'h9af;
        src77 <= 12'hcbb;
        src78 <= 12'hc4;
        src79 <= 12'hae3;
        src80 <= 12'h16c;
        src81 <= 12'h4ff;
        src82 <= 12'h3f1;
        src83 <= 12'ha06;
        src84 <= 12'hade;
        src85 <= 12'h295;
        src86 <= 12'hbb9;
        src87 <= 12'h6e9;
        src88 <= 12'h83f;
        src89 <= 12'h656;
        src90 <= 12'h20e;
        src91 <= 12'h137;
        src92 <= 12'h14a;
        src93 <= 12'h44;
        src94 <= 12'h22e;
        src95 <= 12'h200;
        src96 <= 12'h9e9;
        src97 <= 12'hf79;
        src98 <= 12'he14;
        src99 <= 12'hbd6;
        src100 <= 12'hd9c;
        src101 <= 12'hb70;
        src102 <= 12'h6d3;
        src103 <= 12'h1b0;
        src104 <= 12'hd0c;
        src105 <= 12'hdec;
        src106 <= 12'hdb9;
        src107 <= 12'hb08;
        src108 <= 12'h63;
        src109 <= 12'h54b;
        src110 <= 12'hc1;
        src111 <= 12'hafe;
        src112 <= 12'heed;
        src113 <= 12'h672;
        src114 <= 12'hc52;
        src115 <= 12'h1a4;
        src116 <= 12'h678;
        src117 <= 12'haac;
        src118 <= 12'h52c;
        src119 <= 12'h527;
        src120 <= 12'h7af;
        src121 <= 12'h41d;
        src122 <= 12'h113;
        src123 <= 12'hac1;
        src124 <= 12'hfe3;
        src125 <= 12'hbfb;
        src126 <= 12'h227;
        src127 <= 12'h8d7;
        src128 <= 12'ha67;
        src129 <= 12'haa8;
        src130 <= 12'ha10;
        src131 <= 12'hebd;
        src132 <= 12'h5bd;
        src133 <= 12'h914;
        src134 <= 12'h70e;
        src135 <= 12'hd4b;
        src136 <= 12'h8de;
        src137 <= 12'hdd8;
        src138 <= 12'h93;
        src139 <= 12'ha2c;
        src140 <= 12'h8ff;
        src141 <= 12'hbbf;
        src142 <= 12'h1e3;
        src143 <= 12'hd06;
        src144 <= 12'h52c;
        src145 <= 12'h292;
        src146 <= 12'hd8;
        src147 <= 12'he51;
        src148 <= 12'h53e;
        src149 <= 12'h475;
        src150 <= 12'hbbb;
        src151 <= 12'h60d;
        src152 <= 12'h3d6;
        src153 <= 12'h94b;
        src154 <= 12'h11;
        src155 <= 12'h617;
        src156 <= 12'hbac;
        src157 <= 12'h700;
        src158 <= 12'hee9;
        src159 <= 12'h63c;
        src160 <= 12'hf8e;
        src161 <= 12'hfdf;
        src162 <= 12'h896;
        src163 <= 12'ha91;
        src164 <= 12'hb7f;
        src165 <= 12'h491;
        src166 <= 12'h1a5;
        src167 <= 12'hb82;
        src168 <= 12'hbab;
        src169 <= 12'h274;
        src170 <= 12'ha4d;
        src171 <= 12'h716;
        src172 <= 12'h3d5;
        src173 <= 12'h5f5;
        src174 <= 12'h16c;
        src175 <= 12'hb3c;
        src176 <= 12'h1dc;
        src177 <= 12'h94b;
        src178 <= 12'h442;
        src179 <= 12'h5d9;
        src180 <= 12'hfd2;
        src181 <= 12'h79e;
        src182 <= 12'h58f;
        src183 <= 12'hd89;
        src184 <= 12'h59b;
        src185 <= 12'hdf8;
        src186 <= 12'he76;
        src187 <= 12'h4a0;
        src188 <= 12'hc01;
        exp <= 20'h5f77d;
        #1
        src0 <= 12'hd8d;
        src1 <= 12'hb71;
        src2 <= 12'h71b;
        src3 <= 12'ha03;
        src4 <= 12'hba4;
        src5 <= 12'h6d4;
        src6 <= 12'h16d;
        src7 <= 12'h8b6;
        src8 <= 12'hea;
        src9 <= 12'hedf;
        src10 <= 12'h238;
        src11 <= 12'h781;
        src12 <= 12'h883;
        src13 <= 12'h1a8;
        src14 <= 12'h4b8;
        src15 <= 12'h5d;
        src16 <= 12'h806;
        src17 <= 12'h2fb;
        src18 <= 12'h6e;
        src19 <= 12'h572;
        src20 <= 12'h919;
        src21 <= 12'h7c5;
        src22 <= 12'he36;
        src23 <= 12'h8b6;
        src24 <= 12'h46b;
        src25 <= 12'h596;
        src26 <= 12'h8d0;
        src27 <= 12'hc16;
        src28 <= 12'h3ba;
        src29 <= 12'haa7;
        src30 <= 12'h7bd;
        src31 <= 12'h28;
        src32 <= 12'h1c2;
        src33 <= 12'h1ad;
        src34 <= 12'hd0;
        src35 <= 12'h82c;
        src36 <= 12'h985;
        src37 <= 12'h16c;
        src38 <= 12'he3f;
        src39 <= 12'hb8a;
        src40 <= 12'h1f;
        src41 <= 12'hc82;
        src42 <= 12'hbe6;
        src43 <= 12'h2f7;
        src44 <= 12'h945;
        src45 <= 12'hca3;
        src46 <= 12'hb18;
        src47 <= 12'h3b1;
        src48 <= 12'hef2;
        src49 <= 12'h8d5;
        src50 <= 12'h8f6;
        src51 <= 12'hf7;
        src52 <= 12'hc42;
        src53 <= 12'h86;
        src54 <= 12'h3f1;
        src55 <= 12'h469;
        src56 <= 12'hc70;
        src57 <= 12'ha83;
        src58 <= 12'hb39;
        src59 <= 12'h915;
        src60 <= 12'hba4;
        src61 <= 12'h688;
        src62 <= 12'hff4;
        src63 <= 12'hded;
        src64 <= 12'h8cc;
        src65 <= 12'hb7;
        src66 <= 12'h7b8;
        src67 <= 12'hd43;
        src68 <= 12'h76e;
        src69 <= 12'h46e;
        src70 <= 12'haf7;
        src71 <= 12'he42;
        src72 <= 12'hacf;
        src73 <= 12'hcd7;
        src74 <= 12'h1b7;
        src75 <= 12'hd9a;
        src76 <= 12'ha9f;
        src77 <= 12'h7b4;
        src78 <= 12'h435;
        src79 <= 12'hadb;
        src80 <= 12'hf1f;
        src81 <= 12'h198;
        src82 <= 12'hc2;
        src83 <= 12'hf1f;
        src84 <= 12'h2a1;
        src85 <= 12'hbef;
        src86 <= 12'hd9a;
        src87 <= 12'h8c2;
        src88 <= 12'h8af;
        src89 <= 12'h46c;
        src90 <= 12'h234;
        src91 <= 12'hf36;
        src92 <= 12'h7d0;
        src93 <= 12'h591;
        src94 <= 12'hd32;
        src95 <= 12'hafb;
        src96 <= 12'h4b9;
        src97 <= 12'hf0;
        src98 <= 12'h3f6;
        src99 <= 12'hd91;
        src100 <= 12'hccb;
        src101 <= 12'h906;
        src102 <= 12'h170;
        src103 <= 12'hf3;
        src104 <= 12'haf8;
        src105 <= 12'h304;
        src106 <= 12'h1bd;
        src107 <= 12'h753;
        src108 <= 12'h459;
        src109 <= 12'hc96;
        src110 <= 12'ha74;
        src111 <= 12'h8dd;
        src112 <= 12'h13b;
        src113 <= 12'h846;
        src114 <= 12'hdb2;
        src115 <= 12'h7ee;
        src116 <= 12'h539;
        src117 <= 12'hbbe;
        src118 <= 12'h673;
        src119 <= 12'hc48;
        src120 <= 12'hf0a;
        src121 <= 12'h35e;
        src122 <= 12'h301;
        src123 <= 12'h96a;
        src124 <= 12'h9e1;
        src125 <= 12'h3ba;
        src126 <= 12'h201;
        src127 <= 12'h7b0;
        src128 <= 12'ha58;
        src129 <= 12'ha;
        src130 <= 12'h8e0;
        src131 <= 12'hda3;
        src132 <= 12'h732;
        src133 <= 12'h2a4;
        src134 <= 12'h6;
        src135 <= 12'h2a4;
        src136 <= 12'h3;
        src137 <= 12'h3c1;
        src138 <= 12'h9d6;
        src139 <= 12'h62e;
        src140 <= 12'h2ef;
        src141 <= 12'h9fb;
        src142 <= 12'h2a3;
        src143 <= 12'h5a1;
        src144 <= 12'h83f;
        src145 <= 12'h2ec;
        src146 <= 12'hd5c;
        src147 <= 12'h1c;
        src148 <= 12'h286;
        src149 <= 12'hc96;
        src150 <= 12'hc60;
        src151 <= 12'ha92;
        src152 <= 12'h4ba;
        src153 <= 12'h304;
        src154 <= 12'h573;
        src155 <= 12'h258;
        src156 <= 12'hf73;
        src157 <= 12'h776;
        src158 <= 12'h828;
        src159 <= 12'hc4e;
        src160 <= 12'h8ba;
        src161 <= 12'hb52;
        src162 <= 12'h4ec;
        src163 <= 12'h223;
        src164 <= 12'h5bc;
        src165 <= 12'h41f;
        src166 <= 12'he76;
        src167 <= 12'h9f6;
        src168 <= 12'h881;
        src169 <= 12'h2d2;
        src170 <= 12'h4d9;
        src171 <= 12'hb88;
        src172 <= 12'hfea;
        src173 <= 12'hdfd;
        src174 <= 12'he29;
        src175 <= 12'ha0a;
        src176 <= 12'h8fb;
        src177 <= 12'hfb7;
        src178 <= 12'hc2;
        src179 <= 12'h479;
        src180 <= 12'he52;
        src181 <= 12'h7ec;
        src182 <= 12'h211;
        src183 <= 12'h148;
        src184 <= 12'h3bd;
        src185 <= 12'h4b6;
        src186 <= 12'h899;
        src187 <= 12'h76f;
        src188 <= 12'hf18;
        exp <= 20'h5982a;
        #1
        src0 <= 12'hc69;
        src1 <= 12'h9e2;
        src2 <= 12'hd8d;
        src3 <= 12'he5d;
        src4 <= 12'h9dc;
        src5 <= 12'h85e;
        src6 <= 12'h60c;
        src7 <= 12'h1b3;
        src8 <= 12'h605;
        src9 <= 12'hc6d;
        src10 <= 12'hb62;
        src11 <= 12'h620;
        src12 <= 12'h8ec;
        src13 <= 12'h37;
        src14 <= 12'h6e7;
        src15 <= 12'hdab;
        src16 <= 12'h954;
        src17 <= 12'h3db;
        src18 <= 12'h535;
        src19 <= 12'h163;
        src20 <= 12'h909;
        src21 <= 12'h88a;
        src22 <= 12'hab8;
        src23 <= 12'h30e;
        src24 <= 12'h5b0;
        src25 <= 12'hd57;
        src26 <= 12'hf6d;
        src27 <= 12'hf9;
        src28 <= 12'hcf0;
        src29 <= 12'hc47;
        src30 <= 12'h644;
        src31 <= 12'h981;
        src32 <= 12'hdd7;
        src33 <= 12'h5e7;
        src34 <= 12'hbd8;
        src35 <= 12'h73;
        src36 <= 12'h601;
        src37 <= 12'h697;
        src38 <= 12'hf17;
        src39 <= 12'h66e;
        src40 <= 12'h3aa;
        src41 <= 12'h4b4;
        src42 <= 12'heb3;
        src43 <= 12'hd4e;
        src44 <= 12'hb13;
        src45 <= 12'hc6d;
        src46 <= 12'h322;
        src47 <= 12'h671;
        src48 <= 12'h5a9;
        src49 <= 12'hfee;
        src50 <= 12'h6f9;
        src51 <= 12'hb3c;
        src52 <= 12'hbff;
        src53 <= 12'h5b9;
        src54 <= 12'h245;
        src55 <= 12'hd0b;
        src56 <= 12'ha47;
        src57 <= 12'h5fb;
        src58 <= 12'h605;
        src59 <= 12'hf8;
        src60 <= 12'h95b;
        src61 <= 12'h2c7;
        src62 <= 12'hfcd;
        src63 <= 12'h224;
        src64 <= 12'hc3e;
        src65 <= 12'h40b;
        src66 <= 12'hc2c;
        src67 <= 12'hf11;
        src68 <= 12'hee2;
        src69 <= 12'h71b;
        src70 <= 12'hb0f;
        src71 <= 12'h812;
        src72 <= 12'h191;
        src73 <= 12'hd91;
        src74 <= 12'h8de;
        src75 <= 12'h7b;
        src76 <= 12'h382;
        src77 <= 12'hb0;
        src78 <= 12'h96;
        src79 <= 12'h407;
        src80 <= 12'hc1d;
        src81 <= 12'h6da;
        src82 <= 12'h8ac;
        src83 <= 12'h6d7;
        src84 <= 12'h962;
        src85 <= 12'h48b;
        src86 <= 12'hea1;
        src87 <= 12'h1ff;
        src88 <= 12'hec;
        src89 <= 12'he1d;
        src90 <= 12'h82b;
        src91 <= 12'hc64;
        src92 <= 12'hcbb;
        src93 <= 12'h28c;
        src94 <= 12'h795;
        src95 <= 12'hb72;
        src96 <= 12'h242;
        src97 <= 12'h7e6;
        src98 <= 12'h72a;
        src99 <= 12'hade;
        src100 <= 12'h6ce;
        src101 <= 12'h9f4;
        src102 <= 12'ha8f;
        src103 <= 12'h1f9;
        src104 <= 12'h9fe;
        src105 <= 12'h9a8;
        src106 <= 12'h432;
        src107 <= 12'ha39;
        src108 <= 12'ha05;
        src109 <= 12'h5b1;
        src110 <= 12'hf1d;
        src111 <= 12'hbeb;
        src112 <= 12'ha95;
        src113 <= 12'h46f;
        src114 <= 12'h3b6;
        src115 <= 12'hd73;
        src116 <= 12'h1f4;
        src117 <= 12'h587;
        src118 <= 12'h6de;
        src119 <= 12'hf68;
        src120 <= 12'hbe3;
        src121 <= 12'hbeb;
        src122 <= 12'hf60;
        src123 <= 12'hbf6;
        src124 <= 12'hb51;
        src125 <= 12'h1e4;
        src126 <= 12'hac4;
        src127 <= 12'hb7c;
        src128 <= 12'h6d8;
        src129 <= 12'h5f7;
        src130 <= 12'h10f;
        src131 <= 12'h79;
        src132 <= 12'h4c5;
        src133 <= 12'h63f;
        src134 <= 12'h31b;
        src135 <= 12'h878;
        src136 <= 12'hf54;
        src137 <= 12'h459;
        src138 <= 12'h3ac;
        src139 <= 12'h76;
        src140 <= 12'hcfc;
        src141 <= 12'hc72;
        src142 <= 12'h63d;
        src143 <= 12'h67b;
        src144 <= 12'hcf4;
        src145 <= 12'hc2d;
        src146 <= 12'he33;
        src147 <= 12'h7a;
        src148 <= 12'hcf7;
        src149 <= 12'h82f;
        src150 <= 12'h60c;
        src151 <= 12'h2fe;
        src152 <= 12'hc02;
        src153 <= 12'ha21;
        src154 <= 12'h586;
        src155 <= 12'h14f;
        src156 <= 12'hb3d;
        src157 <= 12'hfdf;
        src158 <= 12'hec9;
        src159 <= 12'h56e;
        src160 <= 12'h927;
        src161 <= 12'hb19;
        src162 <= 12'h7b2;
        src163 <= 12'hec8;
        src164 <= 12'h11c;
        src165 <= 12'h59a;
        src166 <= 12'h67d;
        src167 <= 12'h9bc;
        src168 <= 12'heea;
        src169 <= 12'h53d;
        src170 <= 12'hc50;
        src171 <= 12'he93;
        src172 <= 12'h56a;
        src173 <= 12'h732;
        src174 <= 12'h218;
        src175 <= 12'h45e;
        src176 <= 12'h41f;
        src177 <= 12'h1ea;
        src178 <= 12'h72a;
        src179 <= 12'hc77;
        src180 <= 12'h25b;
        src181 <= 12'h961;
        src182 <= 12'h324;
        src183 <= 12'h40;
        src184 <= 12'h54f;
        src185 <= 12'h43f;
        src186 <= 12'hef4;
        src187 <= 12'h80b;
        src188 <= 12'h472;
        exp <= 20'h5f183;
        #1
        src0 <= 12'h2e3;
        src1 <= 12'h837;
        src2 <= 12'hf7c;
        src3 <= 12'hb5f;
        src4 <= 12'hfd9;
        src5 <= 12'h999;
        src6 <= 12'hfb;
        src7 <= 12'h6f7;
        src8 <= 12'h74d;
        src9 <= 12'h8a3;
        src10 <= 12'hc92;
        src11 <= 12'hef4;
        src12 <= 12'h9cb;
        src13 <= 12'h758;
        src14 <= 12'h61b;
        src15 <= 12'hbb2;
        src16 <= 12'h7f2;
        src17 <= 12'h826;
        src18 <= 12'h4e;
        src19 <= 12'h635;
        src20 <= 12'hc83;
        src21 <= 12'h618;
        src22 <= 12'ha5b;
        src23 <= 12'ha51;
        src24 <= 12'h34d;
        src25 <= 12'hdb4;
        src26 <= 12'h5a4;
        src27 <= 12'h837;
        src28 <= 12'h29d;
        src29 <= 12'h263;
        src30 <= 12'heb6;
        src31 <= 12'h1a1;
        src32 <= 12'hd3c;
        src33 <= 12'h666;
        src34 <= 12'hfbe;
        src35 <= 12'hc6a;
        src36 <= 12'hee0;
        src37 <= 12'h767;
        src38 <= 12'h6;
        src39 <= 12'h38e;
        src40 <= 12'h17b;
        src41 <= 12'h1cc;
        src42 <= 12'hafb;
        src43 <= 12'hae2;
        src44 <= 12'hd51;
        src45 <= 12'h43b;
        src46 <= 12'h5c;
        src47 <= 12'h872;
        src48 <= 12'h75a;
        src49 <= 12'h456;
        src50 <= 12'hf86;
        src51 <= 12'hfd4;
        src52 <= 12'hfb3;
        src53 <= 12'hc29;
        src54 <= 12'h184;
        src55 <= 12'he30;
        src56 <= 12'h505;
        src57 <= 12'h29f;
        src58 <= 12'haa8;
        src59 <= 12'hd48;
        src60 <= 12'h2a2;
        src61 <= 12'haa4;
        src62 <= 12'he21;
        src63 <= 12'hf37;
        src64 <= 12'hbda;
        src65 <= 12'h43;
        src66 <= 12'h31a;
        src67 <= 12'h19e;
        src68 <= 12'h81c;
        src69 <= 12'hbce;
        src70 <= 12'h41e;
        src71 <= 12'hb8e;
        src72 <= 12'he05;
        src73 <= 12'hd8c;
        src74 <= 12'h4ff;
        src75 <= 12'h37;
        src76 <= 12'h230;
        src77 <= 12'h49d;
        src78 <= 12'h2a;
        src79 <= 12'hc2a;
        src80 <= 12'h1b2;
        src81 <= 12'hbe1;
        src82 <= 12'h117;
        src83 <= 12'h497;
        src84 <= 12'hfc0;
        src85 <= 12'hffb;
        src86 <= 12'ha18;
        src87 <= 12'h842;
        src88 <= 12'h595;
        src89 <= 12'hd96;
        src90 <= 12'ha65;
        src91 <= 12'h3fb;
        src92 <= 12'h321;
        src93 <= 12'hb15;
        src94 <= 12'h540;
        src95 <= 12'h9d;
        src96 <= 12'h1b7;
        src97 <= 12'h69c;
        src98 <= 12'he58;
        src99 <= 12'h6b5;
        src100 <= 12'hdb7;
        src101 <= 12'h70e;
        src102 <= 12'hf9;
        src103 <= 12'hb1f;
        src104 <= 12'h3d5;
        src105 <= 12'he37;
        src106 <= 12'hb2a;
        src107 <= 12'haf2;
        src108 <= 12'h91a;
        src109 <= 12'h130;
        src110 <= 12'ha7e;
        src111 <= 12'h343;
        src112 <= 12'heb2;
        src113 <= 12'hae2;
        src114 <= 12'he79;
        src115 <= 12'hedb;
        src116 <= 12'haa7;
        src117 <= 12'he9;
        src118 <= 12'h200;
        src119 <= 12'hb01;
        src120 <= 12'h8b4;
        src121 <= 12'he2;
        src122 <= 12'h8d7;
        src123 <= 12'h179;
        src124 <= 12'hb18;
        src125 <= 12'h16b;
        src126 <= 12'hce7;
        src127 <= 12'h41f;
        src128 <= 12'h80b;
        src129 <= 12'h802;
        src130 <= 12'ha0b;
        src131 <= 12'h9b8;
        src132 <= 12'hb49;
        src133 <= 12'h266;
        src134 <= 12'h2b5;
        src135 <= 12'h52c;
        src136 <= 12'h6b8;
        src137 <= 12'h5a;
        src138 <= 12'h99;
        src139 <= 12'h71b;
        src140 <= 12'h1b;
        src141 <= 12'head;
        src142 <= 12'h555;
        src143 <= 12'h85c;
        src144 <= 12'h73a;
        src145 <= 12'ha66;
        src146 <= 12'h7e2;
        src147 <= 12'h8d;
        src148 <= 12'hd9c;
        src149 <= 12'h430;
        src150 <= 12'h490;
        src151 <= 12'ha06;
        src152 <= 12'hd22;
        src153 <= 12'hbcc;
        src154 <= 12'h376;
        src155 <= 12'h3f3;
        src156 <= 12'h54c;
        src157 <= 12'h873;
        src158 <= 12'h371;
        src159 <= 12'h317;
        src160 <= 12'h204;
        src161 <= 12'ha2f;
        src162 <= 12'ha97;
        src163 <= 12'h38c;
        src164 <= 12'h744;
        src165 <= 12'hf2c;
        src166 <= 12'h750;
        src167 <= 12'he5b;
        src168 <= 12'h7a0;
        src169 <= 12'ha48;
        src170 <= 12'h5cb;
        src171 <= 12'hd5;
        src172 <= 12'h528;
        src173 <= 12'h1ce;
        src174 <= 12'h56e;
        src175 <= 12'hda2;
        src176 <= 12'he3f;
        src177 <= 12'h1b1;
        src178 <= 12'hf65;
        src179 <= 12'h1e;
        src180 <= 12'h9db;
        src181 <= 12'h1a2;
        src182 <= 12'h6f9;
        src183 <= 12'h889;
        src184 <= 12'h679;
        src185 <= 12'h244;
        src186 <= 12'hbc3;
        src187 <= 12'h2b3;
        src188 <= 12'h243;
        exp <= 20'h5a8f7;
        #1
        src0 <= 12'he88;
        src1 <= 12'h365;
        src2 <= 12'h15b;
        src3 <= 12'h34f;
        src4 <= 12'h4ea;
        src5 <= 12'hac7;
        src6 <= 12'h3b9;
        src7 <= 12'hfd1;
        src8 <= 12'hdb;
        src9 <= 12'h62f;
        src10 <= 12'hc1a;
        src11 <= 12'h606;
        src12 <= 12'h40e;
        src13 <= 12'hbf6;
        src14 <= 12'h446;
        src15 <= 12'hb40;
        src16 <= 12'hbb0;
        src17 <= 12'hb18;
        src18 <= 12'ha0e;
        src19 <= 12'h16a;
        src20 <= 12'h14e;
        src21 <= 12'hfe5;
        src22 <= 12'h89c;
        src23 <= 12'h495;
        src24 <= 12'h516;
        src25 <= 12'h668;
        src26 <= 12'hdc;
        src27 <= 12'ha9c;
        src28 <= 12'hee7;
        src29 <= 12'hb54;
        src30 <= 12'hc4a;
        src31 <= 12'h640;
        src32 <= 12'h890;
        src33 <= 12'h570;
        src34 <= 12'h6bd;
        src35 <= 12'h46f;
        src36 <= 12'hcc9;
        src37 <= 12'hac1;
        src38 <= 12'h9c5;
        src39 <= 12'hc;
        src40 <= 12'hd46;
        src41 <= 12'h2b;
        src42 <= 12'h679;
        src43 <= 12'hd19;
        src44 <= 12'h68c;
        src45 <= 12'h2d0;
        src46 <= 12'h98e;
        src47 <= 12'h4dc;
        src48 <= 12'he;
        src49 <= 12'h16;
        src50 <= 12'he15;
        src51 <= 12'hf0f;
        src52 <= 12'hfa3;
        src53 <= 12'h81a;
        src54 <= 12'h380;
        src55 <= 12'h868;
        src56 <= 12'hb6b;
        src57 <= 12'h2e8;
        src58 <= 12'h5cb;
        src59 <= 12'h2a9;
        src60 <= 12'h7ba;
        src61 <= 12'h15f;
        src62 <= 12'hbfb;
        src63 <= 12'h9fc;
        src64 <= 12'hee5;
        src65 <= 12'h5ed;
        src66 <= 12'h93e;
        src67 <= 12'hfe5;
        src68 <= 12'h6c2;
        src69 <= 12'h1eb;
        src70 <= 12'h51e;
        src71 <= 12'ha25;
        src72 <= 12'hc31;
        src73 <= 12'hf89;
        src74 <= 12'h157;
        src75 <= 12'h2ea;
        src76 <= 12'h6f9;
        src77 <= 12'hd16;
        src78 <= 12'hdb;
        src79 <= 12'h4a;
        src80 <= 12'hb89;
        src81 <= 12'hc67;
        src82 <= 12'h986;
        src83 <= 12'h6da;
        src84 <= 12'h297;
        src85 <= 12'hc91;
        src86 <= 12'h96e;
        src87 <= 12'hec1;
        src88 <= 12'h9e7;
        src89 <= 12'hc69;
        src90 <= 12'h54;
        src91 <= 12'h7ee;
        src92 <= 12'h89c;
        src93 <= 12'h5fd;
        src94 <= 12'h9bf;
        src95 <= 12'h312;
        src96 <= 12'h3a1;
        src97 <= 12'hc7f;
        src98 <= 12'h1c4;
        src99 <= 12'h77f;
        src100 <= 12'h66c;
        src101 <= 12'hc8f;
        src102 <= 12'he7f;
        src103 <= 12'h108;
        src104 <= 12'h2ce;
        src105 <= 12'h24e;
        src106 <= 12'hfd9;
        src107 <= 12'he1f;
        src108 <= 12'hb47;
        src109 <= 12'h8f9;
        src110 <= 12'h8e1;
        src111 <= 12'h714;
        src112 <= 12'h509;
        src113 <= 12'h180;
        src114 <= 12'h93f;
        src115 <= 12'h345;
        src116 <= 12'ha9d;
        src117 <= 12'ha4c;
        src118 <= 12'h8bd;
        src119 <= 12'he9f;
        src120 <= 12'ha1c;
        src121 <= 12'h852;
        src122 <= 12'h4e3;
        src123 <= 12'haf3;
        src124 <= 12'h686;
        src125 <= 12'ha8f;
        src126 <= 12'h399;
        src127 <= 12'h3ae;
        src128 <= 12'h31f;
        src129 <= 12'hfe9;
        src130 <= 12'hace;
        src131 <= 12'h1ea;
        src132 <= 12'h524;
        src133 <= 12'h670;
        src134 <= 12'h6e0;
        src135 <= 12'h1f8;
        src136 <= 12'h82d;
        src137 <= 12'h325;
        src138 <= 12'h9fc;
        src139 <= 12'ha56;
        src140 <= 12'hdc9;
        src141 <= 12'h739;
        src142 <= 12'h1f1;
        src143 <= 12'hbdc;
        src144 <= 12'hdb9;
        src145 <= 12'hb93;
        src146 <= 12'hf41;
        src147 <= 12'h2c6;
        src148 <= 12'h3fe;
        src149 <= 12'ha06;
        src150 <= 12'h46b;
        src151 <= 12'h22e;
        src152 <= 12'hbda;
        src153 <= 12'h100;
        src154 <= 12'hc30;
        src155 <= 12'h1a2;
        src156 <= 12'h414;
        src157 <= 12'hd16;
        src158 <= 12'h320;
        src159 <= 12'hfb2;
        src160 <= 12'h5a8;
        src161 <= 12'h8b8;
        src162 <= 12'hfe4;
        src163 <= 12'hfb6;
        src164 <= 12'h201;
        src165 <= 12'hbf0;
        src166 <= 12'h468;
        src167 <= 12'he3b;
        src168 <= 12'h304;
        src169 <= 12'he5e;
        src170 <= 12'hf02;
        src171 <= 12'h9e1;
        src172 <= 12'h17e;
        src173 <= 12'h753;
        src174 <= 12'h65b;
        src175 <= 12'h715;
        src176 <= 12'hd46;
        src177 <= 12'h831;
        src178 <= 12'hdfc;
        src179 <= 12'hf2d;
        src180 <= 12'hc3;
        src181 <= 12'h164;
        src182 <= 12'h1a7;
        src183 <= 12'hd48;
        src184 <= 12'hc13;
        src185 <= 12'h700;
        src186 <= 12'h1bc;
        src187 <= 12'h588;
        src188 <= 12'h876;
        exp <= 20'h5cd9e;
        #1
        src0 <= 12'h54b;
        src1 <= 12'h2ed;
        src2 <= 12'hf3;
        src3 <= 12'h1f4;
        src4 <= 12'hc3e;
        src5 <= 12'h52a;
        src6 <= 12'h7a4;
        src7 <= 12'h6a9;
        src8 <= 12'hf1e;
        src9 <= 12'hccf;
        src10 <= 12'h482;
        src11 <= 12'hfcb;
        src12 <= 12'h17;
        src13 <= 12'h92;
        src14 <= 12'h96;
        src15 <= 12'hb9b;
        src16 <= 12'h67d;
        src17 <= 12'h45b;
        src18 <= 12'h396;
        src19 <= 12'h337;
        src20 <= 12'hcf3;
        src21 <= 12'hff;
        src22 <= 12'hf51;
        src23 <= 12'h18c;
        src24 <= 12'hbf1;
        src25 <= 12'h86d;
        src26 <= 12'h96f;
        src27 <= 12'h4d3;
        src28 <= 12'h995;
        src29 <= 12'ha68;
        src30 <= 12'h885;
        src31 <= 12'h709;
        src32 <= 12'h3c1;
        src33 <= 12'h257;
        src34 <= 12'hb86;
        src35 <= 12'hb78;
        src36 <= 12'h408;
        src37 <= 12'hf5f;
        src38 <= 12'hd58;
        src39 <= 12'h38;
        src40 <= 12'ha3f;
        src41 <= 12'h21e;
        src42 <= 12'h122;
        src43 <= 12'h4e;
        src44 <= 12'h214;
        src45 <= 12'hccc;
        src46 <= 12'hbc5;
        src47 <= 12'hd92;
        src48 <= 12'h84b;
        src49 <= 12'hfa6;
        src50 <= 12'hcf5;
        src51 <= 12'h305;
        src52 <= 12'ha2d;
        src53 <= 12'hadd;
        src54 <= 12'h9e;
        src55 <= 12'hea7;
        src56 <= 12'h97b;
        src57 <= 12'ha91;
        src58 <= 12'he20;
        src59 <= 12'hbd5;
        src60 <= 12'ha83;
        src61 <= 12'h427;
        src62 <= 12'hb87;
        src63 <= 12'hb3;
        src64 <= 12'h266;
        src65 <= 12'h63c;
        src66 <= 12'hce2;
        src67 <= 12'hb8e;
        src68 <= 12'hf2a;
        src69 <= 12'hf1f;
        src70 <= 12'h88d;
        src71 <= 12'hc36;
        src72 <= 12'h26d;
        src73 <= 12'ha4;
        src74 <= 12'hfc9;
        src75 <= 12'hc24;
        src76 <= 12'h743;
        src77 <= 12'h919;
        src78 <= 12'hd56;
        src79 <= 12'hd88;
        src80 <= 12'hbb1;
        src81 <= 12'h18a;
        src82 <= 12'hafa;
        src83 <= 12'h7da;
        src84 <= 12'h14e;
        src85 <= 12'hcfd;
        src86 <= 12'h236;
        src87 <= 12'h756;
        src88 <= 12'h4c7;
        src89 <= 12'h1cb;
        src90 <= 12'h603;
        src91 <= 12'h11;
        src92 <= 12'h870;
        src93 <= 12'hbb4;
        src94 <= 12'h22a;
        src95 <= 12'h725;
        src96 <= 12'h9b6;
        src97 <= 12'h8a;
        src98 <= 12'hbc0;
        src99 <= 12'h26e;
        src100 <= 12'he6f;
        src101 <= 12'h60;
        src102 <= 12'h33f;
        src103 <= 12'hd84;
        src104 <= 12'hfe3;
        src105 <= 12'hdc2;
        src106 <= 12'ha1;
        src107 <= 12'he51;
        src108 <= 12'hbcf;
        src109 <= 12'h8f7;
        src110 <= 12'h599;
        src111 <= 12'he03;
        src112 <= 12'hcc2;
        src113 <= 12'h6ce;
        src114 <= 12'ha;
        src115 <= 12'h736;
        src116 <= 12'hb41;
        src117 <= 12'h429;
        src118 <= 12'h23b;
        src119 <= 12'hed7;
        src120 <= 12'h9d9;
        src121 <= 12'h30a;
        src122 <= 12'h188;
        src123 <= 12'he30;
        src124 <= 12'h649;
        src125 <= 12'h946;
        src126 <= 12'h645;
        src127 <= 12'h110;
        src128 <= 12'h906;
        src129 <= 12'hc38;
        src130 <= 12'hc43;
        src131 <= 12'hdd7;
        src132 <= 12'h7ff;
        src133 <= 12'had9;
        src134 <= 12'h98a;
        src135 <= 12'h6c5;
        src136 <= 12'hb1e;
        src137 <= 12'hd45;
        src138 <= 12'hba;
        src139 <= 12'h5ec;
        src140 <= 12'h4dd;
        src141 <= 12'hc0c;
        src142 <= 12'h997;
        src143 <= 12'h98e;
        src144 <= 12'hd49;
        src145 <= 12'hd8b;
        src146 <= 12'h176;
        src147 <= 12'h728;
        src148 <= 12'h9fb;
        src149 <= 12'hd3e;
        src150 <= 12'h93d;
        src151 <= 12'hbe;
        src152 <= 12'h3fc;
        src153 <= 12'hc57;
        src154 <= 12'h286;
        src155 <= 12'h648;
        src156 <= 12'h7ba;
        src157 <= 12'ha30;
        src158 <= 12'h28b;
        src159 <= 12'h4c7;
        src160 <= 12'ha10;
        src161 <= 12'hc2f;
        src162 <= 12'h1d5;
        src163 <= 12'hbd6;
        src164 <= 12'h92e;
        src165 <= 12'h49a;
        src166 <= 12'h99f;
        src167 <= 12'h77d;
        src168 <= 12'hc68;
        src169 <= 12'he78;
        src170 <= 12'h469;
        src171 <= 12'h7a6;
        src172 <= 12'h9e2;
        src173 <= 12'h131;
        src174 <= 12'h4bb;
        src175 <= 12'ha0;
        src176 <= 12'h1ff;
        src177 <= 12'hea6;
        src178 <= 12'hf90;
        src179 <= 12'hf28;
        src180 <= 12'h669;
        src181 <= 12'h3e5;
        src182 <= 12'h6b1;
        src183 <= 12'h792;
        src184 <= 12'h22a;
        src185 <= 12'hc92;
        src186 <= 12'hd3;
        src187 <= 12'h44f;
        src188 <= 12'hdce;
        exp <= 20'h5d42e;
        #1
        src0 <= 12'haa7;
        src1 <= 12'h1cb;
        src2 <= 12'h46a;
        src3 <= 12'h4e5;
        src4 <= 12'hc84;
        src5 <= 12'h4e8;
        src6 <= 12'h2fb;
        src7 <= 12'h58e;
        src8 <= 12'h6cb;
        src9 <= 12'h7c9;
        src10 <= 12'h33a;
        src11 <= 12'hcf;
        src12 <= 12'h269;
        src13 <= 12'h30d;
        src14 <= 12'h42f;
        src15 <= 12'h38f;
        src16 <= 12'hb8;
        src17 <= 12'h8d4;
        src18 <= 12'h7ac;
        src19 <= 12'he14;
        src20 <= 12'h43d;
        src21 <= 12'h74a;
        src22 <= 12'h21;
        src23 <= 12'h594;
        src24 <= 12'h982;
        src25 <= 12'h616;
        src26 <= 12'h294;
        src27 <= 12'h1a;
        src28 <= 12'hdf;
        src29 <= 12'h176;
        src30 <= 12'h4b2;
        src31 <= 12'hfec;
        src32 <= 12'h47d;
        src33 <= 12'hb4a;
        src34 <= 12'he98;
        src35 <= 12'hdb2;
        src36 <= 12'ha2e;
        src37 <= 12'hd99;
        src38 <= 12'h48a;
        src39 <= 12'h4fa;
        src40 <= 12'h3e7;
        src41 <= 12'h452;
        src42 <= 12'he87;
        src43 <= 12'haba;
        src44 <= 12'h88d;
        src45 <= 12'h9e7;
        src46 <= 12'he6f;
        src47 <= 12'hfc6;
        src48 <= 12'h3e9;
        src49 <= 12'h715;
        src50 <= 12'h482;
        src51 <= 12'hd58;
        src52 <= 12'hedb;
        src53 <= 12'h452;
        src54 <= 12'ha84;
        src55 <= 12'h442;
        src56 <= 12'h975;
        src57 <= 12'he8f;
        src58 <= 12'h2fe;
        src59 <= 12'h916;
        src60 <= 12'h670;
        src61 <= 12'h66e;
        src62 <= 12'h9b;
        src63 <= 12'h254;
        src64 <= 12'hec6;
        src65 <= 12'h8d9;
        src66 <= 12'h344;
        src67 <= 12'h4a2;
        src68 <= 12'h8d6;
        src69 <= 12'h7b6;
        src70 <= 12'h885;
        src71 <= 12'h829;
        src72 <= 12'h70a;
        src73 <= 12'hbda;
        src74 <= 12'h605;
        src75 <= 12'h744;
        src76 <= 12'h5af;
        src77 <= 12'h2e0;
        src78 <= 12'hd81;
        src79 <= 12'h2ae;
        src80 <= 12'hfe2;
        src81 <= 12'hf90;
        src82 <= 12'haed;
        src83 <= 12'h45;
        src84 <= 12'h2ef;
        src85 <= 12'hca0;
        src86 <= 12'h138;
        src87 <= 12'h540;
        src88 <= 12'hcc2;
        src89 <= 12'h8a5;
        src90 <= 12'h30;
        src91 <= 12'h705;
        src92 <= 12'hf75;
        src93 <= 12'hccc;
        src94 <= 12'hb60;
        src95 <= 12'hdc3;
        src96 <= 12'haea;
        src97 <= 12'h749;
        src98 <= 12'h785;
        src99 <= 12'hb5e;
        src100 <= 12'h69a;
        src101 <= 12'h300;
        src102 <= 12'hda6;
        src103 <= 12'hbbd;
        src104 <= 12'h826;
        src105 <= 12'h9e5;
        src106 <= 12'hff6;
        src107 <= 12'h24d;
        src108 <= 12'hf0e;
        src109 <= 12'hd10;
        src110 <= 12'h7fd;
        src111 <= 12'hb52;
        src112 <= 12'h2be;
        src113 <= 12'h42f;
        src114 <= 12'ha79;
        src115 <= 12'hcf1;
        src116 <= 12'hb7d;
        src117 <= 12'h8be;
        src118 <= 12'h63c;
        src119 <= 12'h749;
        src120 <= 12'hb40;
        src121 <= 12'hc0b;
        src122 <= 12'h283;
        src123 <= 12'h9d0;
        src124 <= 12'h557;
        src125 <= 12'hea;
        src126 <= 12'h700;
        src127 <= 12'h775;
        src128 <= 12'hf78;
        src129 <= 12'hb5a;
        src130 <= 12'hd2c;
        src131 <= 12'hc36;
        src132 <= 12'hcc5;
        src133 <= 12'h95d;
        src134 <= 12'h52b;
        src135 <= 12'h850;
        src136 <= 12'h88c;
        src137 <= 12'h7ad;
        src138 <= 12'hafc;
        src139 <= 12'h6c9;
        src140 <= 12'h9f6;
        src141 <= 12'hb1e;
        src142 <= 12'he95;
        src143 <= 12'h7d4;
        src144 <= 12'h6f6;
        src145 <= 12'h421;
        src146 <= 12'h2a4;
        src147 <= 12'hf3b;
        src148 <= 12'hba7;
        src149 <= 12'h6a3;
        src150 <= 12'hc2;
        src151 <= 12'h31b;
        src152 <= 12'hfdc;
        src153 <= 12'hd16;
        src154 <= 12'h21;
        src155 <= 12'h371;
        src156 <= 12'hd76;
        src157 <= 12'h274;
        src158 <= 12'h413;
        src159 <= 12'hf1c;
        src160 <= 12'h4a9;
        src161 <= 12'h610;
        src162 <= 12'hf4d;
        src163 <= 12'h28f;
        src164 <= 12'hdac;
        src165 <= 12'h5e0;
        src166 <= 12'h6f6;
        src167 <= 12'ha75;
        src168 <= 12'h8e2;
        src169 <= 12'hc4a;
        src170 <= 12'h4c0;
        src171 <= 12'h23c;
        src172 <= 12'h501;
        src173 <= 12'hefe;
        src174 <= 12'h50c;
        src175 <= 12'h853;
        src176 <= 12'h143;
        src177 <= 12'h167;
        src178 <= 12'h45d;
        src179 <= 12'hbdf;
        src180 <= 12'h23b;
        src181 <= 12'h6e8;
        src182 <= 12'h640;
        src183 <= 12'h992;
        src184 <= 12'h448;
        src185 <= 12'hc5b;
        src186 <= 12'h5d6;
        src187 <= 12'hbe5;
        src188 <= 12'hfad;
        exp <= 20'h5d503;
        #1
        src0 <= 12'h78e;
        src1 <= 12'h8e6;
        src2 <= 12'h76c;
        src3 <= 12'h33;
        src4 <= 12'h5bb;
        src5 <= 12'hf33;
        src6 <= 12'h950;
        src7 <= 12'h28b;
        src8 <= 12'hba3;
        src9 <= 12'hb31;
        src10 <= 12'h65a;
        src11 <= 12'h4c8;
        src12 <= 12'hcb3;
        src13 <= 12'h925;
        src14 <= 12'h31f;
        src15 <= 12'h3e4;
        src16 <= 12'h19;
        src17 <= 12'h502;
        src18 <= 12'h80c;
        src19 <= 12'h612;
        src20 <= 12'hae6;
        src21 <= 12'h139;
        src22 <= 12'h607;
        src23 <= 12'h87b;
        src24 <= 12'hd9d;
        src25 <= 12'h181;
        src26 <= 12'h886;
        src27 <= 12'hf9a;
        src28 <= 12'hf34;
        src29 <= 12'h993;
        src30 <= 12'hefe;
        src31 <= 12'hafa;
        src32 <= 12'hf7b;
        src33 <= 12'h264;
        src34 <= 12'h727;
        src35 <= 12'hcc0;
        src36 <= 12'h81d;
        src37 <= 12'hc5;
        src38 <= 12'h73e;
        src39 <= 12'ha24;
        src40 <= 12'h724;
        src41 <= 12'hbd5;
        src42 <= 12'hb48;
        src43 <= 12'ha37;
        src44 <= 12'h92;
        src45 <= 12'h777;
        src46 <= 12'h117;
        src47 <= 12'hf79;
        src48 <= 12'h426;
        src49 <= 12'h82;
        src50 <= 12'h530;
        src51 <= 12'h79d;
        src52 <= 12'h35d;
        src53 <= 12'h96b;
        src54 <= 12'hed9;
        src55 <= 12'hac2;
        src56 <= 12'h599;
        src57 <= 12'h5d5;
        src58 <= 12'had5;
        src59 <= 12'ha2a;
        src60 <= 12'h563;
        src61 <= 12'he9f;
        src62 <= 12'he19;
        src63 <= 12'h9fc;
        src64 <= 12'h80d;
        src65 <= 12'h60f;
        src66 <= 12'h438;
        src67 <= 12'hed;
        src68 <= 12'h61d;
        src69 <= 12'hb6c;
        src70 <= 12'h92c;
        src71 <= 12'h610;
        src72 <= 12'hfa7;
        src73 <= 12'h924;
        src74 <= 12'h460;
        src75 <= 12'h21f;
        src76 <= 12'hee2;
        src77 <= 12'h7be;
        src78 <= 12'h9ea;
        src79 <= 12'hf01;
        src80 <= 12'hc35;
        src81 <= 12'hf67;
        src82 <= 12'hc46;
        src83 <= 12'h299;
        src84 <= 12'hfb2;
        src85 <= 12'h929;
        src86 <= 12'h577;
        src87 <= 12'hdbe;
        src88 <= 12'h9d4;
        src89 <= 12'h6d5;
        src90 <= 12'hd77;
        src91 <= 12'ha4f;
        src92 <= 12'h48;
        src93 <= 12'h9df;
        src94 <= 12'h423;
        src95 <= 12'h508;
        src96 <= 12'h949;
        src97 <= 12'hd43;
        src98 <= 12'hea1;
        src99 <= 12'h446;
        src100 <= 12'hb42;
        src101 <= 12'h3a;
        src102 <= 12'hfab;
        src103 <= 12'h1ba;
        src104 <= 12'hc3a;
        src105 <= 12'h59b;
        src106 <= 12'h93c;
        src107 <= 12'hfdc;
        src108 <= 12'h553;
        src109 <= 12'h61b;
        src110 <= 12'hbe8;
        src111 <= 12'h8cc;
        src112 <= 12'h133;
        src113 <= 12'hcc9;
        src114 <= 12'h8fe;
        src115 <= 12'hb0b;
        src116 <= 12'he03;
        src117 <= 12'hfee;
        src118 <= 12'h376;
        src119 <= 12'h5fd;
        src120 <= 12'hf2d;
        src121 <= 12'h860;
        src122 <= 12'h251;
        src123 <= 12'hc0f;
        src124 <= 12'hd3;
        src125 <= 12'h62a;
        src126 <= 12'h5ee;
        src127 <= 12'h536;
        src128 <= 12'h39d;
        src129 <= 12'h3a5;
        src130 <= 12'h992;
        src131 <= 12'h1bd;
        src132 <= 12'h800;
        src133 <= 12'haa0;
        src134 <= 12'hcd2;
        src135 <= 12'h604;
        src136 <= 12'h670;
        src137 <= 12'h94e;
        src138 <= 12'h777;
        src139 <= 12'he0d;
        src140 <= 12'h48c;
        src141 <= 12'h55b;
        src142 <= 12'h983;
        src143 <= 12'h95c;
        src144 <= 12'h663;
        src145 <= 12'h44e;
        src146 <= 12'h7c0;
        src147 <= 12'had;
        src148 <= 12'ha68;
        src149 <= 12'haf6;
        src150 <= 12'h169;
        src151 <= 12'h330;
        src152 <= 12'hb1d;
        src153 <= 12'hbf;
        src154 <= 12'h6ac;
        src155 <= 12'h438;
        src156 <= 12'hcad;
        src157 <= 12'h256;
        src158 <= 12'h482;
        src159 <= 12'h20;
        src160 <= 12'h2bd;
        src161 <= 12'h390;
        src162 <= 12'h8d2;
        src163 <= 12'h10c;
        src164 <= 12'h3a9;
        src165 <= 12'hff2;
        src166 <= 12'h446;
        src167 <= 12'he0e;
        src168 <= 12'h844;
        src169 <= 12'hf20;
        src170 <= 12'h2aa;
        src171 <= 12'h5ee;
        src172 <= 12'hc40;
        src173 <= 12'h750;
        src174 <= 12'hcb;
        src175 <= 12'hf3e;
        src176 <= 12'h616;
        src177 <= 12'h345;
        src178 <= 12'hf56;
        src179 <= 12'h31;
        src180 <= 12'heba;
        src181 <= 12'h35a;
        src182 <= 12'h454;
        src183 <= 12'h591;
        src184 <= 12'h8e;
        src185 <= 12'h2ba;
        src186 <= 12'h679;
        src187 <= 12'h3e0;
        src188 <= 12'hfe4;
        exp <= 20'h5ca94;
        #1
        src0 <= 12'h9ab;
        src1 <= 12'h7b1;
        src2 <= 12'h6b6;
        src3 <= 12'h203;
        src4 <= 12'h4b3;
        src5 <= 12'h71e;
        src6 <= 12'h258;
        src7 <= 12'h44d;
        src8 <= 12'hcf0;
        src9 <= 12'h594;
        src10 <= 12'h62b;
        src11 <= 12'hc21;
        src12 <= 12'hee5;
        src13 <= 12'ha07;
        src14 <= 12'h31a;
        src15 <= 12'hdfa;
        src16 <= 12'hded;
        src17 <= 12'heac;
        src18 <= 12'ha2a;
        src19 <= 12'hf66;
        src20 <= 12'hf2e;
        src21 <= 12'heb4;
        src22 <= 12'h883;
        src23 <= 12'h371;
        src24 <= 12'h72;
        src25 <= 12'h9e;
        src26 <= 12'he18;
        src27 <= 12'hfd7;
        src28 <= 12'hb24;
        src29 <= 12'hca3;
        src30 <= 12'h9d6;
        src31 <= 12'h84e;
        src32 <= 12'h24a;
        src33 <= 12'h7ca;
        src34 <= 12'h8ed;
        src35 <= 12'hff6;
        src36 <= 12'h8d4;
        src37 <= 12'h79;
        src38 <= 12'hb38;
        src39 <= 12'h512;
        src40 <= 12'h543;
        src41 <= 12'h889;
        src42 <= 12'h1b5;
        src43 <= 12'h4aa;
        src44 <= 12'hb8a;
        src45 <= 12'h670;
        src46 <= 12'h80e;
        src47 <= 12'hd27;
        src48 <= 12'h523;
        src49 <= 12'hf5;
        src50 <= 12'hb13;
        src51 <= 12'h384;
        src52 <= 12'hb9f;
        src53 <= 12'h30;
        src54 <= 12'hbd5;
        src55 <= 12'h8ca;
        src56 <= 12'hcf8;
        src57 <= 12'hc03;
        src58 <= 12'h312;
        src59 <= 12'h96c;
        src60 <= 12'h14;
        src61 <= 12'h873;
        src62 <= 12'hc86;
        src63 <= 12'hb77;
        src64 <= 12'h17a;
        src65 <= 12'he0a;
        src66 <= 12'hd9a;
        src67 <= 12'hcb4;
        src68 <= 12'hd60;
        src69 <= 12'hef9;
        src70 <= 12'hc22;
        src71 <= 12'hdd;
        src72 <= 12'h68a;
        src73 <= 12'h579;
        src74 <= 12'h8ef;
        src75 <= 12'he33;
        src76 <= 12'hce6;
        src77 <= 12'h53e;
        src78 <= 12'h90d;
        src79 <= 12'h4d7;
        src80 <= 12'h67;
        src81 <= 12'h83a;
        src82 <= 12'h83b;
        src83 <= 12'hd50;
        src84 <= 12'hb7d;
        src85 <= 12'h5ea;
        src86 <= 12'h98f;
        src87 <= 12'h11b;
        src88 <= 12'h70e;
        src89 <= 12'hb6e;
        src90 <= 12'haaa;
        src91 <= 12'hc79;
        src92 <= 12'h75d;
        src93 <= 12'h324;
        src94 <= 12'h95e;
        src95 <= 12'hbf8;
        src96 <= 12'h630;
        src97 <= 12'hceb;
        src98 <= 12'h73c;
        src99 <= 12'h4d6;
        src100 <= 12'hcd5;
        src101 <= 12'hd2d;
        src102 <= 12'h768;
        src103 <= 12'h837;
        src104 <= 12'h51c;
        src105 <= 12'h2aa;
        src106 <= 12'hd31;
        src107 <= 12'ha48;
        src108 <= 12'h73d;
        src109 <= 12'hab2;
        src110 <= 12'h4c9;
        src111 <= 12'hbfe;
        src112 <= 12'h138;
        src113 <= 12'he04;
        src114 <= 12'h2cd;
        src115 <= 12'h239;
        src116 <= 12'h2ed;
        src117 <= 12'h2c7;
        src118 <= 12'hd05;
        src119 <= 12'h3e0;
        src120 <= 12'ha1a;
        src121 <= 12'ha78;
        src122 <= 12'h9ea;
        src123 <= 12'hcbc;
        src124 <= 12'hfe2;
        src125 <= 12'h40e;
        src126 <= 12'ha1b;
        src127 <= 12'hf74;
        src128 <= 12'h151;
        src129 <= 12'h42d;
        src130 <= 12'h66f;
        src131 <= 12'h335;
        src132 <= 12'h4b2;
        src133 <= 12'h9e9;
        src134 <= 12'hc06;
        src135 <= 12'hb69;
        src136 <= 12'hede;
        src137 <= 12'h6f3;
        src138 <= 12'hf86;
        src139 <= 12'hcfc;
        src140 <= 12'h899;
        src141 <= 12'hf68;
        src142 <= 12'h2d2;
        src143 <= 12'h1cd;
        src144 <= 12'hdc6;
        src145 <= 12'hd03;
        src146 <= 12'h7e;
        src147 <= 12'h8e8;
        src148 <= 12'hd50;
        src149 <= 12'hf3d;
        src150 <= 12'hf95;
        src151 <= 12'h6d2;
        src152 <= 12'ha2e;
        src153 <= 12'h88b;
        src154 <= 12'h92f;
        src155 <= 12'h65;
        src156 <= 12'h3d6;
        src157 <= 12'h42b;
        src158 <= 12'h92c;
        src159 <= 12'h220;
        src160 <= 12'h979;
        src161 <= 12'h1ed;
        src162 <= 12'hd36;
        src163 <= 12'h4c4;
        src164 <= 12'h673;
        src165 <= 12'h3c7;
        src166 <= 12'hadf;
        src167 <= 12'hb09;
        src168 <= 12'hb9a;
        src169 <= 12'hb5e;
        src170 <= 12'h66b;
        src171 <= 12'hbf1;
        src172 <= 12'h1e5;
        src173 <= 12'hb98;
        src174 <= 12'hfac;
        src175 <= 12'h885;
        src176 <= 12'hbef;
        src177 <= 12'hbf0;
        src178 <= 12'h450;
        src179 <= 12'hc8d;
        src180 <= 12'hd4d;
        src181 <= 12'he11;
        src182 <= 12'hf25;
        src183 <= 12'h107;
        src184 <= 12'h6bc;
        src185 <= 12'hb02;
        src186 <= 12'hf78;
        src187 <= 12'h594;
        src188 <= 12'hdbe;
        exp <= 20'h65fd3;
        #1
        src0 <= 12'h5b8;
        src1 <= 12'h3ba;
        src2 <= 12'h8e0;
        src3 <= 12'hc4e;
        src4 <= 12'h32f;
        src5 <= 12'h12f;
        src6 <= 12'hf52;
        src7 <= 12'hc70;
        src8 <= 12'h603;
        src9 <= 12'h167;
        src10 <= 12'hf5b;
        src11 <= 12'h124;
        src12 <= 12'h520;
        src13 <= 12'hb10;
        src14 <= 12'h9d2;
        src15 <= 12'h47a;
        src16 <= 12'hd1d;
        src17 <= 12'h22f;
        src18 <= 12'hb03;
        src19 <= 12'h3b1;
        src20 <= 12'h250;
        src21 <= 12'h8b1;
        src22 <= 12'h7d8;
        src23 <= 12'he60;
        src24 <= 12'h209;
        src25 <= 12'h734;
        src26 <= 12'h995;
        src27 <= 12'h114;
        src28 <= 12'h704;
        src29 <= 12'he41;
        src30 <= 12'hfd5;
        src31 <= 12'he7b;
        src32 <= 12'h81c;
        src33 <= 12'h693;
        src34 <= 12'he5d;
        src35 <= 12'h487;
        src36 <= 12'h33a;
        src37 <= 12'h661;
        src38 <= 12'h553;
        src39 <= 12'h394;
        src40 <= 12'h51e;
        src41 <= 12'hfdf;
        src42 <= 12'he06;
        src43 <= 12'h548;
        src44 <= 12'he07;
        src45 <= 12'h4f1;
        src46 <= 12'hd35;
        src47 <= 12'h4c3;
        src48 <= 12'h4af;
        src49 <= 12'hbb8;
        src50 <= 12'h727;
        src51 <= 12'hfa2;
        src52 <= 12'h7e;
        src53 <= 12'h364;
        src54 <= 12'hda7;
        src55 <= 12'h767;
        src56 <= 12'ha8d;
        src57 <= 12'h3d2;
        src58 <= 12'h445;
        src59 <= 12'hdc3;
        src60 <= 12'h7d;
        src61 <= 12'he01;
        src62 <= 12'h7ba;
        src63 <= 12'h706;
        src64 <= 12'h4dd;
        src65 <= 12'hac0;
        src66 <= 12'hf1e;
        src67 <= 12'h3c9;
        src68 <= 12'h776;
        src69 <= 12'h4b0;
        src70 <= 12'h78c;
        src71 <= 12'h8a5;
        src72 <= 12'hc5e;
        src73 <= 12'h44d;
        src74 <= 12'h38b;
        src75 <= 12'he6c;
        src76 <= 12'h21;
        src77 <= 12'hd4a;
        src78 <= 12'he00;
        src79 <= 12'hbd3;
        src80 <= 12'h6bb;
        src81 <= 12'hf59;
        src82 <= 12'h6cf;
        src83 <= 12'hf66;
        src84 <= 12'hcc5;
        src85 <= 12'h393;
        src86 <= 12'h493;
        src87 <= 12'hd25;
        src88 <= 12'hb4b;
        src89 <= 12'h303;
        src90 <= 12'h2e6;
        src91 <= 12'h69f;
        src92 <= 12'h1b;
        src93 <= 12'hb7a;
        src94 <= 12'he7d;
        src95 <= 12'hd95;
        src96 <= 12'h1cb;
        src97 <= 12'h41f;
        src98 <= 12'hf0c;
        src99 <= 12'h657;
        src100 <= 12'h5a1;
        src101 <= 12'h9eb;
        src102 <= 12'h3df;
        src103 <= 12'hd9f;
        src104 <= 12'hcef;
        src105 <= 12'h4a0;
        src106 <= 12'h719;
        src107 <= 12'h661;
        src108 <= 12'h49a;
        src109 <= 12'he53;
        src110 <= 12'h28c;
        src111 <= 12'h4f0;
        src112 <= 12'he4c;
        src113 <= 12'h5cb;
        src114 <= 12'h2eb;
        src115 <= 12'hf2;
        src116 <= 12'h4f1;
        src117 <= 12'h735;
        src118 <= 12'hdc1;
        src119 <= 12'hde7;
        src120 <= 12'h6f8;
        src121 <= 12'h2d5;
        src122 <= 12'h26;
        src123 <= 12'h566;
        src124 <= 12'h177;
        src125 <= 12'h966;
        src126 <= 12'hebc;
        src127 <= 12'hba3;
        src128 <= 12'h6c4;
        src129 <= 12'h62d;
        src130 <= 12'hf8c;
        src131 <= 12'h42;
        src132 <= 12'hd66;
        src133 <= 12'h3ee;
        src134 <= 12'h8ce;
        src135 <= 12'hd76;
        src136 <= 12'hec1;
        src137 <= 12'hd0a;
        src138 <= 12'h6ab;
        src139 <= 12'hef2;
        src140 <= 12'h6ab;
        src141 <= 12'he59;
        src142 <= 12'h543;
        src143 <= 12'h2f;
        src144 <= 12'he68;
        src145 <= 12'h84;
        src146 <= 12'h3c3;
        src147 <= 12'he48;
        src148 <= 12'h4d9;
        src149 <= 12'hf78;
        src150 <= 12'hc5c;
        src151 <= 12'hf8f;
        src152 <= 12'h768;
        src153 <= 12'h83b;
        src154 <= 12'h928;
        src155 <= 12'h4b5;
        src156 <= 12'h5f2;
        src157 <= 12'h32f;
        src158 <= 12'h7f0;
        src159 <= 12'hfc3;
        src160 <= 12'h4ea;
        src161 <= 12'h95f;
        src162 <= 12'he6c;
        src163 <= 12'hbfe;
        src164 <= 12'h16d;
        src165 <= 12'hbc0;
        src166 <= 12'ha32;
        src167 <= 12'hfcc;
        src168 <= 12'h559;
        src169 <= 12'hb24;
        src170 <= 12'h21a;
        src171 <= 12'h603;
        src172 <= 12'h5f5;
        src173 <= 12'hac8;
        src174 <= 12'h84a;
        src175 <= 12'h774;
        src176 <= 12'hbb7;
        src177 <= 12'h534;
        src178 <= 12'ha8f;
        src179 <= 12'h21d;
        src180 <= 12'h72a;
        src181 <= 12'h70c;
        src182 <= 12'h9a4;
        src183 <= 12'h837;
        src184 <= 12'hb41;
        src185 <= 12'h93d;
        src186 <= 12'h521;
        src187 <= 12'h311;
        src188 <= 12'h813;
        exp <= 20'h606b6;
        #1
        src0 <= 12'hdda;
        src1 <= 12'hca8;
        src2 <= 12'hccb;
        src3 <= 12'hcd4;
        src4 <= 12'hcbf;
        src5 <= 12'hb9c;
        src6 <= 12'h9e5;
        src7 <= 12'hdf4;
        src8 <= 12'hca;
        src9 <= 12'h47f;
        src10 <= 12'h14f;
        src11 <= 12'he51;
        src12 <= 12'h405;
        src13 <= 12'h7cc;
        src14 <= 12'h6d9;
        src15 <= 12'h890;
        src16 <= 12'h159;
        src17 <= 12'h5f5;
        src18 <= 12'h51c;
        src19 <= 12'h2af;
        src20 <= 12'h8;
        src21 <= 12'h472;
        src22 <= 12'h89;
        src23 <= 12'hafa;
        src24 <= 12'h296;
        src25 <= 12'ha60;
        src26 <= 12'h90d;
        src27 <= 12'h3d;
        src28 <= 12'h494;
        src29 <= 12'h46c;
        src30 <= 12'hd6b;
        src31 <= 12'hd05;
        src32 <= 12'h1a9;
        src33 <= 12'h4a;
        src34 <= 12'h28e;
        src35 <= 12'h485;
        src36 <= 12'hda2;
        src37 <= 12'h99f;
        src38 <= 12'hfd;
        src39 <= 12'h899;
        src40 <= 12'h5fc;
        src41 <= 12'hcd3;
        src42 <= 12'heee;
        src43 <= 12'haab;
        src44 <= 12'h16;
        src45 <= 12'h947;
        src46 <= 12'hb47;
        src47 <= 12'h1e0;
        src48 <= 12'hc7d;
        src49 <= 12'h1db;
        src50 <= 12'h31b;
        src51 <= 12'h385;
        src52 <= 12'hb2d;
        src53 <= 12'hb3f;
        src54 <= 12'hd9d;
        src55 <= 12'hf26;
        src56 <= 12'hd79;
        src57 <= 12'h21f;
        src58 <= 12'hab;
        src59 <= 12'hfcb;
        src60 <= 12'hb01;
        src61 <= 12'h3dc;
        src62 <= 12'hf29;
        src63 <= 12'h733;
        src64 <= 12'hfdd;
        src65 <= 12'h570;
        src66 <= 12'h829;
        src67 <= 12'h183;
        src68 <= 12'hd11;
        src69 <= 12'he22;
        src70 <= 12'h98d;
        src71 <= 12'hbd0;
        src72 <= 12'h4cc;
        src73 <= 12'hbfa;
        src74 <= 12'hc25;
        src75 <= 12'hf6;
        src76 <= 12'h1cf;
        src77 <= 12'h46;
        src78 <= 12'h2e0;
        src79 <= 12'hdc;
        src80 <= 12'he2b;
        src81 <= 12'h1d5;
        src82 <= 12'hf58;
        src83 <= 12'hd3a;
        src84 <= 12'h99b;
        src85 <= 12'ha3a;
        src86 <= 12'hbfd;
        src87 <= 12'haf5;
        src88 <= 12'h3cc;
        src89 <= 12'h2f1;
        src90 <= 12'he03;
        src91 <= 12'h452;
        src92 <= 12'h301;
        src93 <= 12'hb66;
        src94 <= 12'h371;
        src95 <= 12'h46e;
        src96 <= 12'h9c5;
        src97 <= 12'had;
        src98 <= 12'h70d;
        src99 <= 12'h62;
        src100 <= 12'ha89;
        src101 <= 12'h794;
        src102 <= 12'h814;
        src103 <= 12'hb71;
        src104 <= 12'h830;
        src105 <= 12'h592;
        src106 <= 12'h8c0;
        src107 <= 12'h609;
        src108 <= 12'h18a;
        src109 <= 12'h8d0;
        src110 <= 12'hc36;
        src111 <= 12'hd2;
        src112 <= 12'h621;
        src113 <= 12'h239;
        src114 <= 12'he90;
        src115 <= 12'hfda;
        src116 <= 12'hca9;
        src117 <= 12'h4f0;
        src118 <= 12'h51d;
        src119 <= 12'h3c2;
        src120 <= 12'hf02;
        src121 <= 12'he50;
        src122 <= 12'he0e;
        src123 <= 12'hf9;
        src124 <= 12'ha4c;
        src125 <= 12'hd19;
        src126 <= 12'hf1b;
        src127 <= 12'h3db;
        src128 <= 12'hff5;
        src129 <= 12'hb02;
        src130 <= 12'h126;
        src131 <= 12'h2ce;
        src132 <= 12'h1f;
        src133 <= 12'h291;
        src134 <= 12'ha39;
        src135 <= 12'h39c;
        src136 <= 12'h23;
        src137 <= 12'hfbb;
        src138 <= 12'ha1e;
        src139 <= 12'h7ce;
        src140 <= 12'hfa9;
        src141 <= 12'h7d7;
        src142 <= 12'h124;
        src143 <= 12'h33d;
        src144 <= 12'h260;
        src145 <= 12'h530;
        src146 <= 12'h42b;
        src147 <= 12'hdba;
        src148 <= 12'ha2a;
        src149 <= 12'h228;
        src150 <= 12'h14;
        src151 <= 12'h14c;
        src152 <= 12'h8d2;
        src153 <= 12'hd4b;
        src154 <= 12'hc5;
        src155 <= 12'h75f;
        src156 <= 12'h81a;
        src157 <= 12'h53f;
        src158 <= 12'h77d;
        src159 <= 12'hcec;
        src160 <= 12'hecc;
        src161 <= 12'h390;
        src162 <= 12'h7f7;
        src163 <= 12'h9e8;
        src164 <= 12'hbf;
        src165 <= 12'he43;
        src166 <= 12'hc8e;
        src167 <= 12'ha8c;
        src168 <= 12'h8cb;
        src169 <= 12'h55a;
        src170 <= 12'h8e3;
        src171 <= 12'h6db;
        src172 <= 12'h48d;
        src173 <= 12'h21e;
        src174 <= 12'hf74;
        src175 <= 12'ha;
        src176 <= 12'h72b;
        src177 <= 12'h7d9;
        src178 <= 12'ha30;
        src179 <= 12'h6d0;
        src180 <= 12'hefd;
        src181 <= 12'h923;
        src182 <= 12'h7f5;
        src183 <= 12'h963;
        src184 <= 12'h5af;
        src185 <= 12'h92e;
        src186 <= 12'h116;
        src187 <= 12'ha62;
        src188 <= 12'hda5;
        exp <= 20'h5a8df;
        #1
        src0 <= 12'h532;
        src1 <= 12'h8d5;
        src2 <= 12'h7eb;
        src3 <= 12'h944;
        src4 <= 12'h3d6;
        src5 <= 12'hba;
        src6 <= 12'h9ed;
        src7 <= 12'ha74;
        src8 <= 12'hd23;
        src9 <= 12'h5ac;
        src10 <= 12'h1ef;
        src11 <= 12'h57;
        src12 <= 12'ha1c;
        src13 <= 12'h938;
        src14 <= 12'h392;
        src15 <= 12'hb53;
        src16 <= 12'h4b2;
        src17 <= 12'hf49;
        src18 <= 12'h8b9;
        src19 <= 12'h12c;
        src20 <= 12'h11b;
        src21 <= 12'h85b;
        src22 <= 12'hf89;
        src23 <= 12'he3e;
        src24 <= 12'ha39;
        src25 <= 12'h118;
        src26 <= 12'h163;
        src27 <= 12'h4f5;
        src28 <= 12'h859;
        src29 <= 12'he34;
        src30 <= 12'h13c;
        src31 <= 12'hcb8;
        src32 <= 12'h9dc;
        src33 <= 12'h4b;
        src34 <= 12'h516;
        src35 <= 12'ha99;
        src36 <= 12'h7e;
        src37 <= 12'hf03;
        src38 <= 12'hc03;
        src39 <= 12'h1d3;
        src40 <= 12'hc92;
        src41 <= 12'h331;
        src42 <= 12'hc9d;
        src43 <= 12'h951;
        src44 <= 12'hcbd;
        src45 <= 12'h625;
        src46 <= 12'h9cd;
        src47 <= 12'h20d;
        src48 <= 12'h8bd;
        src49 <= 12'hf9d;
        src50 <= 12'h3ee;
        src51 <= 12'h42c;
        src52 <= 12'hd24;
        src53 <= 12'h4d6;
        src54 <= 12'hcad;
        src55 <= 12'h74e;
        src56 <= 12'h6d6;
        src57 <= 12'h9df;
        src58 <= 12'h70c;
        src59 <= 12'h905;
        src60 <= 12'h45b;
        src61 <= 12'hc01;
        src62 <= 12'hfb0;
        src63 <= 12'h39d;
        src64 <= 12'hfae;
        src65 <= 12'h4b1;
        src66 <= 12'h802;
        src67 <= 12'h7e1;
        src68 <= 12'h67b;
        src69 <= 12'he11;
        src70 <= 12'h37f;
        src71 <= 12'h112;
        src72 <= 12'h4d;
        src73 <= 12'h872;
        src74 <= 12'hc49;
        src75 <= 12'h349;
        src76 <= 12'h429;
        src77 <= 12'h8ba;
        src78 <= 12'hf51;
        src79 <= 12'h1df;
        src80 <= 12'he2e;
        src81 <= 12'hf99;
        src82 <= 12'h273;
        src83 <= 12'h1aa;
        src84 <= 12'h48c;
        src85 <= 12'hde7;
        src86 <= 12'h9e4;
        src87 <= 12'h7af;
        src88 <= 12'hec6;
        src89 <= 12'h966;
        src90 <= 12'hcd3;
        src91 <= 12'h100;
        src92 <= 12'h2bb;
        src93 <= 12'h237;
        src94 <= 12'h36c;
        src95 <= 12'h129;
        src96 <= 12'h5ba;
        src97 <= 12'hd66;
        src98 <= 12'h6f6;
        src99 <= 12'he4f;
        src100 <= 12'h16f;
        src101 <= 12'h853;
        src102 <= 12'h737;
        src103 <= 12'hde7;
        src104 <= 12'hce7;
        src105 <= 12'h2e2;
        src106 <= 12'hd25;
        src107 <= 12'h688;
        src108 <= 12'h2a0;
        src109 <= 12'h51;
        src110 <= 12'hbfe;
        src111 <= 12'hfcf;
        src112 <= 12'h829;
        src113 <= 12'h40e;
        src114 <= 12'h339;
        src115 <= 12'h30c;
        src116 <= 12'hc1d;
        src117 <= 12'hb2d;
        src118 <= 12'h893;
        src119 <= 12'he9b;
        src120 <= 12'hde4;
        src121 <= 12'h106;
        src122 <= 12'hc56;
        src123 <= 12'he0d;
        src124 <= 12'h812;
        src125 <= 12'h2c5;
        src126 <= 12'h2c5;
        src127 <= 12'hfaf;
        src128 <= 12'h620;
        src129 <= 12'h378;
        src130 <= 12'h3c3;
        src131 <= 12'h414;
        src132 <= 12'h7ee;
        src133 <= 12'h54e;
        src134 <= 12'h44b;
        src135 <= 12'h94c;
        src136 <= 12'h7cd;
        src137 <= 12'hafa;
        src138 <= 12'h7da;
        src139 <= 12'hef0;
        src140 <= 12'hb68;
        src141 <= 12'hd73;
        src142 <= 12'h4dc;
        src143 <= 12'h78e;
        src144 <= 12'h60a;
        src145 <= 12'hb2f;
        src146 <= 12'h6e8;
        src147 <= 12'h400;
        src148 <= 12'h749;
        src149 <= 12'h669;
        src150 <= 12'h247;
        src151 <= 12'h4af;
        src152 <= 12'h1a8;
        src153 <= 12'he36;
        src154 <= 12'h543;
        src155 <= 12'hfb1;
        src156 <= 12'h81c;
        src157 <= 12'hb7b;
        src158 <= 12'hfd3;
        src159 <= 12'hfaa;
        src160 <= 12'h26f;
        src161 <= 12'h39;
        src162 <= 12'hab7;
        src163 <= 12'h545;
        src164 <= 12'h3f2;
        src165 <= 12'hde3;
        src166 <= 12'h279;
        src167 <= 12'had8;
        src168 <= 12'ha87;
        src169 <= 12'h384;
        src170 <= 12'hb52;
        src171 <= 12'hacb;
        src172 <= 12'he1;
        src173 <= 12'h4f7;
        src174 <= 12'h970;
        src175 <= 12'h6fd;
        src176 <= 12'h968;
        src177 <= 12'hebe;
        src178 <= 12'h1ac;
        src179 <= 12'hcff;
        src180 <= 12'hd5a;
        src181 <= 12'h883;
        src182 <= 12'hc1;
        src183 <= 12'h87a;
        src184 <= 12'h870;
        src185 <= 12'h58b;
        src186 <= 12'hb56;
        src187 <= 12'h45c;
        src188 <= 12'h385;
        exp <= 20'h5c27f;
        #1
        src0 <= 12'h95d;
        src1 <= 12'h810;
        src2 <= 12'hb44;
        src3 <= 12'h2e4;
        src4 <= 12'h669;
        src5 <= 12'hc1f;
        src6 <= 12'h69e;
        src7 <= 12'h95b;
        src8 <= 12'h18a;
        src9 <= 12'he48;
        src10 <= 12'h9d6;
        src11 <= 12'hc0d;
        src12 <= 12'h15e;
        src13 <= 12'hb8b;
        src14 <= 12'he53;
        src15 <= 12'hd6b;
        src16 <= 12'h83;
        src17 <= 12'he2c;
        src18 <= 12'he15;
        src19 <= 12'hb73;
        src20 <= 12'h6e;
        src21 <= 12'h2b4;
        src22 <= 12'hda3;
        src23 <= 12'h353;
        src24 <= 12'hd6a;
        src25 <= 12'hcea;
        src26 <= 12'h593;
        src27 <= 12'hdc8;
        src28 <= 12'h3c7;
        src29 <= 12'hdc;
        src30 <= 12'h74;
        src31 <= 12'he95;
        src32 <= 12'hb15;
        src33 <= 12'h87;
        src34 <= 12'hb69;
        src35 <= 12'hc28;
        src36 <= 12'hafe;
        src37 <= 12'h57d;
        src38 <= 12'h3b4;
        src39 <= 12'h578;
        src40 <= 12'hb3;
        src41 <= 12'h2bd;
        src42 <= 12'h767;
        src43 <= 12'h3a;
        src44 <= 12'h4e7;
        src45 <= 12'hfea;
        src46 <= 12'h846;
        src47 <= 12'hf6b;
        src48 <= 12'he7f;
        src49 <= 12'h1c;
        src50 <= 12'h98f;
        src51 <= 12'h678;
        src52 <= 12'heff;
        src53 <= 12'h753;
        src54 <= 12'hd56;
        src55 <= 12'h9b3;
        src56 <= 12'hf0f;
        src57 <= 12'h4;
        src58 <= 12'hf46;
        src59 <= 12'habe;
        src60 <= 12'h7b6;
        src61 <= 12'h9a7;
        src62 <= 12'h295;
        src63 <= 12'h13;
        src64 <= 12'h830;
        src65 <= 12'hb69;
        src66 <= 12'h9bc;
        src67 <= 12'h253;
        src68 <= 12'hbf7;
        src69 <= 12'hc20;
        src70 <= 12'h456;
        src71 <= 12'hdf8;
        src72 <= 12'h44e;
        src73 <= 12'h661;
        src74 <= 12'hf54;
        src75 <= 12'hfda;
        src76 <= 12'h754;
        src77 <= 12'h10;
        src78 <= 12'h3fc;
        src79 <= 12'h812;
        src80 <= 12'h839;
        src81 <= 12'h57;
        src82 <= 12'habd;
        src83 <= 12'haa3;
        src84 <= 12'hff6;
        src85 <= 12'hf79;
        src86 <= 12'h8dc;
        src87 <= 12'h77e;
        src88 <= 12'hbc7;
        src89 <= 12'hcdd;
        src90 <= 12'heb2;
        src91 <= 12'hba7;
        src92 <= 12'h749;
        src93 <= 12'hcc2;
        src94 <= 12'h461;
        src95 <= 12'hcb;
        src96 <= 12'h8dd;
        src97 <= 12'h876;
        src98 <= 12'hae9;
        src99 <= 12'hb54;
        src100 <= 12'h898;
        src101 <= 12'h797;
        src102 <= 12'h8ea;
        src103 <= 12'h2a7;
        src104 <= 12'heda;
        src105 <= 12'h534;
        src106 <= 12'hceb;
        src107 <= 12'h6d2;
        src108 <= 12'h29e;
        src109 <= 12'hd39;
        src110 <= 12'ha8d;
        src111 <= 12'h6d;
        src112 <= 12'h1ee;
        src113 <= 12'h86c;
        src114 <= 12'h8fb;
        src115 <= 12'h53e;
        src116 <= 12'hb0b;
        src117 <= 12'h820;
        src118 <= 12'hb54;
        src119 <= 12'hf13;
        src120 <= 12'h1b4;
        src121 <= 12'h737;
        src122 <= 12'h126;
        src123 <= 12'h273;
        src124 <= 12'h311;
        src125 <= 12'h658;
        src126 <= 12'h82e;
        src127 <= 12'hee4;
        src128 <= 12'ha62;
        src129 <= 12'hf60;
        src130 <= 12'h52f;
        src131 <= 12'h396;
        src132 <= 12'h1e4;
        src133 <= 12'h678;
        src134 <= 12'h3ae;
        src135 <= 12'h2a3;
        src136 <= 12'h532;
        src137 <= 12'h1a3;
        src138 <= 12'h686;
        src139 <= 12'had8;
        src140 <= 12'h9fb;
        src141 <= 12'hb8e;
        src142 <= 12'hd47;
        src143 <= 12'h21c;
        src144 <= 12'h35e;
        src145 <= 12'hb89;
        src146 <= 12'h66d;
        src147 <= 12'he28;
        src148 <= 12'hff0;
        src149 <= 12'hb5;
        src150 <= 12'h427;
        src151 <= 12'hf82;
        src152 <= 12'h768;
        src153 <= 12'h6e6;
        src154 <= 12'hd2;
        src155 <= 12'h666;
        src156 <= 12'h670;
        src157 <= 12'hb68;
        src158 <= 12'hbf3;
        src159 <= 12'h148;
        src160 <= 12'h74a;
        src161 <= 12'he91;
        src162 <= 12'h4d0;
        src163 <= 12'hb37;
        src164 <= 12'h36;
        src165 <= 12'h433;
        src166 <= 12'h386;
        src167 <= 12'h805;
        src168 <= 12'h5b4;
        src169 <= 12'h93c;
        src170 <= 12'h512;
        src171 <= 12'h49e;
        src172 <= 12'hce3;
        src173 <= 12'hba1;
        src174 <= 12'h3e;
        src175 <= 12'h409;
        src176 <= 12'hb38;
        src177 <= 12'hb3b;
        src178 <= 12'hda6;
        src179 <= 12'hf49;
        src180 <= 12'h486;
        src181 <= 12'h4ea;
        src182 <= 12'ha42;
        src183 <= 12'h18c;
        src184 <= 12'h726;
        src185 <= 12'h434;
        src186 <= 12'hf3c;
        src187 <= 12'ha30;
        src188 <= 12'ha0b;
        exp <= 20'h5f35d;
        #1
        src0 <= 12'h4c7;
        src1 <= 12'h35b;
        src2 <= 12'h1fb;
        src3 <= 12'hfbe;
        src4 <= 12'h825;
        src5 <= 12'h606;
        src6 <= 12'hc5c;
        src7 <= 12'hf5b;
        src8 <= 12'hab9;
        src9 <= 12'h7f7;
        src10 <= 12'h6d6;
        src11 <= 12'h1e5;
        src12 <= 12'h18e;
        src13 <= 12'h9d2;
        src14 <= 12'hed1;
        src15 <= 12'hcab;
        src16 <= 12'h17c;
        src17 <= 12'hc6b;
        src18 <= 12'h315;
        src19 <= 12'hb42;
        src20 <= 12'hd1e;
        src21 <= 12'h719;
        src22 <= 12'h39f;
        src23 <= 12'ha2;
        src24 <= 12'hbfa;
        src25 <= 12'he81;
        src26 <= 12'heb2;
        src27 <= 12'h751;
        src28 <= 12'h3c3;
        src29 <= 12'hd76;
        src30 <= 12'h852;
        src31 <= 12'h8a4;
        src32 <= 12'h9c1;
        src33 <= 12'hb76;
        src34 <= 12'haba;
        src35 <= 12'hcfa;
        src36 <= 12'h6a9;
        src37 <= 12'h291;
        src38 <= 12'h3f5;
        src39 <= 12'h511;
        src40 <= 12'h961;
        src41 <= 12'h43c;
        src42 <= 12'ha83;
        src43 <= 12'heb7;
        src44 <= 12'h311;
        src45 <= 12'h9d8;
        src46 <= 12'hb8a;
        src47 <= 12'hc64;
        src48 <= 12'hdd2;
        src49 <= 12'hfde;
        src50 <= 12'h646;
        src51 <= 12'hdd5;
        src52 <= 12'h25b;
        src53 <= 12'h5ad;
        src54 <= 12'h526;
        src55 <= 12'hf9d;
        src56 <= 12'h3df;
        src57 <= 12'h1a5;
        src58 <= 12'h20f;
        src59 <= 12'hf38;
        src60 <= 12'h158;
        src61 <= 12'h683;
        src62 <= 12'h442;
        src63 <= 12'h606;
        src64 <= 12'hb4d;
        src65 <= 12'h7ea;
        src66 <= 12'hcde;
        src67 <= 12'hca7;
        src68 <= 12'h38;
        src69 <= 12'h74c;
        src70 <= 12'ha5b;
        src71 <= 12'hbea;
        src72 <= 12'heaf;
        src73 <= 12'he27;
        src74 <= 12'h7bb;
        src75 <= 12'hf4c;
        src76 <= 12'hef7;
        src77 <= 12'h96a;
        src78 <= 12'h15c;
        src79 <= 12'hb27;
        src80 <= 12'h254;
        src81 <= 12'h23d;
        src82 <= 12'ha2c;
        src83 <= 12'h271;
        src84 <= 12'h57f;
        src85 <= 12'hd05;
        src86 <= 12'h1d8;
        src87 <= 12'h3a8;
        src88 <= 12'hbdf;
        src89 <= 12'h428;
        src90 <= 12'h9cc;
        src91 <= 12'h2be;
        src92 <= 12'h7c0;
        src93 <= 12'hc54;
        src94 <= 12'h392;
        src95 <= 12'h690;
        src96 <= 12'h935;
        src97 <= 12'h3d9;
        src98 <= 12'h737;
        src99 <= 12'hf44;
        src100 <= 12'h9ec;
        src101 <= 12'he6f;
        src102 <= 12'h7;
        src103 <= 12'h5db;
        src104 <= 12'h475;
        src105 <= 12'hedf;
        src106 <= 12'h543;
        src107 <= 12'hed5;
        src108 <= 12'h93a;
        src109 <= 12'hd87;
        src110 <= 12'hba7;
        src111 <= 12'hf85;
        src112 <= 12'h2e8;
        src113 <= 12'hfa1;
        src114 <= 12'h3cf;
        src115 <= 12'hb8f;
        src116 <= 12'h39b;
        src117 <= 12'hf4e;
        src118 <= 12'hd91;
        src119 <= 12'hae;
        src120 <= 12'h493;
        src121 <= 12'h438;
        src122 <= 12'h4ed;
        src123 <= 12'hb7;
        src124 <= 12'h9b4;
        src125 <= 12'hf2e;
        src126 <= 12'hf58;
        src127 <= 12'hb31;
        src128 <= 12'h762;
        src129 <= 12'ha2e;
        src130 <= 12'h2b1;
        src131 <= 12'hb63;
        src132 <= 12'h50c;
        src133 <= 12'hc76;
        src134 <= 12'h817;
        src135 <= 12'hb8d;
        src136 <= 12'h69a;
        src137 <= 12'h4a8;
        src138 <= 12'ha58;
        src139 <= 12'h476;
        src140 <= 12'h477;
        src141 <= 12'h97;
        src142 <= 12'h3e0;
        src143 <= 12'ha7a;
        src144 <= 12'hb86;
        src145 <= 12'h148;
        src146 <= 12'hb2d;
        src147 <= 12'he6e;
        src148 <= 12'he15;
        src149 <= 12'h3f5;
        src150 <= 12'hc48;
        src151 <= 12'h602;
        src152 <= 12'hf08;
        src153 <= 12'h1b2;
        src154 <= 12'h51b;
        src155 <= 12'h10e;
        src156 <= 12'h769;
        src157 <= 12'he32;
        src158 <= 12'hcfa;
        src159 <= 12'h554;
        src160 <= 12'hfef;
        src161 <= 12'hb58;
        src162 <= 12'hdcc;
        src163 <= 12'h418;
        src164 <= 12'h5b4;
        src165 <= 12'h629;
        src166 <= 12'h602;
        src167 <= 12'h1eb;
        src168 <= 12'h5c3;
        src169 <= 12'h58a;
        src170 <= 12'h840;
        src171 <= 12'h4f4;
        src172 <= 12'h9f3;
        src173 <= 12'he1f;
        src174 <= 12'hc83;
        src175 <= 12'h98e;
        src176 <= 12'h9bc;
        src177 <= 12'hbd4;
        src178 <= 12'h8dc;
        src179 <= 12'h47f;
        src180 <= 12'hce0;
        src181 <= 12'h797;
        src182 <= 12'hef2;
        src183 <= 12'h586;
        src184 <= 12'h99e;
        src185 <= 12'had0;
        src186 <= 12'hec;
        src187 <= 12'h87;
        src188 <= 12'h92b;
        exp <= 20'h62555;
        #1
        src0 <= 12'h683;
        src1 <= 12'h992;
        src2 <= 12'hd62;
        src3 <= 12'h8a5;
        src4 <= 12'hd4e;
        src5 <= 12'hed2;
        src6 <= 12'hd08;
        src7 <= 12'hcd5;
        src8 <= 12'hb05;
        src9 <= 12'h82b;
        src10 <= 12'h338;
        src11 <= 12'hbe8;
        src12 <= 12'h754;
        src13 <= 12'h477;
        src14 <= 12'hfed;
        src15 <= 12'hf0f;
        src16 <= 12'h757;
        src17 <= 12'hebe;
        src18 <= 12'hfe4;
        src19 <= 12'h5cf;
        src20 <= 12'hf2d;
        src21 <= 12'hbad;
        src22 <= 12'haeb;
        src23 <= 12'h749;
        src24 <= 12'h617;
        src25 <= 12'h901;
        src26 <= 12'h99e;
        src27 <= 12'h7b8;
        src28 <= 12'h2;
        src29 <= 12'hd39;
        src30 <= 12'h482;
        src31 <= 12'h927;
        src32 <= 12'h71c;
        src33 <= 12'hfd0;
        src34 <= 12'h5a5;
        src35 <= 12'h365;
        src36 <= 12'h328;
        src37 <= 12'h279;
        src38 <= 12'ha48;
        src39 <= 12'h12;
        src40 <= 12'h9b4;
        src41 <= 12'haf5;
        src42 <= 12'hc06;
        src43 <= 12'h557;
        src44 <= 12'haae;
        src45 <= 12'h7b6;
        src46 <= 12'h27d;
        src47 <= 12'hae0;
        src48 <= 12'h4d4;
        src49 <= 12'h76e;
        src50 <= 12'h289;
        src51 <= 12'h2af;
        src52 <= 12'hb9;
        src53 <= 12'h7d1;
        src54 <= 12'hd91;
        src55 <= 12'h5ef;
        src56 <= 12'h977;
        src57 <= 12'h87f;
        src58 <= 12'h71b;
        src59 <= 12'h17b;
        src60 <= 12'hac6;
        src61 <= 12'h154;
        src62 <= 12'ha6d;
        src63 <= 12'h5c8;
        src64 <= 12'hcf;
        src65 <= 12'hec9;
        src66 <= 12'h309;
        src67 <= 12'hf65;
        src68 <= 12'h173;
        src69 <= 12'ha6f;
        src70 <= 12'h8b4;
        src71 <= 12'hda2;
        src72 <= 12'h814;
        src73 <= 12'hff4;
        src74 <= 12'h84a;
        src75 <= 12'hf4e;
        src76 <= 12'hb19;
        src77 <= 12'h17e;
        src78 <= 12'h125;
        src79 <= 12'h752;
        src80 <= 12'hcca;
        src81 <= 12'hefa;
        src82 <= 12'h576;
        src83 <= 12'hfa8;
        src84 <= 12'hf60;
        src85 <= 12'h7ad;
        src86 <= 12'h30f;
        src87 <= 12'h7ce;
        src88 <= 12'hf16;
        src89 <= 12'h609;
        src90 <= 12'h2a5;
        src91 <= 12'hb04;
        src92 <= 12'h765;
        src93 <= 12'h28f;
        src94 <= 12'h4fe;
        src95 <= 12'hcd5;
        src96 <= 12'h87b;
        src97 <= 12'h1ff;
        src98 <= 12'h560;
        src99 <= 12'ha50;
        src100 <= 12'h93e;
        src101 <= 12'h9b8;
        src102 <= 12'h524;
        src103 <= 12'hd00;
        src104 <= 12'hf36;
        src105 <= 12'hecd;
        src106 <= 12'h12c;
        src107 <= 12'ha4f;
        src108 <= 12'haf8;
        src109 <= 12'h492;
        src110 <= 12'h37d;
        src111 <= 12'h9a9;
        src112 <= 12'ha52;
        src113 <= 12'h1f5;
        src114 <= 12'hb3c;
        src115 <= 12'hac9;
        src116 <= 12'ha96;
        src117 <= 12'hf3d;
        src118 <= 12'h679;
        src119 <= 12'h189;
        src120 <= 12'hb8e;
        src121 <= 12'hd75;
        src122 <= 12'h610;
        src123 <= 12'ha2f;
        src124 <= 12'h951;
        src125 <= 12'ha13;
        src126 <= 12'h521;
        src127 <= 12'h6d8;
        src128 <= 12'h1;
        src129 <= 12'hb12;
        src130 <= 12'h533;
        src131 <= 12'h35f;
        src132 <= 12'h5c8;
        src133 <= 12'hd36;
        src134 <= 12'h1fa;
        src135 <= 12'h83d;
        src136 <= 12'h229;
        src137 <= 12'hd8b;
        src138 <= 12'h3b5;
        src139 <= 12'h82;
        src140 <= 12'hbf2;
        src141 <= 12'h872;
        src142 <= 12'hf17;
        src143 <= 12'h60;
        src144 <= 12'hf4b;
        src145 <= 12'h966;
        src146 <= 12'h72;
        src147 <= 12'h1cb;
        src148 <= 12'haeb;
        src149 <= 12'h3a5;
        src150 <= 12'he0b;
        src151 <= 12'h7c4;
        src152 <= 12'h8a2;
        src153 <= 12'h3c4;
        src154 <= 12'hcf6;
        src155 <= 12'h5e7;
        src156 <= 12'h95;
        src157 <= 12'h8fe;
        src158 <= 12'hdad;
        src159 <= 12'h518;
        src160 <= 12'hca1;
        src161 <= 12'h824;
        src162 <= 12'hdcf;
        src163 <= 12'h488;
        src164 <= 12'h5d7;
        src165 <= 12'h421;
        src166 <= 12'h194;
        src167 <= 12'hefd;
        src168 <= 12'hc58;
        src169 <= 12'h487;
        src170 <= 12'h6dc;
        src171 <= 12'hcb6;
        src172 <= 12'hce7;
        src173 <= 12'h27d;
        src174 <= 12'ha0e;
        src175 <= 12'he4d;
        src176 <= 12'h378;
        src177 <= 12'h4f5;
        src178 <= 12'h392;
        src179 <= 12'hdff;
        src180 <= 12'h38e;
        src181 <= 12'hb6a;
        src182 <= 12'hd4b;
        src183 <= 12'h1d5;
        src184 <= 12'hb29;
        src185 <= 12'hb2;
        src186 <= 12'hec3;
        src187 <= 12'h79f;
        src188 <= 12'h138;
        exp <= 20'h610d0;
        #1
        src0 <= 12'h500;
        src1 <= 12'he27;
        src2 <= 12'h997;
        src3 <= 12'h3da;
        src4 <= 12'h106;
        src5 <= 12'h48d;
        src6 <= 12'h8bb;
        src7 <= 12'hedf;
        src8 <= 12'h76e;
        src9 <= 12'hd78;
        src10 <= 12'hffa;
        src11 <= 12'ha1e;
        src12 <= 12'he7b;
        src13 <= 12'hbd8;
        src14 <= 12'h98c;
        src15 <= 12'hc3d;
        src16 <= 12'hbb3;
        src17 <= 12'h49;
        src18 <= 12'h857;
        src19 <= 12'hf87;
        src20 <= 12'hfb7;
        src21 <= 12'h391;
        src22 <= 12'h7a6;
        src23 <= 12'hd7;
        src24 <= 12'he65;
        src25 <= 12'h4be;
        src26 <= 12'hebd;
        src27 <= 12'hedb;
        src28 <= 12'hcf9;
        src29 <= 12'h924;
        src30 <= 12'h1e1;
        src31 <= 12'hb0;
        src32 <= 12'h513;
        src33 <= 12'ha20;
        src34 <= 12'habd;
        src35 <= 12'hd62;
        src36 <= 12'hc93;
        src37 <= 12'h5d1;
        src38 <= 12'h909;
        src39 <= 12'h257;
        src40 <= 12'ha38;
        src41 <= 12'hbc2;
        src42 <= 12'hcfc;
        src43 <= 12'hd3d;
        src44 <= 12'h6bb;
        src45 <= 12'he24;
        src46 <= 12'h659;
        src47 <= 12'h97a;
        src48 <= 12'h958;
        src49 <= 12'h77;
        src50 <= 12'h719;
        src51 <= 12'h8ae;
        src52 <= 12'h50d;
        src53 <= 12'hd0d;
        src54 <= 12'hb8;
        src55 <= 12'hacb;
        src56 <= 12'h651;
        src57 <= 12'h8a2;
        src58 <= 12'ha91;
        src59 <= 12'hbbb;
        src60 <= 12'hde5;
        src61 <= 12'hbed;
        src62 <= 12'hcf0;
        src63 <= 12'hdab;
        src64 <= 12'hde3;
        src65 <= 12'h235;
        src66 <= 12'hb0b;
        src67 <= 12'haee;
        src68 <= 12'h71a;
        src69 <= 12'h526;
        src70 <= 12'hba;
        src71 <= 12'h465;
        src72 <= 12'hdd7;
        src73 <= 12'he69;
        src74 <= 12'h62;
        src75 <= 12'ha8c;
        src76 <= 12'h132;
        src77 <= 12'h5c0;
        src78 <= 12'h563;
        src79 <= 12'hc05;
        src80 <= 12'h294;
        src81 <= 12'h439;
        src82 <= 12'h930;
        src83 <= 12'hb7d;
        src84 <= 12'h2fc;
        src85 <= 12'h4d3;
        src86 <= 12'hc0;
        src87 <= 12'hde0;
        src88 <= 12'h868;
        src89 <= 12'h580;
        src90 <= 12'h7ac;
        src91 <= 12'h3a6;
        src92 <= 12'h681;
        src93 <= 12'h733;
        src94 <= 12'hf84;
        src95 <= 12'hf40;
        src96 <= 12'h681;
        src97 <= 12'h44b;
        src98 <= 12'hbe1;
        src99 <= 12'hb32;
        src100 <= 12'h9ae;
        src101 <= 12'ha3;
        src102 <= 12'hb2c;
        src103 <= 12'h19d;
        src104 <= 12'h943;
        src105 <= 12'h288;
        src106 <= 12'h3f4;
        src107 <= 12'hb79;
        src108 <= 12'haad;
        src109 <= 12'h577;
        src110 <= 12'hd46;
        src111 <= 12'h2ca;
        src112 <= 12'hfd6;
        src113 <= 12'hd03;
        src114 <= 12'hcf0;
        src115 <= 12'h7f1;
        src116 <= 12'h9f1;
        src117 <= 12'hda0;
        src118 <= 12'h418;
        src119 <= 12'h589;
        src120 <= 12'h60e;
        src121 <= 12'hb1f;
        src122 <= 12'h615;
        src123 <= 12'ha;
        src124 <= 12'h7e4;
        src125 <= 12'h6a;
        src126 <= 12'h400;
        src127 <= 12'h13e;
        src128 <= 12'hf0a;
        src129 <= 12'hb85;
        src130 <= 12'h98b;
        src131 <= 12'h306;
        src132 <= 12'hcb1;
        src133 <= 12'h4f9;
        src134 <= 12'hd08;
        src135 <= 12'h6bd;
        src136 <= 12'h58c;
        src137 <= 12'hcae;
        src138 <= 12'h294;
        src139 <= 12'h5b1;
        src140 <= 12'hcf8;
        src141 <= 12'h4df;
        src142 <= 12'h1ee;
        src143 <= 12'h7e;
        src144 <= 12'hc7;
        src145 <= 12'hbe9;
        src146 <= 12'h2f4;
        src147 <= 12'ha94;
        src148 <= 12'h3d9;
        src149 <= 12'h829;
        src150 <= 12'h7ae;
        src151 <= 12'hc96;
        src152 <= 12'hdcb;
        src153 <= 12'haff;
        src154 <= 12'hbb7;
        src155 <= 12'h97d;
        src156 <= 12'h3fb;
        src157 <= 12'he76;
        src158 <= 12'h281;
        src159 <= 12'ha74;
        src160 <= 12'h8b6;
        src161 <= 12'h53e;
        src162 <= 12'h408;
        src163 <= 12'hfd0;
        src164 <= 12'hce5;
        src165 <= 12'hd69;
        src166 <= 12'h5d3;
        src167 <= 12'h12f;
        src168 <= 12'h3e8;
        src169 <= 12'hf6c;
        src170 <= 12'hac3;
        src171 <= 12'hd6e;
        src172 <= 12'h6fc;
        src173 <= 12'h84c;
        src174 <= 12'hdf9;
        src175 <= 12'h451;
        src176 <= 12'hc13;
        src177 <= 12'h2d5;
        src178 <= 12'h7ff;
        src179 <= 12'h2df;
        src180 <= 12'h5b9;
        src181 <= 12'h129;
        src182 <= 12'h971;
        src183 <= 12'h612;
        src184 <= 12'h18b;
        src185 <= 12'h915;
        src186 <= 12'h820;
        src187 <= 12'hb63;
        src188 <= 12'h414;
        exp <= 20'h61145;
        #1
        src0 <= 12'h49c;
        src1 <= 12'h20;
        src2 <= 12'h209;
        src3 <= 12'h9d1;
        src4 <= 12'h295;
        src5 <= 12'h87b;
        src6 <= 12'h1a;
        src7 <= 12'h58c;
        src8 <= 12'hfbf;
        src9 <= 12'hb54;
        src10 <= 12'h562;
        src11 <= 12'h3d5;
        src12 <= 12'hd00;
        src13 <= 12'hcd7;
        src14 <= 12'ha71;
        src15 <= 12'h46d;
        src16 <= 12'h440;
        src17 <= 12'h146;
        src18 <= 12'h598;
        src19 <= 12'h928;
        src20 <= 12'hf89;
        src21 <= 12'h2;
        src22 <= 12'hf86;
        src23 <= 12'h6f9;
        src24 <= 12'h79f;
        src25 <= 12'hafe;
        src26 <= 12'h2ab;
        src27 <= 12'h5b;
        src28 <= 12'h32;
        src29 <= 12'ha33;
        src30 <= 12'hdef;
        src31 <= 12'h4c0;
        src32 <= 12'h427;
        src33 <= 12'hc26;
        src34 <= 12'h983;
        src35 <= 12'h1c2;
        src36 <= 12'h286;
        src37 <= 12'hab2;
        src38 <= 12'h4fd;
        src39 <= 12'h3f6;
        src40 <= 12'hf17;
        src41 <= 12'hbc4;
        src42 <= 12'h601;
        src43 <= 12'ha0e;
        src44 <= 12'h3e7;
        src45 <= 12'h2b0;
        src46 <= 12'hb4a;
        src47 <= 12'h9dc;
        src48 <= 12'hbec;
        src49 <= 12'h115;
        src50 <= 12'hff8;
        src51 <= 12'h22;
        src52 <= 12'h598;
        src53 <= 12'h22;
        src54 <= 12'h81f;
        src55 <= 12'h4da;
        src56 <= 12'h993;
        src57 <= 12'h801;
        src58 <= 12'he01;
        src59 <= 12'h330;
        src60 <= 12'h383;
        src61 <= 12'h122;
        src62 <= 12'h231;
        src63 <= 12'h33f;
        src64 <= 12'h622;
        src65 <= 12'h236;
        src66 <= 12'hb04;
        src67 <= 12'h887;
        src68 <= 12'h3fb;
        src69 <= 12'h25d;
        src70 <= 12'h829;
        src71 <= 12'hd8b;
        src72 <= 12'hd9f;
        src73 <= 12'h5ac;
        src74 <= 12'hbdc;
        src75 <= 12'hd64;
        src76 <= 12'h80;
        src77 <= 12'h2ac;
        src78 <= 12'h534;
        src79 <= 12'hc2f;
        src80 <= 12'heb7;
        src81 <= 12'h2c;
        src82 <= 12'hb3d;
        src83 <= 12'h189;
        src84 <= 12'h9c1;
        src85 <= 12'h3a3;
        src86 <= 12'hca5;
        src87 <= 12'hf1d;
        src88 <= 12'hf5b;
        src89 <= 12'h3da;
        src90 <= 12'h651;
        src91 <= 12'h591;
        src92 <= 12'hea9;
        src93 <= 12'hb2d;
        src94 <= 12'h948;
        src95 <= 12'h2e2;
        src96 <= 12'h8e3;
        src97 <= 12'ha2a;
        src98 <= 12'hb23;
        src99 <= 12'h366;
        src100 <= 12'hed4;
        src101 <= 12'h958;
        src102 <= 12'h46e;
        src103 <= 12'h83a;
        src104 <= 12'h875;
        src105 <= 12'h81d;
        src106 <= 12'hcf1;
        src107 <= 12'hee3;
        src108 <= 12'hccd;
        src109 <= 12'haaf;
        src110 <= 12'h6b4;
        src111 <= 12'h113;
        src112 <= 12'h51a;
        src113 <= 12'h1d0;
        src114 <= 12'h721;
        src115 <= 12'h17a;
        src116 <= 12'ha57;
        src117 <= 12'hae;
        src118 <= 12'h13c;
        src119 <= 12'he31;
        src120 <= 12'h373;
        src121 <= 12'h599;
        src122 <= 12'h858;
        src123 <= 12'hd6b;
        src124 <= 12'hb35;
        src125 <= 12'hc66;
        src126 <= 12'h1c2;
        src127 <= 12'h3d8;
        src128 <= 12'hf97;
        src129 <= 12'he07;
        src130 <= 12'hc44;
        src131 <= 12'hc26;
        src132 <= 12'hd80;
        src133 <= 12'hd8f;
        src134 <= 12'h93b;
        src135 <= 12'h8e9;
        src136 <= 12'h683;
        src137 <= 12'h4a8;
        src138 <= 12'h71f;
        src139 <= 12'h624;
        src140 <= 12'hde5;
        src141 <= 12'hfc1;
        src142 <= 12'h76e;
        src143 <= 12'h356;
        src144 <= 12'hfcd;
        src145 <= 12'h29f;
        src146 <= 12'hb;
        src147 <= 12'hcfe;
        src148 <= 12'he37;
        src149 <= 12'hc26;
        src150 <= 12'hbf2;
        src151 <= 12'h508;
        src152 <= 12'h977;
        src153 <= 12'hf56;
        src154 <= 12'h7b7;
        src155 <= 12'h443;
        src156 <= 12'hed6;
        src157 <= 12'h224;
        src158 <= 12'h770;
        src159 <= 12'h811;
        src160 <= 12'h65b;
        src161 <= 12'hf6d;
        src162 <= 12'h9b2;
        src163 <= 12'h7a1;
        src164 <= 12'h715;
        src165 <= 12'h30d;
        src166 <= 12'h50b;
        src167 <= 12'h2d6;
        src168 <= 12'hdc9;
        src169 <= 12'hd4b;
        src170 <= 12'h159;
        src171 <= 12'h170;
        src172 <= 12'hddc;
        src173 <= 12'h3da;
        src174 <= 12'hfd9;
        src175 <= 12'h48e;
        src176 <= 12'h92a;
        src177 <= 12'he26;
        src178 <= 12'hfd4;
        src179 <= 12'h741;
        src180 <= 12'hb12;
        src181 <= 12'h626;
        src182 <= 12'h911;
        src183 <= 12'h816;
        src184 <= 12'h6c8;
        src185 <= 12'h7c4;
        src186 <= 12'h376;
        src187 <= 12'h761;
        src188 <= 12'h9c7;
        exp <= 20'h5d082;
        #1
        src0 <= 12'h885;
        src1 <= 12'ha55;
        src2 <= 12'h286;
        src3 <= 12'h5d8;
        src4 <= 12'hff6;
        src5 <= 12'hb45;
        src6 <= 12'hcb6;
        src7 <= 12'hce2;
        src8 <= 12'h567;
        src9 <= 12'hf05;
        src10 <= 12'h890;
        src11 <= 12'heec;
        src12 <= 12'h2f3;
        src13 <= 12'h7f4;
        src14 <= 12'h510;
        src15 <= 12'h4a3;
        src16 <= 12'hc0d;
        src17 <= 12'hdd9;
        src18 <= 12'h52a;
        src19 <= 12'h14a;
        src20 <= 12'he9e;
        src21 <= 12'hd84;
        src22 <= 12'h268;
        src23 <= 12'hdd;
        src24 <= 12'h99c;
        src25 <= 12'h717;
        src26 <= 12'hc0f;
        src27 <= 12'h7d3;
        src28 <= 12'h2a3;
        src29 <= 12'hc5d;
        src30 <= 12'h28c;
        src31 <= 12'heee;
        src32 <= 12'h775;
        src33 <= 12'h31f;
        src34 <= 12'h8e2;
        src35 <= 12'h5dc;
        src36 <= 12'hcb9;
        src37 <= 12'h574;
        src38 <= 12'hcb5;
        src39 <= 12'h798;
        src40 <= 12'hce6;
        src41 <= 12'h94e;
        src42 <= 12'hbbd;
        src43 <= 12'h36e;
        src44 <= 12'hf2e;
        src45 <= 12'h21f;
        src46 <= 12'h679;
        src47 <= 12'hef1;
        src48 <= 12'had7;
        src49 <= 12'h92c;
        src50 <= 12'hde8;
        src51 <= 12'h770;
        src52 <= 12'ha9a;
        src53 <= 12'h754;
        src54 <= 12'heb;
        src55 <= 12'h14b;
        src56 <= 12'h136;
        src57 <= 12'hc61;
        src58 <= 12'hde8;
        src59 <= 12'h684;
        src60 <= 12'h323;
        src61 <= 12'hc75;
        src62 <= 12'h265;
        src63 <= 12'hb97;
        src64 <= 12'hc3f;
        src65 <= 12'ha2;
        src66 <= 12'h7e4;
        src67 <= 12'h6ad;
        src68 <= 12'h4ea;
        src69 <= 12'h7c4;
        src70 <= 12'h263;
        src71 <= 12'h971;
        src72 <= 12'h9b1;
        src73 <= 12'hafb;
        src74 <= 12'h589;
        src75 <= 12'h5fb;
        src76 <= 12'h9aa;
        src77 <= 12'h84a;
        src78 <= 12'hce1;
        src79 <= 12'h8;
        src80 <= 12'hcc8;
        src81 <= 12'h470;
        src82 <= 12'h43a;
        src83 <= 12'h9c5;
        src84 <= 12'h3b4;
        src85 <= 12'h264;
        src86 <= 12'he9d;
        src87 <= 12'ha4a;
        src88 <= 12'h44f;
        src89 <= 12'h74d;
        src90 <= 12'h59e;
        src91 <= 12'h46d;
        src92 <= 12'he08;
        src93 <= 12'ha80;
        src94 <= 12'h20b;
        src95 <= 12'h8e3;
        src96 <= 12'h2e7;
        src97 <= 12'h566;
        src98 <= 12'hfee;
        src99 <= 12'h12f;
        src100 <= 12'h90a;
        src101 <= 12'h20b;
        src102 <= 12'h3da;
        src103 <= 12'h362;
        src104 <= 12'h9f5;
        src105 <= 12'h148;
        src106 <= 12'h384;
        src107 <= 12'h9a7;
        src108 <= 12'hc4d;
        src109 <= 12'h669;
        src110 <= 12'hd6;
        src111 <= 12'h23c;
        src112 <= 12'h3ea;
        src113 <= 12'h424;
        src114 <= 12'h5b8;
        src115 <= 12'h73c;
        src116 <= 12'h717;
        src117 <= 12'he0;
        src118 <= 12'h8cd;
        src119 <= 12'hc8c;
        src120 <= 12'he08;
        src121 <= 12'hffb;
        src122 <= 12'hdfe;
        src123 <= 12'he77;
        src124 <= 12'hc90;
        src125 <= 12'hc69;
        src126 <= 12'h48c;
        src127 <= 12'h6e1;
        src128 <= 12'hf90;
        src129 <= 12'he48;
        src130 <= 12'hba5;
        src131 <= 12'hb8e;
        src132 <= 12'h7e9;
        src133 <= 12'hfb7;
        src134 <= 12'hd65;
        src135 <= 12'hc80;
        src136 <= 12'h370;
        src137 <= 12'hdd4;
        src138 <= 12'h1ab;
        src139 <= 12'h804;
        src140 <= 12'h96a;
        src141 <= 12'h8a2;
        src142 <= 12'h26e;
        src143 <= 12'h33b;
        src144 <= 12'hc07;
        src145 <= 12'h7f3;
        src146 <= 12'hf9c;
        src147 <= 12'ha2e;
        src148 <= 12'hed4;
        src149 <= 12'h147;
        src150 <= 12'h544;
        src151 <= 12'h66e;
        src152 <= 12'hc90;
        src153 <= 12'h1a;
        src154 <= 12'h3e8;
        src155 <= 12'h51;
        src156 <= 12'hc92;
        src157 <= 12'hf8;
        src158 <= 12'hc77;
        src159 <= 12'h658;
        src160 <= 12'h13b;
        src161 <= 12'hebd;
        src162 <= 12'hd9c;
        src163 <= 12'hb2;
        src164 <= 12'h930;
        src165 <= 12'he89;
        src166 <= 12'hbf6;
        src167 <= 12'h99e;
        src168 <= 12'h897;
        src169 <= 12'h3b9;
        src170 <= 12'h2f6;
        src171 <= 12'he9c;
        src172 <= 12'h8a1;
        src173 <= 12'hed8;
        src174 <= 12'h2b2;
        src175 <= 12'h9c;
        src176 <= 12'ha1d;
        src177 <= 12'hff7;
        src178 <= 12'hf81;
        src179 <= 12'h4ac;
        src180 <= 12'hdcb;
        src181 <= 12'h225;
        src182 <= 12'hcc1;
        src183 <= 12'hf05;
        src184 <= 12'hf47;
        src185 <= 12'hcdf;
        src186 <= 12'h11c;
        src187 <= 12'h16e;
        src188 <= 12'he06;
        exp <= 20'h612b2;
        #1
        src0 <= 12'h6e7;
        src1 <= 12'hfba;
        src2 <= 12'h4db;
        src3 <= 12'h5e;
        src4 <= 12'hf46;
        src5 <= 12'he1d;
        src6 <= 12'h90b;
        src7 <= 12'he9e;
        src8 <= 12'ha5c;
        src9 <= 12'he38;
        src10 <= 12'h60c;
        src11 <= 12'hf51;
        src12 <= 12'h3d1;
        src13 <= 12'he43;
        src14 <= 12'h566;
        src15 <= 12'h6be;
        src16 <= 12'h8b6;
        src17 <= 12'h67a;
        src18 <= 12'h985;
        src19 <= 12'h62a;
        src20 <= 12'h980;
        src21 <= 12'hd96;
        src22 <= 12'hf48;
        src23 <= 12'h715;
        src24 <= 12'hb9e;
        src25 <= 12'h133;
        src26 <= 12'h6c8;
        src27 <= 12'heaa;
        src28 <= 12'h70c;
        src29 <= 12'h4ed;
        src30 <= 12'hc69;
        src31 <= 12'hdce;
        src32 <= 12'h35d;
        src33 <= 12'h2c1;
        src34 <= 12'h77a;
        src35 <= 12'h8ae;
        src36 <= 12'h869;
        src37 <= 12'ha20;
        src38 <= 12'hf48;
        src39 <= 12'h1d4;
        src40 <= 12'h98;
        src41 <= 12'he12;
        src42 <= 12'h616;
        src43 <= 12'h3e6;
        src44 <= 12'h44b;
        src45 <= 12'h5f1;
        src46 <= 12'hb7a;
        src47 <= 12'hdee;
        src48 <= 12'hd8d;
        src49 <= 12'hacc;
        src50 <= 12'h445;
        src51 <= 12'hed3;
        src52 <= 12'h277;
        src53 <= 12'h2ad;
        src54 <= 12'hb10;
        src55 <= 12'h285;
        src56 <= 12'h715;
        src57 <= 12'h13;
        src58 <= 12'h8b8;
        src59 <= 12'h42a;
        src60 <= 12'h38;
        src61 <= 12'he23;
        src62 <= 12'h40c;
        src63 <= 12'h860;
        src64 <= 12'hd80;
        src65 <= 12'hd1d;
        src66 <= 12'h100;
        src67 <= 12'h97;
        src68 <= 12'hb1a;
        src69 <= 12'h1eb;
        src70 <= 12'hfd5;
        src71 <= 12'h88f;
        src72 <= 12'h187;
        src73 <= 12'h424;
        src74 <= 12'hbee;
        src75 <= 12'h47b;
        src76 <= 12'h3f9;
        src77 <= 12'h26e;
        src78 <= 12'h956;
        src79 <= 12'hddf;
        src80 <= 12'h4c3;
        src81 <= 12'h7d5;
        src82 <= 12'habe;
        src83 <= 12'h32;
        src84 <= 12'he80;
        src85 <= 12'hfd4;
        src86 <= 12'hee6;
        src87 <= 12'h654;
        src88 <= 12'h6f1;
        src89 <= 12'h5b3;
        src90 <= 12'h7e8;
        src91 <= 12'h77;
        src92 <= 12'h2a2;
        src93 <= 12'h357;
        src94 <= 12'he6b;
        src95 <= 12'hd83;
        src96 <= 12'hfd7;
        src97 <= 12'h47b;
        src98 <= 12'h6a3;
        src99 <= 12'hb3;
        src100 <= 12'h12d;
        src101 <= 12'h60e;
        src102 <= 12'h38c;
        src103 <= 12'h6b4;
        src104 <= 12'haa1;
        src105 <= 12'ha01;
        src106 <= 12'h6a3;
        src107 <= 12'hfe0;
        src108 <= 12'hce1;
        src109 <= 12'h417;
        src110 <= 12'h787;
        src111 <= 12'h80b;
        src112 <= 12'h23f;
        src113 <= 12'hd0d;
        src114 <= 12'h39f;
        src115 <= 12'hc2;
        src116 <= 12'h338;
        src117 <= 12'hec0;
        src118 <= 12'h9bc;
        src119 <= 12'hcb7;
        src120 <= 12'h909;
        src121 <= 12'h208;
        src122 <= 12'h42b;
        src123 <= 12'hf0e;
        src124 <= 12'hfba;
        src125 <= 12'h8f7;
        src126 <= 12'hdfc;
        src127 <= 12'hd6e;
        src128 <= 12'heb9;
        src129 <= 12'h4a9;
        src130 <= 12'h948;
        src131 <= 12'h511;
        src132 <= 12'h52f;
        src133 <= 12'h4a2;
        src134 <= 12'h611;
        src135 <= 12'haba;
        src136 <= 12'h6a0;
        src137 <= 12'h70b;
        src138 <= 12'hc1a;
        src139 <= 12'hc36;
        src140 <= 12'hd2;
        src141 <= 12'h9df;
        src142 <= 12'hf00;
        src143 <= 12'h64a;
        src144 <= 12'h3fc;
        src145 <= 12'hb24;
        src146 <= 12'h84b;
        src147 <= 12'hc3f;
        src148 <= 12'h33f;
        src149 <= 12'h281;
        src150 <= 12'h2eb;
        src151 <= 12'h646;
        src152 <= 12'hacd;
        src153 <= 12'h739;
        src154 <= 12'h660;
        src155 <= 12'hfee;
        src156 <= 12'he90;
        src157 <= 12'h68a;
        src158 <= 12'hd88;
        src159 <= 12'h7f3;
        src160 <= 12'h174;
        src161 <= 12'h24e;
        src162 <= 12'h637;
        src163 <= 12'h5e3;
        src164 <= 12'h85a;
        src165 <= 12'hf4b;
        src166 <= 12'hcc5;
        src167 <= 12'h191;
        src168 <= 12'h123;
        src169 <= 12'hf63;
        src170 <= 12'hfce;
        src171 <= 12'h7c5;
        src172 <= 12'h8c3;
        src173 <= 12'h5da;
        src174 <= 12'hc0;
        src175 <= 12'heb6;
        src176 <= 12'h331;
        src177 <= 12'h636;
        src178 <= 12'h283;
        src179 <= 12'h362;
        src180 <= 12'he09;
        src181 <= 12'h538;
        src182 <= 12'h205;
        src183 <= 12'h4e5;
        src184 <= 12'h18f;
        src185 <= 12'hf25;
        src186 <= 12'h3ce;
        src187 <= 12'h2e1;
        src188 <= 12'hf7a;
        exp <= 20'h5e7c8;
        #1
        src0 <= 12'h1f3;
        src1 <= 12'hfd4;
        src2 <= 12'ha2;
        src3 <= 12'h509;
        src4 <= 12'h607;
        src5 <= 12'hee;
        src6 <= 12'h9e5;
        src7 <= 12'hf96;
        src8 <= 12'h426;
        src9 <= 12'h438;
        src10 <= 12'h904;
        src11 <= 12'hd66;
        src12 <= 12'h253;
        src13 <= 12'h42d;
        src14 <= 12'h8a7;
        src15 <= 12'hf11;
        src16 <= 12'he11;
        src17 <= 12'hcdc;
        src18 <= 12'hd84;
        src19 <= 12'heca;
        src20 <= 12'h905;
        src21 <= 12'hb25;
        src22 <= 12'hb00;
        src23 <= 12'h73e;
        src24 <= 12'h429;
        src25 <= 12'hd54;
        src26 <= 12'h8f;
        src27 <= 12'h655;
        src28 <= 12'h90b;
        src29 <= 12'hdff;
        src30 <= 12'hc1a;
        src31 <= 12'h72d;
        src32 <= 12'hc7f;
        src33 <= 12'h9d2;
        src34 <= 12'h485;
        src35 <= 12'h61b;
        src36 <= 12'he46;
        src37 <= 12'h3db;
        src38 <= 12'h7c1;
        src39 <= 12'h287;
        src40 <= 12'h59;
        src41 <= 12'h23e;
        src42 <= 12'h9db;
        src43 <= 12'hc17;
        src44 <= 12'h25d;
        src45 <= 12'hb57;
        src46 <= 12'h9fb;
        src47 <= 12'h608;
        src48 <= 12'hf3c;
        src49 <= 12'h5db;
        src50 <= 12'hcb0;
        src51 <= 12'he3b;
        src52 <= 12'ha6a;
        src53 <= 12'h1fd;
        src54 <= 12'h6f2;
        src55 <= 12'h6d7;
        src56 <= 12'he11;
        src57 <= 12'hbe6;
        src58 <= 12'hfdc;
        src59 <= 12'h42f;
        src60 <= 12'hca8;
        src61 <= 12'hca8;
        src62 <= 12'h2f;
        src63 <= 12'h562;
        src64 <= 12'h92d;
        src65 <= 12'hd15;
        src66 <= 12'ha41;
        src67 <= 12'hdd3;
        src68 <= 12'h1ac;
        src69 <= 12'hd2c;
        src70 <= 12'h68d;
        src71 <= 12'hb20;
        src72 <= 12'hcd3;
        src73 <= 12'h2a7;
        src74 <= 12'h5b1;
        src75 <= 12'h390;
        src76 <= 12'hfa2;
        src77 <= 12'ha27;
        src78 <= 12'hfc2;
        src79 <= 12'h851;
        src80 <= 12'hacf;
        src81 <= 12'h888;
        src82 <= 12'h1c3;
        src83 <= 12'h286;
        src84 <= 12'h34;
        src85 <= 12'hb8f;
        src86 <= 12'h6f2;
        src87 <= 12'h9e6;
        src88 <= 12'hbb9;
        src89 <= 12'hb31;
        src90 <= 12'h1a8;
        src91 <= 12'hf9c;
        src92 <= 12'h5d0;
        src93 <= 12'hf50;
        src94 <= 12'hc9e;
        src95 <= 12'hdb;
        src96 <= 12'hbf2;
        src97 <= 12'hb4b;
        src98 <= 12'h195;
        src99 <= 12'hf0f;
        src100 <= 12'h21;
        src101 <= 12'h128;
        src102 <= 12'hd13;
        src103 <= 12'hbd6;
        src104 <= 12'h3f1;
        src105 <= 12'h4c9;
        src106 <= 12'h92b;
        src107 <= 12'h8f;
        src108 <= 12'hf4d;
        src109 <= 12'h354;
        src110 <= 12'h3a6;
        src111 <= 12'h57e;
        src112 <= 12'heed;
        src113 <= 12'hf13;
        src114 <= 12'h542;
        src115 <= 12'hc8c;
        src116 <= 12'hc05;
        src117 <= 12'hf6;
        src118 <= 12'h366;
        src119 <= 12'h38;
        src120 <= 12'h89a;
        src121 <= 12'hbb4;
        src122 <= 12'h521;
        src123 <= 12'h841;
        src124 <= 12'ha37;
        src125 <= 12'h919;
        src126 <= 12'h6b1;
        src127 <= 12'h31d;
        src128 <= 12'h15a;
        src129 <= 12'hb0;
        src130 <= 12'hc32;
        src131 <= 12'h17;
        src132 <= 12'h25c;
        src133 <= 12'h5d8;
        src134 <= 12'h7fe;
        src135 <= 12'ha10;
        src136 <= 12'h2eb;
        src137 <= 12'hd46;
        src138 <= 12'hfb8;
        src139 <= 12'h7f1;
        src140 <= 12'h8e3;
        src141 <= 12'h830;
        src142 <= 12'h843;
        src143 <= 12'h98b;
        src144 <= 12'h54c;
        src145 <= 12'h34;
        src146 <= 12'h530;
        src147 <= 12'hce;
        src148 <= 12'hd47;
        src149 <= 12'h38b;
        src150 <= 12'hd63;
        src151 <= 12'h5e7;
        src152 <= 12'h1ad;
        src153 <= 12'hbc4;
        src154 <= 12'h3ca;
        src155 <= 12'h8c7;
        src156 <= 12'ha09;
        src157 <= 12'h596;
        src158 <= 12'hff3;
        src159 <= 12'h1d5;
        src160 <= 12'haf8;
        src161 <= 12'h95b;
        src162 <= 12'h943;
        src163 <= 12'hcc0;
        src164 <= 12'hd76;
        src165 <= 12'hea1;
        src166 <= 12'h2b;
        src167 <= 12'hd79;
        src168 <= 12'hed1;
        src169 <= 12'hf98;
        src170 <= 12'hb4;
        src171 <= 12'hb04;
        src172 <= 12'h174;
        src173 <= 12'hbcc;
        src174 <= 12'hc07;
        src175 <= 12'h16a;
        src176 <= 12'hb46;
        src177 <= 12'h613;
        src178 <= 12'hbf5;
        src179 <= 12'ha30;
        src180 <= 12'hce0;
        src181 <= 12'hf6b;
        src182 <= 12'h6f;
        src183 <= 12'h29b;
        src184 <= 12'he04;
        src185 <= 12'h33f;
        src186 <= 12'h28;
        src187 <= 12'h902;
        src188 <= 12'h8fe;
        exp <= 20'h6094f;
        #1
        src0 <= 12'h436;
        src1 <= 12'h7d4;
        src2 <= 12'h113;
        src3 <= 12'h4b5;
        src4 <= 12'h26c;
        src5 <= 12'hdcd;
        src6 <= 12'h2dc;
        src7 <= 12'h387;
        src8 <= 12'h5d7;
        src9 <= 12'h6c1;
        src10 <= 12'ha0f;
        src11 <= 12'h790;
        src12 <= 12'h32b;
        src13 <= 12'hb79;
        src14 <= 12'ha02;
        src15 <= 12'h4b0;
        src16 <= 12'h314;
        src17 <= 12'h7c9;
        src18 <= 12'h34a;
        src19 <= 12'h39b;
        src20 <= 12'h5a7;
        src21 <= 12'h6f2;
        src22 <= 12'h223;
        src23 <= 12'hd9a;
        src24 <= 12'h76d;
        src25 <= 12'h61f;
        src26 <= 12'h854;
        src27 <= 12'hda5;
        src28 <= 12'hc7f;
        src29 <= 12'h33;
        src30 <= 12'h72;
        src31 <= 12'he58;
        src32 <= 12'h513;
        src33 <= 12'hca9;
        src34 <= 12'h54e;
        src35 <= 12'hc3b;
        src36 <= 12'h81;
        src37 <= 12'h18e;
        src38 <= 12'h8ef;
        src39 <= 12'h1fb;
        src40 <= 12'h9b7;
        src41 <= 12'ha9d;
        src42 <= 12'h4bb;
        src43 <= 12'h6a5;
        src44 <= 12'h881;
        src45 <= 12'hdaa;
        src46 <= 12'h372;
        src47 <= 12'ha9f;
        src48 <= 12'hb35;
        src49 <= 12'h195;
        src50 <= 12'hdac;
        src51 <= 12'hfc3;
        src52 <= 12'h723;
        src53 <= 12'hd01;
        src54 <= 12'h5f6;
        src55 <= 12'hd58;
        src56 <= 12'h4cf;
        src57 <= 12'h689;
        src58 <= 12'h769;
        src59 <= 12'ha85;
        src60 <= 12'h252;
        src61 <= 12'h31d;
        src62 <= 12'h111;
        src63 <= 12'he2a;
        src64 <= 12'hd88;
        src65 <= 12'h8df;
        src66 <= 12'he88;
        src67 <= 12'h610;
        src68 <= 12'h29b;
        src69 <= 12'ha67;
        src70 <= 12'h66f;
        src71 <= 12'h7d7;
        src72 <= 12'h311;
        src73 <= 12'h932;
        src74 <= 12'hb7d;
        src75 <= 12'h8ed;
        src76 <= 12'h124;
        src77 <= 12'h20f;
        src78 <= 12'h864;
        src79 <= 12'hdbb;
        src80 <= 12'h5c7;
        src81 <= 12'h51f;
        src82 <= 12'h5da;
        src83 <= 12'he33;
        src84 <= 12'hb6d;
        src85 <= 12'h241;
        src86 <= 12'hdde;
        src87 <= 12'hf07;
        src88 <= 12'h6d7;
        src89 <= 12'h4e4;
        src90 <= 12'he8a;
        src91 <= 12'h33;
        src92 <= 12'hdab;
        src93 <= 12'h125;
        src94 <= 12'hb1a;
        src95 <= 12'h8b9;
        src96 <= 12'hcb3;
        src97 <= 12'ha27;
        src98 <= 12'h47e;
        src99 <= 12'h481;
        src100 <= 12'h723;
        src101 <= 12'h508;
        src102 <= 12'h53;
        src103 <= 12'h433;
        src104 <= 12'hfea;
        src105 <= 12'h1a3;
        src106 <= 12'h80b;
        src107 <= 12'h7c7;
        src108 <= 12'h8db;
        src109 <= 12'h13e;
        src110 <= 12'hee2;
        src111 <= 12'hf7e;
        src112 <= 12'hc6e;
        src113 <= 12'ha77;
        src114 <= 12'hddb;
        src115 <= 12'h472;
        src116 <= 12'hec0;
        src117 <= 12'hd07;
        src118 <= 12'h95f;
        src119 <= 12'h93f;
        src120 <= 12'hfbb;
        src121 <= 12'h32c;
        src122 <= 12'h749;
        src123 <= 12'h8b;
        src124 <= 12'h41e;
        src125 <= 12'h64d;
        src126 <= 12'h2cd;
        src127 <= 12'heca;
        src128 <= 12'h83a;
        src129 <= 12'hed2;
        src130 <= 12'he0b;
        src131 <= 12'hf34;
        src132 <= 12'hf61;
        src133 <= 12'h6d4;
        src134 <= 12'h7cb;
        src135 <= 12'hf6e;
        src136 <= 12'h62d;
        src137 <= 12'h2cb;
        src138 <= 12'hf17;
        src139 <= 12'h7e5;
        src140 <= 12'h82;
        src141 <= 12'h49d;
        src142 <= 12'h8fc;
        src143 <= 12'h8ee;
        src144 <= 12'h20f;
        src145 <= 12'ha20;
        src146 <= 12'h4dd;
        src147 <= 12'hf30;
        src148 <= 12'hae1;
        src149 <= 12'hcd6;
        src150 <= 12'h397;
        src151 <= 12'h616;
        src152 <= 12'hbb8;
        src153 <= 12'h3de;
        src154 <= 12'h927;
        src155 <= 12'h1b6;
        src156 <= 12'h5e9;
        src157 <= 12'hf5a;
        src158 <= 12'h8d5;
        src159 <= 12'hca4;
        src160 <= 12'h575;
        src161 <= 12'h7d7;
        src162 <= 12'hdab;
        src163 <= 12'h7aa;
        src164 <= 12'h6d4;
        src165 <= 12'he62;
        src166 <= 12'hfe7;
        src167 <= 12'hbb3;
        src168 <= 12'h10c;
        src169 <= 12'he2f;
        src170 <= 12'he45;
        src171 <= 12'h7f4;
        src172 <= 12'h865;
        src173 <= 12'h2c5;
        src174 <= 12'ha9d;
        src175 <= 12'hbb8;
        src176 <= 12'h2f4;
        src177 <= 12'h21e;
        src178 <= 12'hd85;
        src179 <= 12'hb1d;
        src180 <= 12'h3f9;
        src181 <= 12'h76d;
        src182 <= 12'h575;
        src183 <= 12'h71a;
        src184 <= 12'h8d5;
        src185 <= 12'hafc;
        src186 <= 12'hd2f;
        src187 <= 12'h38c;
        src188 <= 12'h4da;
        exp <= 20'h5f172;
        #1
        src0 <= 12'h560;
        src1 <= 12'h352;
        src2 <= 12'h6b9;
        src3 <= 12'h856;
        src4 <= 12'h9f7;
        src5 <= 12'h76f;
        src6 <= 12'hd9f;
        src7 <= 12'hbac;
        src8 <= 12'he22;
        src9 <= 12'hb3;
        src10 <= 12'hc01;
        src11 <= 12'he3e;
        src12 <= 12'hab1;
        src13 <= 12'h7c4;
        src14 <= 12'h797;
        src15 <= 12'h3f8;
        src16 <= 12'h19;
        src17 <= 12'hcf8;
        src18 <= 12'he8f;
        src19 <= 12'h4fa;
        src20 <= 12'hda1;
        src21 <= 12'h9ff;
        src22 <= 12'h4cf;
        src23 <= 12'h72;
        src24 <= 12'hfa7;
        src25 <= 12'hbdb;
        src26 <= 12'h31e;
        src27 <= 12'h32b;
        src28 <= 12'hd82;
        src29 <= 12'h188;
        src30 <= 12'h18a;
        src31 <= 12'h9fe;
        src32 <= 12'h369;
        src33 <= 12'h18e;
        src34 <= 12'h22a;
        src35 <= 12'h374;
        src36 <= 12'h129;
        src37 <= 12'hcd1;
        src38 <= 12'h9f4;
        src39 <= 12'h5d2;
        src40 <= 12'h736;
        src41 <= 12'hd75;
        src42 <= 12'h40b;
        src43 <= 12'h6b;
        src44 <= 12'h2e5;
        src45 <= 12'h45a;
        src46 <= 12'hef6;
        src47 <= 12'h731;
        src48 <= 12'h922;
        src49 <= 12'h8d3;
        src50 <= 12'h329;
        src51 <= 12'h3d0;
        src52 <= 12'h752;
        src53 <= 12'hc43;
        src54 <= 12'h397;
        src55 <= 12'haca;
        src56 <= 12'hc19;
        src57 <= 12'hf04;
        src58 <= 12'h3d7;
        src59 <= 12'hca7;
        src60 <= 12'h288;
        src61 <= 12'h15e;
        src62 <= 12'h442;
        src63 <= 12'hdbf;
        src64 <= 12'habc;
        src65 <= 12'h198;
        src66 <= 12'h102;
        src67 <= 12'h926;
        src68 <= 12'ha8b;
        src69 <= 12'h284;
        src70 <= 12'hd16;
        src71 <= 12'h137;
        src72 <= 12'h4bd;
        src73 <= 12'h353;
        src74 <= 12'h31;
        src75 <= 12'hd69;
        src76 <= 12'h3ba;
        src77 <= 12'h85a;
        src78 <= 12'hc0a;
        src79 <= 12'he35;
        src80 <= 12'h282;
        src81 <= 12'hc7b;
        src82 <= 12'h71c;
        src83 <= 12'hae2;
        src84 <= 12'he91;
        src85 <= 12'h15b;
        src86 <= 12'h83;
        src87 <= 12'hbaa;
        src88 <= 12'h12e;
        src89 <= 12'h8d6;
        src90 <= 12'h6e3;
        src91 <= 12'h5fc;
        src92 <= 12'h880;
        src93 <= 12'h50f;
        src94 <= 12'hda0;
        src95 <= 12'heee;
        src96 <= 12'ha56;
        src97 <= 12'h669;
        src98 <= 12'haa3;
        src99 <= 12'hb27;
        src100 <= 12'hb37;
        src101 <= 12'hb5;
        src102 <= 12'h58a;
        src103 <= 12'hadd;
        src104 <= 12'h59c;
        src105 <= 12'h46;
        src106 <= 12'h2c1;
        src107 <= 12'hfbb;
        src108 <= 12'hcc6;
        src109 <= 12'h757;
        src110 <= 12'h3e2;
        src111 <= 12'h657;
        src112 <= 12'h3a9;
        src113 <= 12'h8fc;
        src114 <= 12'ha39;
        src115 <= 12'hb86;
        src116 <= 12'h133;
        src117 <= 12'hb14;
        src118 <= 12'haa3;
        src119 <= 12'h3ba;
        src120 <= 12'ha25;
        src121 <= 12'h913;
        src122 <= 12'h147;
        src123 <= 12'hcf0;
        src124 <= 12'h71;
        src125 <= 12'hdb8;
        src126 <= 12'h640;
        src127 <= 12'hb26;
        src128 <= 12'h4e;
        src129 <= 12'h214;
        src130 <= 12'hc8c;
        src131 <= 12'h398;
        src132 <= 12'h496;
        src133 <= 12'h103;
        src134 <= 12'ha7c;
        src135 <= 12'ha0;
        src136 <= 12'ha8d;
        src137 <= 12'h373;
        src138 <= 12'h4b;
        src139 <= 12'hf7d;
        src140 <= 12'h30b;
        src141 <= 12'h913;
        src142 <= 12'h8dd;
        src143 <= 12'h879;
        src144 <= 12'h33a;
        src145 <= 12'hba1;
        src146 <= 12'hbbb;
        src147 <= 12'h4be;
        src148 <= 12'h846;
        src149 <= 12'h7fd;
        src150 <= 12'hfa3;
        src151 <= 12'he84;
        src152 <= 12'hdab;
        src153 <= 12'h815;
        src154 <= 12'h444;
        src155 <= 12'h45;
        src156 <= 12'h5f3;
        src157 <= 12'h1c7;
        src158 <= 12'hfc7;
        src159 <= 12'h6c1;
        src160 <= 12'h680;
        src161 <= 12'h3cc;
        src162 <= 12'h391;
        src163 <= 12'haea;
        src164 <= 12'h774;
        src165 <= 12'h438;
        src166 <= 12'h81c;
        src167 <= 12'h43f;
        src168 <= 12'h67e;
        src169 <= 12'h6ae;
        src170 <= 12'h3f6;
        src171 <= 12'h43;
        src172 <= 12'hb7b;
        src173 <= 12'h70b;
        src174 <= 12'h178;
        src175 <= 12'h37;
        src176 <= 12'h6b8;
        src177 <= 12'h8bd;
        src178 <= 12'h8b8;
        src179 <= 12'h410;
        src180 <= 12'hf9a;
        src181 <= 12'h408;
        src182 <= 12'h5fb;
        src183 <= 12'hf80;
        src184 <= 12'hc31;
        src185 <= 12'h585;
        src186 <= 12'h616;
        src187 <= 12'h3a6;
        src188 <= 12'h555;
        exp <= 20'h5636c;
        #1
        src0 <= 12'h2c5;
        src1 <= 12'h965;
        src2 <= 12'h28e;
        src3 <= 12'h3b6;
        src4 <= 12'h90b;
        src5 <= 12'h2a2;
        src6 <= 12'h68b;
        src7 <= 12'h8a5;
        src8 <= 12'h984;
        src9 <= 12'hf2c;
        src10 <= 12'h288;
        src11 <= 12'h451;
        src12 <= 12'h72;
        src13 <= 12'h821;
        src14 <= 12'h785;
        src15 <= 12'h8ca;
        src16 <= 12'hcef;
        src17 <= 12'hbd6;
        src18 <= 12'h8ea;
        src19 <= 12'h81d;
        src20 <= 12'h3dc;
        src21 <= 12'hbc2;
        src22 <= 12'h946;
        src23 <= 12'h9a5;
        src24 <= 12'h9f9;
        src25 <= 12'h8c1;
        src26 <= 12'haa;
        src27 <= 12'he2e;
        src28 <= 12'h7d8;
        src29 <= 12'he0f;
        src30 <= 12'h409;
        src31 <= 12'h49b;
        src32 <= 12'hafa;
        src33 <= 12'hf32;
        src34 <= 12'hcad;
        src35 <= 12'h7c4;
        src36 <= 12'h4cb;
        src37 <= 12'h1fc;
        src38 <= 12'h17d;
        src39 <= 12'h799;
        src40 <= 12'h54;
        src41 <= 12'h121;
        src42 <= 12'h35b;
        src43 <= 12'h338;
        src44 <= 12'h749;
        src45 <= 12'h84d;
        src46 <= 12'h5ab;
        src47 <= 12'hd19;
        src48 <= 12'h550;
        src49 <= 12'he95;
        src50 <= 12'he5d;
        src51 <= 12'hfed;
        src52 <= 12'h71b;
        src53 <= 12'h5c5;
        src54 <= 12'h143;
        src55 <= 12'hc55;
        src56 <= 12'h37;
        src57 <= 12'h786;
        src58 <= 12'h6d5;
        src59 <= 12'hd0f;
        src60 <= 12'h5bb;
        src61 <= 12'h37d;
        src62 <= 12'hd36;
        src63 <= 12'hc4d;
        src64 <= 12'hf12;
        src65 <= 12'hb41;
        src66 <= 12'h94b;
        src67 <= 12'hdfe;
        src68 <= 12'h525;
        src69 <= 12'h53c;
        src70 <= 12'h4fb;
        src71 <= 12'h83d;
        src72 <= 12'hcf1;
        src73 <= 12'h6cb;
        src74 <= 12'hf47;
        src75 <= 12'ha8f;
        src76 <= 12'hec9;
        src77 <= 12'h545;
        src78 <= 12'h11a;
        src79 <= 12'h138;
        src80 <= 12'hb5b;
        src81 <= 12'ha49;
        src82 <= 12'h1fd;
        src83 <= 12'h975;
        src84 <= 12'h2a5;
        src85 <= 12'h76b;
        src86 <= 12'h645;
        src87 <= 12'h748;
        src88 <= 12'haef;
        src89 <= 12'h69f;
        src90 <= 12'hc19;
        src91 <= 12'he94;
        src92 <= 12'hdc7;
        src93 <= 12'h315;
        src94 <= 12'h839;
        src95 <= 12'hfcf;
        src96 <= 12'h33e;
        src97 <= 12'h306;
        src98 <= 12'hfc7;
        src99 <= 12'h326;
        src100 <= 12'ha2d;
        src101 <= 12'hc05;
        src102 <= 12'hca1;
        src103 <= 12'hd02;
        src104 <= 12'hcd3;
        src105 <= 12'had9;
        src106 <= 12'he3a;
        src107 <= 12'h2e7;
        src108 <= 12'h66a;
        src109 <= 12'h2e7;
        src110 <= 12'h1ec;
        src111 <= 12'h707;
        src112 <= 12'hc37;
        src113 <= 12'hdf2;
        src114 <= 12'h71c;
        src115 <= 12'hf8a;
        src116 <= 12'hb43;
        src117 <= 12'h423;
        src118 <= 12'h4d9;
        src119 <= 12'hacb;
        src120 <= 12'h79;
        src121 <= 12'hd6e;
        src122 <= 12'he6;
        src123 <= 12'hd89;
        src124 <= 12'hce9;
        src125 <= 12'hd08;
        src126 <= 12'heb8;
        src127 <= 12'h893;
        src128 <= 12'h386;
        src129 <= 12'hccf;
        src130 <= 12'h1fd;
        src131 <= 12'h7be;
        src132 <= 12'hb1b;
        src133 <= 12'h714;
        src134 <= 12'hb0c;
        src135 <= 12'hce4;
        src136 <= 12'hf7c;
        src137 <= 12'hbf0;
        src138 <= 12'h1cb;
        src139 <= 12'h735;
        src140 <= 12'h81;
        src141 <= 12'h9e2;
        src142 <= 12'hc12;
        src143 <= 12'had5;
        src144 <= 12'hefd;
        src145 <= 12'haae;
        src146 <= 12'h7ff;
        src147 <= 12'hc2a;
        src148 <= 12'h628;
        src149 <= 12'h4d0;
        src150 <= 12'heff;
        src151 <= 12'hee5;
        src152 <= 12'h44e;
        src153 <= 12'h58c;
        src154 <= 12'hba2;
        src155 <= 12'h58f;
        src156 <= 12'h83b;
        src157 <= 12'h285;
        src158 <= 12'ha87;
        src159 <= 12'h50e;
        src160 <= 12'h4c7;
        src161 <= 12'h91e;
        src162 <= 12'h9b6;
        src163 <= 12'h7ce;
        src164 <= 12'hcd6;
        src165 <= 12'h66e;
        src166 <= 12'he51;
        src167 <= 12'hb6e;
        src168 <= 12'h25d;
        src169 <= 12'ha88;
        src170 <= 12'h62b;
        src171 <= 12'hd4d;
        src172 <= 12'h654;
        src173 <= 12'hcb9;
        src174 <= 12'h8c6;
        src175 <= 12'hbd;
        src176 <= 12'h8b0;
        src177 <= 12'hd57;
        src178 <= 12'hb8b;
        src179 <= 12'hd3a;
        src180 <= 12'he90;
        src181 <= 12'h252;
        src182 <= 12'h15e;
        src183 <= 12'h1cb;
        src184 <= 12'hf5d;
        src185 <= 12'h985;
        src186 <= 12'h5d6;
        src187 <= 12'haea;
        src188 <= 12'hf1b;
        exp <= 20'h63d64;
        #1
        src0 <= 12'hfeb;
        src1 <= 12'h37f;
        src2 <= 12'hd7;
        src3 <= 12'hcae;
        src4 <= 12'h5cf;
        src5 <= 12'hff1;
        src6 <= 12'hf16;
        src7 <= 12'h849;
        src8 <= 12'h23a;
        src9 <= 12'h321;
        src10 <= 12'h50f;
        src11 <= 12'hd29;
        src12 <= 12'h8c0;
        src13 <= 12'h7d6;
        src14 <= 12'h6b9;
        src15 <= 12'h278;
        src16 <= 12'hcb4;
        src17 <= 12'h6a0;
        src18 <= 12'hcdc;
        src19 <= 12'h61;
        src20 <= 12'h2a8;
        src21 <= 12'hcb2;
        src22 <= 12'hf27;
        src23 <= 12'h4d9;
        src24 <= 12'h189;
        src25 <= 12'h409;
        src26 <= 12'h965;
        src27 <= 12'hd4a;
        src28 <= 12'h49;
        src29 <= 12'h71d;
        src30 <= 12'h187;
        src31 <= 12'hf8;
        src32 <= 12'he68;
        src33 <= 12'hc09;
        src34 <= 12'h2de;
        src35 <= 12'h7d6;
        src36 <= 12'hda3;
        src37 <= 12'ha23;
        src38 <= 12'hf84;
        src39 <= 12'hca9;
        src40 <= 12'he5d;
        src41 <= 12'h581;
        src42 <= 12'h85;
        src43 <= 12'hbcf;
        src44 <= 12'ha60;
        src45 <= 12'h781;
        src46 <= 12'h180;
        src47 <= 12'h8bc;
        src48 <= 12'hcc8;
        src49 <= 12'h704;
        src50 <= 12'h695;
        src51 <= 12'hf1b;
        src52 <= 12'h5cf;
        src53 <= 12'h505;
        src54 <= 12'h6e2;
        src55 <= 12'hb16;
        src56 <= 12'hebf;
        src57 <= 12'ha0f;
        src58 <= 12'hf21;
        src59 <= 12'h30a;
        src60 <= 12'hf68;
        src61 <= 12'h39d;
        src62 <= 12'h1d6;
        src63 <= 12'h4ba;
        src64 <= 12'h923;
        src65 <= 12'h86b;
        src66 <= 12'h62c;
        src67 <= 12'h145;
        src68 <= 12'h74f;
        src69 <= 12'he9c;
        src70 <= 12'h498;
        src71 <= 12'h1a1;
        src72 <= 12'h3c1;
        src73 <= 12'ha47;
        src74 <= 12'hbfa;
        src75 <= 12'hf71;
        src76 <= 12'hb73;
        src77 <= 12'h63b;
        src78 <= 12'he55;
        src79 <= 12'h9ee;
        src80 <= 12'h646;
        src81 <= 12'h5a;
        src82 <= 12'hb3a;
        src83 <= 12'h16b;
        src84 <= 12'h78f;
        src85 <= 12'h918;
        src86 <= 12'h37d;
        src87 <= 12'h7be;
        src88 <= 12'hb89;
        src89 <= 12'h977;
        src90 <= 12'h86a;
        src91 <= 12'hda6;
        src92 <= 12'h692;
        src93 <= 12'hb53;
        src94 <= 12'h7c2;
        src95 <= 12'h18c;
        src96 <= 12'ha07;
        src97 <= 12'hb50;
        src98 <= 12'h572;
        src99 <= 12'hf32;
        src100 <= 12'h602;
        src101 <= 12'h8b1;
        src102 <= 12'h13e;
        src103 <= 12'h7f9;
        src104 <= 12'hdc0;
        src105 <= 12'hf78;
        src106 <= 12'h513;
        src107 <= 12'h9d2;
        src108 <= 12'h5c3;
        src109 <= 12'h33c;
        src110 <= 12'h9da;
        src111 <= 12'hb3f;
        src112 <= 12'h21f;
        src113 <= 12'h774;
        src114 <= 12'hf7c;
        src115 <= 12'hd77;
        src116 <= 12'h1b7;
        src117 <= 12'h614;
        src118 <= 12'h3b6;
        src119 <= 12'h450;
        src120 <= 12'h7ad;
        src121 <= 12'hd8d;
        src122 <= 12'hbc;
        src123 <= 12'hc84;
        src124 <= 12'h4b1;
        src125 <= 12'h407;
        src126 <= 12'heee;
        src127 <= 12'ha4c;
        src128 <= 12'hcea;
        src129 <= 12'h1dd;
        src130 <= 12'h32a;
        src131 <= 12'hfb5;
        src132 <= 12'h9eb;
        src133 <= 12'h33a;
        src134 <= 12'h41b;
        src135 <= 12'h1f4;
        src136 <= 12'hf35;
        src137 <= 12'ha09;
        src138 <= 12'hf94;
        src139 <= 12'hced;
        src140 <= 12'h7c;
        src141 <= 12'h692;
        src142 <= 12'h667;
        src143 <= 12'h547;
        src144 <= 12'h90c;
        src145 <= 12'hfb5;
        src146 <= 12'h61b;
        src147 <= 12'h60;
        src148 <= 12'h947;
        src149 <= 12'h3a5;
        src150 <= 12'h720;
        src151 <= 12'h336;
        src152 <= 12'h2a3;
        src153 <= 12'hf85;
        src154 <= 12'he64;
        src155 <= 12'hb88;
        src156 <= 12'h4f0;
        src157 <= 12'he3;
        src158 <= 12'h33;
        src159 <= 12'h61f;
        src160 <= 12'hfb2;
        src161 <= 12'h9b2;
        src162 <= 12'h46e;
        src163 <= 12'he3e;
        src164 <= 12'hee1;
        src165 <= 12'h61;
        src166 <= 12'h9d1;
        src167 <= 12'h5c0;
        src168 <= 12'h544;
        src169 <= 12'h303;
        src170 <= 12'h12;
        src171 <= 12'h1c7;
        src172 <= 12'h67c;
        src173 <= 12'h744;
        src174 <= 12'hbdf;
        src175 <= 12'hea7;
        src176 <= 12'h4b9;
        src177 <= 12'h811;
        src178 <= 12'hb7a;
        src179 <= 12'ha7e;
        src180 <= 12'h920;
        src181 <= 12'he62;
        src182 <= 12'haf0;
        src183 <= 12'hd0d;
        src184 <= 12'hfc6;
        src185 <= 12'h82f;
        src186 <= 12'h73c;
        src187 <= 12'hbd3;
        src188 <= 12'hb17;
        exp <= 20'h60035;
        #1
        src0 <= 12'hec1;
        src1 <= 12'hca8;
        src2 <= 12'h52e;
        src3 <= 12'h9af;
        src4 <= 12'hefc;
        src5 <= 12'h660;
        src6 <= 12'h50b;
        src7 <= 12'h3;
        src8 <= 12'h942;
        src9 <= 12'hd2b;
        src10 <= 12'h8b5;
        src11 <= 12'h9b9;
        src12 <= 12'h149;
        src13 <= 12'hd9f;
        src14 <= 12'h71e;
        src15 <= 12'h5cc;
        src16 <= 12'h66e;
        src17 <= 12'h393;
        src18 <= 12'heb5;
        src19 <= 12'h6f9;
        src20 <= 12'h4f0;
        src21 <= 12'he33;
        src22 <= 12'ha16;
        src23 <= 12'h2d1;
        src24 <= 12'h18e;
        src25 <= 12'h45a;
        src26 <= 12'ha7a;
        src27 <= 12'h919;
        src28 <= 12'h559;
        src29 <= 12'hadd;
        src30 <= 12'h65d;
        src31 <= 12'h8dd;
        src32 <= 12'h25a;
        src33 <= 12'hc24;
        src34 <= 12'h34;
        src35 <= 12'hf11;
        src36 <= 12'hfdb;
        src37 <= 12'ha95;
        src38 <= 12'h175;
        src39 <= 12'hc7c;
        src40 <= 12'he73;
        src41 <= 12'h95c;
        src42 <= 12'hb53;
        src43 <= 12'h6bb;
        src44 <= 12'h4c6;
        src45 <= 12'had4;
        src46 <= 12'h9e;
        src47 <= 12'ha3c;
        src48 <= 12'h45;
        src49 <= 12'he70;
        src50 <= 12'h833;
        src51 <= 12'h694;
        src52 <= 12'ha43;
        src53 <= 12'hb45;
        src54 <= 12'hab2;
        src55 <= 12'h698;
        src56 <= 12'he1;
        src57 <= 12'hc90;
        src58 <= 12'hd4a;
        src59 <= 12'h40;
        src60 <= 12'h32c;
        src61 <= 12'h110;
        src62 <= 12'h84e;
        src63 <= 12'ha64;
        src64 <= 12'h773;
        src65 <= 12'ha5;
        src66 <= 12'hcde;
        src67 <= 12'hb2;
        src68 <= 12'h1ae;
        src69 <= 12'h83d;
        src70 <= 12'h4d6;
        src71 <= 12'hd8b;
        src72 <= 12'ha05;
        src73 <= 12'h738;
        src74 <= 12'h99a;
        src75 <= 12'hba1;
        src76 <= 12'hcbf;
        src77 <= 12'h2fc;
        src78 <= 12'h99e;
        src79 <= 12'h584;
        src80 <= 12'h29e;
        src81 <= 12'hf90;
        src82 <= 12'h5b3;
        src83 <= 12'h136;
        src84 <= 12'hfac;
        src85 <= 12'h1c1;
        src86 <= 12'h434;
        src87 <= 12'h893;
        src88 <= 12'h5f7;
        src89 <= 12'h14b;
        src90 <= 12'hb58;
        src91 <= 12'he26;
        src92 <= 12'h81d;
        src93 <= 12'hc50;
        src94 <= 12'h2;
        src95 <= 12'hbb1;
        src96 <= 12'h830;
        src97 <= 12'he9b;
        src98 <= 12'h32a;
        src99 <= 12'hcb;
        src100 <= 12'h37b;
        src101 <= 12'hedb;
        src102 <= 12'hf00;
        src103 <= 12'ha33;
        src104 <= 12'hbd2;
        src105 <= 12'hbb1;
        src106 <= 12'hf26;
        src107 <= 12'hfe9;
        src108 <= 12'hc41;
        src109 <= 12'h39d;
        src110 <= 12'h3f7;
        src111 <= 12'hebb;
        src112 <= 12'he78;
        src113 <= 12'hd4c;
        src114 <= 12'hed1;
        src115 <= 12'hd4;
        src116 <= 12'h5dc;
        src117 <= 12'hf6;
        src118 <= 12'h273;
        src119 <= 12'h273;
        src120 <= 12'h156;
        src121 <= 12'h2dd;
        src122 <= 12'h3e9;
        src123 <= 12'h792;
        src124 <= 12'h450;
        src125 <= 12'h5c8;
        src126 <= 12'hf7e;
        src127 <= 12'h175;
        src128 <= 12'hadf;
        src129 <= 12'h675;
        src130 <= 12'h1d5;
        src131 <= 12'h6ce;
        src132 <= 12'hef0;
        src133 <= 12'h835;
        src134 <= 12'hc6b;
        src135 <= 12'h988;
        src136 <= 12'h369;
        src137 <= 12'ha7c;
        src138 <= 12'h944;
        src139 <= 12'h4bf;
        src140 <= 12'h7bd;
        src141 <= 12'h473;
        src142 <= 12'hc31;
        src143 <= 12'h827;
        src144 <= 12'hece;
        src145 <= 12'hbd1;
        src146 <= 12'h153;
        src147 <= 12'h270;
        src148 <= 12'h5f0;
        src149 <= 12'h81b;
        src150 <= 12'he4c;
        src151 <= 12'h8d2;
        src152 <= 12'h3ee;
        src153 <= 12'h40e;
        src154 <= 12'h550;
        src155 <= 12'h954;
        src156 <= 12'h1e1;
        src157 <= 12'ha26;
        src158 <= 12'hc98;
        src159 <= 12'he2a;
        src160 <= 12'hfaf;
        src161 <= 12'h675;
        src162 <= 12'h370;
        src163 <= 12'he88;
        src164 <= 12'h172;
        src165 <= 12'hf3;
        src166 <= 12'h3f3;
        src167 <= 12'h32e;
        src168 <= 12'hfe0;
        src169 <= 12'hf6;
        src170 <= 12'h972;
        src171 <= 12'h417;
        src172 <= 12'hd46;
        src173 <= 12'hfca;
        src174 <= 12'hcf3;
        src175 <= 12'h26b;
        src176 <= 12'h30e;
        src177 <= 12'hc78;
        src178 <= 12'h3f7;
        src179 <= 12'hff4;
        src180 <= 12'h947;
        src181 <= 12'h38d;
        src182 <= 12'h2b3;
        src183 <= 12'h659;
        src184 <= 12'h64d;
        src185 <= 12'h695;
        src186 <= 12'h978;
        src187 <= 12'h997;
        src188 <= 12'h78e;
        exp <= 20'h5d518;
        #1
        src0 <= 12'he0e;
        src1 <= 12'h2ee;
        src2 <= 12'h1cb;
        src3 <= 12'hdb7;
        src4 <= 12'h975;
        src5 <= 12'h97a;
        src6 <= 12'h6b2;
        src7 <= 12'h42f;
        src8 <= 12'he3e;
        src9 <= 12'h988;
        src10 <= 12'hf51;
        src11 <= 12'he28;
        src12 <= 12'h84;
        src13 <= 12'h175;
        src14 <= 12'hc71;
        src15 <= 12'h81f;
        src16 <= 12'h492;
        src17 <= 12'hef9;
        src18 <= 12'hf3e;
        src19 <= 12'hd52;
        src20 <= 12'h3d1;
        src21 <= 12'h7c1;
        src22 <= 12'h6b6;
        src23 <= 12'hb42;
        src24 <= 12'h296;
        src25 <= 12'h4ff;
        src26 <= 12'hdc8;
        src27 <= 12'ha65;
        src28 <= 12'hd73;
        src29 <= 12'h9b4;
        src30 <= 12'h48;
        src31 <= 12'h8c3;
        src32 <= 12'hb8a;
        src33 <= 12'hd69;
        src34 <= 12'h168;
        src35 <= 12'h3cc;
        src36 <= 12'hd75;
        src37 <= 12'h621;
        src38 <= 12'hd4b;
        src39 <= 12'h58d;
        src40 <= 12'h3d9;
        src41 <= 12'hb0;
        src42 <= 12'hca9;
        src43 <= 12'h529;
        src44 <= 12'h3d8;
        src45 <= 12'hbb3;
        src46 <= 12'h6e9;
        src47 <= 12'hbac;
        src48 <= 12'habe;
        src49 <= 12'h3d;
        src50 <= 12'h19c;
        src51 <= 12'h21b;
        src52 <= 12'h4f7;
        src53 <= 12'h6ad;
        src54 <= 12'h7b6;
        src55 <= 12'h195;
        src56 <= 12'h892;
        src57 <= 12'hd11;
        src58 <= 12'h65b;
        src59 <= 12'h4a5;
        src60 <= 12'h868;
        src61 <= 12'hef7;
        src62 <= 12'hb5e;
        src63 <= 12'hc00;
        src64 <= 12'hbf4;
        src65 <= 12'h278;
        src66 <= 12'hf38;
        src67 <= 12'hecc;
        src68 <= 12'hcc2;
        src69 <= 12'hc76;
        src70 <= 12'hcc3;
        src71 <= 12'h228;
        src72 <= 12'hf93;
        src73 <= 12'h259;
        src74 <= 12'ha72;
        src75 <= 12'h340;
        src76 <= 12'he8a;
        src77 <= 12'h6d4;
        src78 <= 12'h443;
        src79 <= 12'hd3e;
        src80 <= 12'h807;
        src81 <= 12'hb86;
        src82 <= 12'h6de;
        src83 <= 12'he41;
        src84 <= 12'h99d;
        src85 <= 12'he0f;
        src86 <= 12'h4cd;
        src87 <= 12'h58a;
        src88 <= 12'h633;
        src89 <= 12'hd53;
        src90 <= 12'heaa;
        src91 <= 12'h9b1;
        src92 <= 12'hbef;
        src93 <= 12'h44d;
        src94 <= 12'h555;
        src95 <= 12'h234;
        src96 <= 12'h3ac;
        src97 <= 12'h871;
        src98 <= 12'hd8d;
        src99 <= 12'hce9;
        src100 <= 12'hb6;
        src101 <= 12'h9c;
        src102 <= 12'hf4d;
        src103 <= 12'hbd5;
        src104 <= 12'h32c;
        src105 <= 12'h3e3;
        src106 <= 12'hf2d;
        src107 <= 12'h497;
        src108 <= 12'hf03;
        src109 <= 12'ha5a;
        src110 <= 12'hfaa;
        src111 <= 12'h8f7;
        src112 <= 12'hfd5;
        src113 <= 12'h3e8;
        src114 <= 12'h103;
        src115 <= 12'h658;
        src116 <= 12'h635;
        src117 <= 12'hd72;
        src118 <= 12'h47a;
        src119 <= 12'h2ff;
        src120 <= 12'hdf1;
        src121 <= 12'h9e8;
        src122 <= 12'hd84;
        src123 <= 12'h310;
        src124 <= 12'hc98;
        src125 <= 12'h372;
        src126 <= 12'hd02;
        src127 <= 12'h285;
        src128 <= 12'hea8;
        src129 <= 12'ha88;
        src130 <= 12'hd8e;
        src131 <= 12'h862;
        src132 <= 12'h169;
        src133 <= 12'hf6c;
        src134 <= 12'hae0;
        src135 <= 12'hb09;
        src136 <= 12'he60;
        src137 <= 12'hefa;
        src138 <= 12'h6;
        src139 <= 12'ha1f;
        src140 <= 12'h8fb;
        src141 <= 12'h331;
        src142 <= 12'he6c;
        src143 <= 12'h897;
        src144 <= 12'hdd;
        src145 <= 12'h8d4;
        src146 <= 12'hed0;
        src147 <= 12'hed4;
        src148 <= 12'h302;
        src149 <= 12'h624;
        src150 <= 12'hc0e;
        src151 <= 12'h845;
        src152 <= 12'h648;
        src153 <= 12'hea1;
        src154 <= 12'h9c2;
        src155 <= 12'ha6c;
        src156 <= 12'h7a2;
        src157 <= 12'h970;
        src158 <= 12'h1fd;
        src159 <= 12'h65;
        src160 <= 12'hd25;
        src161 <= 12'h831;
        src162 <= 12'h62;
        src163 <= 12'h4bf;
        src164 <= 12'hdfe;
        src165 <= 12'h160;
        src166 <= 12'hec5;
        src167 <= 12'h16b;
        src168 <= 12'hc7c;
        src169 <= 12'hb4f;
        src170 <= 12'h3b6;
        src171 <= 12'h242;
        src172 <= 12'h159;
        src173 <= 12'h81;
        src174 <= 12'h620;
        src175 <= 12'hd13;
        src176 <= 12'h65b;
        src177 <= 12'ha7c;
        src178 <= 12'h7d2;
        src179 <= 12'h79d;
        src180 <= 12'h824;
        src181 <= 12'h571;
        src182 <= 12'h9e;
        src183 <= 12'he2f;
        src184 <= 12'h998;
        src185 <= 12'hcae;
        src186 <= 12'hc10;
        src187 <= 12'hd67;
        src188 <= 12'h4b;
        exp <= 20'h63a9d;
        #1
        src0 <= 12'ha88;
        src1 <= 12'h90c;
        src2 <= 12'hb1;
        src3 <= 12'h22d;
        src4 <= 12'h41a;
        src5 <= 12'h1a6;
        src6 <= 12'h5e4;
        src7 <= 12'h4d1;
        src8 <= 12'haec;
        src9 <= 12'h2c7;
        src10 <= 12'hfa3;
        src11 <= 12'he0a;
        src12 <= 12'h454;
        src13 <= 12'hdc6;
        src14 <= 12'h339;
        src15 <= 12'hd54;
        src16 <= 12'hbd2;
        src17 <= 12'hef3;
        src18 <= 12'h704;
        src19 <= 12'h425;
        src20 <= 12'h686;
        src21 <= 12'hf0b;
        src22 <= 12'hd67;
        src23 <= 12'h6c;
        src24 <= 12'hb73;
        src25 <= 12'ha2f;
        src26 <= 12'h37d;
        src27 <= 12'he16;
        src28 <= 12'h57b;
        src29 <= 12'hd94;
        src30 <= 12'ha4f;
        src31 <= 12'h5c9;
        src32 <= 12'h469;
        src33 <= 12'hfeb;
        src34 <= 12'h977;
        src35 <= 12'he73;
        src36 <= 12'hcff;
        src37 <= 12'h73b;
        src38 <= 12'h212;
        src39 <= 12'h726;
        src40 <= 12'ha7f;
        src41 <= 12'h6c2;
        src42 <= 12'ha56;
        src43 <= 12'h606;
        src44 <= 12'hff8;
        src45 <= 12'h400;
        src46 <= 12'hdac;
        src47 <= 12'ha02;
        src48 <= 12'h26c;
        src49 <= 12'hbb5;
        src50 <= 12'ha4d;
        src51 <= 12'hbe;
        src52 <= 12'hce2;
        src53 <= 12'hdf3;
        src54 <= 12'hd94;
        src55 <= 12'hb78;
        src56 <= 12'he41;
        src57 <= 12'hb12;
        src58 <= 12'hba2;
        src59 <= 12'h8c1;
        src60 <= 12'hb85;
        src61 <= 12'hc83;
        src62 <= 12'hc37;
        src63 <= 12'hf95;
        src64 <= 12'h60b;
        src65 <= 12'h97b;
        src66 <= 12'h86f;
        src67 <= 12'hf76;
        src68 <= 12'h9c6;
        src69 <= 12'hc93;
        src70 <= 12'he40;
        src71 <= 12'he02;
        src72 <= 12'he95;
        src73 <= 12'hd48;
        src74 <= 12'h7c9;
        src75 <= 12'had2;
        src76 <= 12'hc20;
        src77 <= 12'h538;
        src78 <= 12'h5f1;
        src79 <= 12'ha67;
        src80 <= 12'hab6;
        src81 <= 12'hfa5;
        src82 <= 12'he82;
        src83 <= 12'h2ff;
        src84 <= 12'ha5a;
        src85 <= 12'h692;
        src86 <= 12'h8d2;
        src87 <= 12'hcd;
        src88 <= 12'h62f;
        src89 <= 12'h4fd;
        src90 <= 12'haab;
        src91 <= 12'hafb;
        src92 <= 12'hee3;
        src93 <= 12'hb8a;
        src94 <= 12'h556;
        src95 <= 12'hc67;
        src96 <= 12'h8cb;
        src97 <= 12'h2cd;
        src98 <= 12'hb;
        src99 <= 12'h43f;
        src100 <= 12'hf62;
        src101 <= 12'h70c;
        src102 <= 12'h5ca;
        src103 <= 12'haca;
        src104 <= 12'h44e;
        src105 <= 12'h716;
        src106 <= 12'h398;
        src107 <= 12'h6cd;
        src108 <= 12'hb20;
        src109 <= 12'hac5;
        src110 <= 12'hb72;
        src111 <= 12'h8cf;
        src112 <= 12'h4f1;
        src113 <= 12'h1f0;
        src114 <= 12'ha99;
        src115 <= 12'he9d;
        src116 <= 12'h3ac;
        src117 <= 12'hfb9;
        src118 <= 12'h10;
        src119 <= 12'h431;
        src120 <= 12'h369;
        src121 <= 12'h7b6;
        src122 <= 12'h4c5;
        src123 <= 12'hbd9;
        src124 <= 12'hd78;
        src125 <= 12'h5ed;
        src126 <= 12'h8c9;
        src127 <= 12'hbd0;
        src128 <= 12'haf8;
        src129 <= 12'h60c;
        src130 <= 12'h1f7;
        src131 <= 12'he31;
        src132 <= 12'hbc9;
        src133 <= 12'h151;
        src134 <= 12'h9b2;
        src135 <= 12'h236;
        src136 <= 12'h7f7;
        src137 <= 12'h855;
        src138 <= 12'h9b0;
        src139 <= 12'h932;
        src140 <= 12'hc45;
        src141 <= 12'hdb2;
        src142 <= 12'he78;
        src143 <= 12'h3ac;
        src144 <= 12'h95b;
        src145 <= 12'he77;
        src146 <= 12'h43e;
        src147 <= 12'h12f;
        src148 <= 12'hb66;
        src149 <= 12'hd9c;
        src150 <= 12'h918;
        src151 <= 12'hcff;
        src152 <= 12'h4c;
        src153 <= 12'h226;
        src154 <= 12'h65c;
        src155 <= 12'h14;
        src156 <= 12'h3da;
        src157 <= 12'h3db;
        src158 <= 12'h306;
        src159 <= 12'hff8;
        src160 <= 12'h4d5;
        src161 <= 12'h460;
        src162 <= 12'hfdb;
        src163 <= 12'h430;
        src164 <= 12'hb22;
        src165 <= 12'hfe8;
        src166 <= 12'h561;
        src167 <= 12'h830;
        src168 <= 12'h473;
        src169 <= 12'hb67;
        src170 <= 12'h497;
        src171 <= 12'he5b;
        src172 <= 12'h9d5;
        src173 <= 12'h543;
        src174 <= 12'h675;
        src175 <= 12'h12a;
        src176 <= 12'h209;
        src177 <= 12'h15f;
        src178 <= 12'h9b9;
        src179 <= 12'h712;
        src180 <= 12'h6b1;
        src181 <= 12'hd29;
        src182 <= 12'h50a;
        src183 <= 12'h449;
        src184 <= 12'he3d;
        src185 <= 12'h173;
        src186 <= 12'h900;
        src187 <= 12'h4d6;
        src188 <= 12'h7d0;
        exp <= 20'h64d7a;
        #1
        src0 <= 12'hb61;
        src1 <= 12'haaa;
        src2 <= 12'hf2d;
        src3 <= 12'h4e7;
        src4 <= 12'hd65;
        src5 <= 12'h70d;
        src6 <= 12'hc4a;
        src7 <= 12'hb00;
        src8 <= 12'h59d;
        src9 <= 12'h28e;
        src10 <= 12'h651;
        src11 <= 12'h1d8;
        src12 <= 12'hbe4;
        src13 <= 12'h4b5;
        src14 <= 12'h3a;
        src15 <= 12'hc12;
        src16 <= 12'h51;
        src17 <= 12'h854;
        src18 <= 12'h61d;
        src19 <= 12'hc6;
        src20 <= 12'h83f;
        src21 <= 12'h161;
        src22 <= 12'h846;
        src23 <= 12'hc56;
        src24 <= 12'h901;
        src25 <= 12'h953;
        src26 <= 12'h285;
        src27 <= 12'h4a7;
        src28 <= 12'h892;
        src29 <= 12'hb6c;
        src30 <= 12'h635;
        src31 <= 12'hf42;
        src32 <= 12'hd35;
        src33 <= 12'haac;
        src34 <= 12'h6b0;
        src35 <= 12'hd6;
        src36 <= 12'hf84;
        src37 <= 12'hd0f;
        src38 <= 12'h4ad;
        src39 <= 12'h194;
        src40 <= 12'h854;
        src41 <= 12'h77b;
        src42 <= 12'h9e2;
        src43 <= 12'hbf1;
        src44 <= 12'h177;
        src45 <= 12'he98;
        src46 <= 12'h967;
        src47 <= 12'hee9;
        src48 <= 12'hebd;
        src49 <= 12'h236;
        src50 <= 12'h7b0;
        src51 <= 12'h4bf;
        src52 <= 12'h46c;
        src53 <= 12'he9f;
        src54 <= 12'hc1c;
        src55 <= 12'hbfb;
        src56 <= 12'hd6;
        src57 <= 12'hfd3;
        src58 <= 12'hbf9;
        src59 <= 12'h754;
        src60 <= 12'h478;
        src61 <= 12'hd42;
        src62 <= 12'ha1d;
        src63 <= 12'he27;
        src64 <= 12'hb2b;
        src65 <= 12'h59e;
        src66 <= 12'h104;
        src67 <= 12'hf92;
        src68 <= 12'h7d6;
        src69 <= 12'hff7;
        src70 <= 12'hf48;
        src71 <= 12'hd51;
        src72 <= 12'h8a3;
        src73 <= 12'hb29;
        src74 <= 12'h738;
        src75 <= 12'h999;
        src76 <= 12'h4;
        src77 <= 12'h3cc;
        src78 <= 12'hf36;
        src79 <= 12'h9a7;
        src80 <= 12'h474;
        src81 <= 12'h33;
        src82 <= 12'hc84;
        src83 <= 12'h910;
        src84 <= 12'hb5;
        src85 <= 12'h2f4;
        src86 <= 12'h41c;
        src87 <= 12'hd1b;
        src88 <= 12'hafb;
        src89 <= 12'h3e;
        src90 <= 12'h32c;
        src91 <= 12'h393;
        src92 <= 12'h285;
        src93 <= 12'h27e;
        src94 <= 12'h774;
        src95 <= 12'hf6;
        src96 <= 12'h759;
        src97 <= 12'hd67;
        src98 <= 12'ha7;
        src99 <= 12'h1bb;
        src100 <= 12'hbdf;
        src101 <= 12'h891;
        src102 <= 12'hc1c;
        src103 <= 12'h977;
        src104 <= 12'h957;
        src105 <= 12'h703;
        src106 <= 12'h666;
        src107 <= 12'h88;
        src108 <= 12'hff7;
        src109 <= 12'hde2;
        src110 <= 12'h3c6;
        src111 <= 12'h3aa;
        src112 <= 12'h9af;
        src113 <= 12'ha5;
        src114 <= 12'he84;
        src115 <= 12'h81;
        src116 <= 12'h556;
        src117 <= 12'h643;
        src118 <= 12'h9fc;
        src119 <= 12'h752;
        src120 <= 12'h540;
        src121 <= 12'h52c;
        src122 <= 12'h6eb;
        src123 <= 12'hbfc;
        src124 <= 12'hc32;
        src125 <= 12'h8ca;
        src126 <= 12'h5df;
        src127 <= 12'h228;
        src128 <= 12'h2c1;
        src129 <= 12'h338;
        src130 <= 12'hbe3;
        src131 <= 12'h9c0;
        src132 <= 12'ha06;
        src133 <= 12'h91;
        src134 <= 12'hfd2;
        src135 <= 12'h8f8;
        src136 <= 12'h298;
        src137 <= 12'hc67;
        src138 <= 12'hb1a;
        src139 <= 12'h9f7;
        src140 <= 12'h206;
        src141 <= 12'h714;
        src142 <= 12'h210;
        src143 <= 12'h4d0;
        src144 <= 12'h2f4;
        src145 <= 12'he87;
        src146 <= 12'h99e;
        src147 <= 12'h965;
        src148 <= 12'h2a9;
        src149 <= 12'h10a;
        src150 <= 12'h88d;
        src151 <= 12'h80b;
        src152 <= 12'hb85;
        src153 <= 12'h167;
        src154 <= 12'h891;
        src155 <= 12'hb0b;
        src156 <= 12'h71a;
        src157 <= 12'ha1d;
        src158 <= 12'hb7b;
        src159 <= 12'h7ba;
        src160 <= 12'heb;
        src161 <= 12'h9f0;
        src162 <= 12'h8ec;
        src163 <= 12'heef;
        src164 <= 12'hf25;
        src165 <= 12'h57a;
        src166 <= 12'hd41;
        src167 <= 12'h4b0;
        src168 <= 12'ha24;
        src169 <= 12'h362;
        src170 <= 12'h961;
        src171 <= 12'h791;
        src172 <= 12'h1b9;
        src173 <= 12'hc80;
        src174 <= 12'hde1;
        src175 <= 12'hab6;
        src176 <= 12'h519;
        src177 <= 12'hd5b;
        src178 <= 12'h154;
        src179 <= 12'h3e1;
        src180 <= 12'hdfb;
        src181 <= 12'h819;
        src182 <= 12'hff1;
        src183 <= 12'ha66;
        src184 <= 12'h996;
        src185 <= 12'hc01;
        src186 <= 12'hf72;
        src187 <= 12'h43c;
        src188 <= 12'hd3;
        exp <= 20'h5dfda;
        #1
        src0 <= 12'h261;
        src1 <= 12'had7;
        src2 <= 12'h163;
        src3 <= 12'h298;
        src4 <= 12'hd94;
        src5 <= 12'h347;
        src6 <= 12'h62d;
        src7 <= 12'h5f2;
        src8 <= 12'hc45;
        src9 <= 12'he4;
        src10 <= 12'hb67;
        src11 <= 12'h8e1;
        src12 <= 12'h2d6;
        src13 <= 12'h1b8;
        src14 <= 12'h37b;
        src15 <= 12'h6e8;
        src16 <= 12'hfa;
        src17 <= 12'hb0f;
        src18 <= 12'hf2e;
        src19 <= 12'h67e;
        src20 <= 12'h106;
        src21 <= 12'h26d;
        src22 <= 12'h6b9;
        src23 <= 12'h433;
        src24 <= 12'h96d;
        src25 <= 12'hf23;
        src26 <= 12'h998;
        src27 <= 12'h2ef;
        src28 <= 12'h2b1;
        src29 <= 12'h1a7;
        src30 <= 12'h1b4;
        src31 <= 12'he28;
        src32 <= 12'h119;
        src33 <= 12'h88c;
        src34 <= 12'h1fb;
        src35 <= 12'h26d;
        src36 <= 12'ha24;
        src37 <= 12'hec2;
        src38 <= 12'h4f9;
        src39 <= 12'h7be;
        src40 <= 12'hbb2;
        src41 <= 12'h4ac;
        src42 <= 12'h746;
        src43 <= 12'hdfc;
        src44 <= 12'h66c;
        src45 <= 12'hdce;
        src46 <= 12'ha00;
        src47 <= 12'h332;
        src48 <= 12'h4a4;
        src49 <= 12'h38a;
        src50 <= 12'h55;
        src51 <= 12'h54f;
        src52 <= 12'h8e8;
        src53 <= 12'h88;
        src54 <= 12'h6d;
        src55 <= 12'h900;
        src56 <= 12'ha28;
        src57 <= 12'h725;
        src58 <= 12'ha87;
        src59 <= 12'h30f;
        src60 <= 12'hbd4;
        src61 <= 12'hf9c;
        src62 <= 12'h17c;
        src63 <= 12'hede;
        src64 <= 12'h8d1;
        src65 <= 12'h19e;
        src66 <= 12'h95b;
        src67 <= 12'h317;
        src68 <= 12'h1e3;
        src69 <= 12'h5ea;
        src70 <= 12'hcd7;
        src71 <= 12'h8cc;
        src72 <= 12'h2d8;
        src73 <= 12'hffb;
        src74 <= 12'hae2;
        src75 <= 12'hae7;
        src76 <= 12'hd0d;
        src77 <= 12'h175;
        src78 <= 12'hb04;
        src79 <= 12'h9f7;
        src80 <= 12'hd98;
        src81 <= 12'h9be;
        src82 <= 12'h1da;
        src83 <= 12'hc8c;
        src84 <= 12'h3a2;
        src85 <= 12'hcaa;
        src86 <= 12'h61a;
        src87 <= 12'h214;
        src88 <= 12'hdb7;
        src89 <= 12'hbb0;
        src90 <= 12'hacf;
        src91 <= 12'he39;
        src92 <= 12'h235;
        src93 <= 12'h10c;
        src94 <= 12'hc9c;
        src95 <= 12'hf7;
        src96 <= 12'h2d;
        src97 <= 12'h5aa;
        src98 <= 12'h955;
        src99 <= 12'h669;
        src100 <= 12'h314;
        src101 <= 12'h9dc;
        src102 <= 12'hbea;
        src103 <= 12'hd6e;
        src104 <= 12'h84c;
        src105 <= 12'h40;
        src106 <= 12'he5;
        src107 <= 12'h82;
        src108 <= 12'h24e;
        src109 <= 12'h453;
        src110 <= 12'h122;
        src111 <= 12'hf5a;
        src112 <= 12'h7e7;
        src113 <= 12'hb44;
        src114 <= 12'hc57;
        src115 <= 12'hdac;
        src116 <= 12'h85e;
        src117 <= 12'h1bf;
        src118 <= 12'h666;
        src119 <= 12'he6a;
        src120 <= 12'h2d4;
        src121 <= 12'hfa5;
        src122 <= 12'h8f7;
        src123 <= 12'h309;
        src124 <= 12'h10d;
        src125 <= 12'h101;
        src126 <= 12'h66c;
        src127 <= 12'ha9f;
        src128 <= 12'hbaa;
        src129 <= 12'h3b3;
        src130 <= 12'hb60;
        src131 <= 12'h62a;
        src132 <= 12'h538;
        src133 <= 12'hda6;
        src134 <= 12'h7b7;
        src135 <= 12'h9a2;
        src136 <= 12'h27d;
        src137 <= 12'hd5b;
        src138 <= 12'hbbd;
        src139 <= 12'hd9f;
        src140 <= 12'h4d4;
        src141 <= 12'hab7;
        src142 <= 12'hd96;
        src143 <= 12'haaf;
        src144 <= 12'hccd;
        src145 <= 12'hb4c;
        src146 <= 12'h5d;
        src147 <= 12'h875;
        src148 <= 12'h310;
        src149 <= 12'h24d;
        src150 <= 12'h191;
        src151 <= 12'h87a;
        src152 <= 12'h7f5;
        src153 <= 12'h746;
        src154 <= 12'h472;
        src155 <= 12'h66f;
        src156 <= 12'h793;
        src157 <= 12'h439;
        src158 <= 12'h790;
        src159 <= 12'hec1;
        src160 <= 12'h4f7;
        src161 <= 12'h2a9;
        src162 <= 12'h115;
        src163 <= 12'h3d;
        src164 <= 12'he4d;
        src165 <= 12'ha27;
        src166 <= 12'h79;
        src167 <= 12'hb3;
        src168 <= 12'h143;
        src169 <= 12'h25e;
        src170 <= 12'h9da;
        src171 <= 12'h5da;
        src172 <= 12'hd15;
        src173 <= 12'h328;
        src174 <= 12'h25c;
        src175 <= 12'h41a;
        src176 <= 12'h54a;
        src177 <= 12'hadf;
        src178 <= 12'hd2f;
        src179 <= 12'h6e4;
        src180 <= 12'h819;
        src181 <= 12'h63c;
        src182 <= 12'h70b;
        src183 <= 12'hdad;
        src184 <= 12'h2cf;
        src185 <= 12'hc81;
        src186 <= 12'h249;
        src187 <= 12'hc44;
        src188 <= 12'hdba;
        exp <= 20'h54ca5;
        #1
        src0 <= 12'h934;
        src1 <= 12'h698;
        src2 <= 12'h4c6;
        src3 <= 12'h993;
        src4 <= 12'hf1b;
        src5 <= 12'h9e6;
        src6 <= 12'h703;
        src7 <= 12'hab4;
        src8 <= 12'ha2b;
        src9 <= 12'h4d5;
        src10 <= 12'h38c;
        src11 <= 12'h1bb;
        src12 <= 12'h4cd;
        src13 <= 12'ha93;
        src14 <= 12'h280;
        src15 <= 12'hda0;
        src16 <= 12'hf84;
        src17 <= 12'hc53;
        src18 <= 12'he3d;
        src19 <= 12'h393;
        src20 <= 12'h164;
        src21 <= 12'hb81;
        src22 <= 12'hbaf;
        src23 <= 12'h685;
        src24 <= 12'hc98;
        src25 <= 12'hf18;
        src26 <= 12'hb97;
        src27 <= 12'h13d;
        src28 <= 12'h21b;
        src29 <= 12'ha73;
        src30 <= 12'h718;
        src31 <= 12'hbb8;
        src32 <= 12'h40;
        src33 <= 12'h7e7;
        src34 <= 12'ha8c;
        src35 <= 12'hbda;
        src36 <= 12'hcc1;
        src37 <= 12'h719;
        src38 <= 12'h454;
        src39 <= 12'h65f;
        src40 <= 12'h5f3;
        src41 <= 12'hb0f;
        src42 <= 12'h1bc;
        src43 <= 12'h7f7;
        src44 <= 12'hfeb;
        src45 <= 12'h2b5;
        src46 <= 12'h9c1;
        src47 <= 12'hce2;
        src48 <= 12'h787;
        src49 <= 12'h2ff;
        src50 <= 12'h98c;
        src51 <= 12'h214;
        src52 <= 12'ha23;
        src53 <= 12'h7db;
        src54 <= 12'h1d8;
        src55 <= 12'h51f;
        src56 <= 12'hd1;
        src57 <= 12'h846;
        src58 <= 12'h6c1;
        src59 <= 12'hec7;
        src60 <= 12'h3c0;
        src61 <= 12'hb50;
        src62 <= 12'h879;
        src63 <= 12'h38c;
        src64 <= 12'h57a;
        src65 <= 12'h14;
        src66 <= 12'hb16;
        src67 <= 12'hcc3;
        src68 <= 12'hd66;
        src69 <= 12'h3ef;
        src70 <= 12'h30b;
        src71 <= 12'h259;
        src72 <= 12'h9ff;
        src73 <= 12'hb7e;
        src74 <= 12'h494;
        src75 <= 12'h250;
        src76 <= 12'hc65;
        src77 <= 12'hb69;
        src78 <= 12'h8ce;
        src79 <= 12'h83f;
        src80 <= 12'h7d3;
        src81 <= 12'he4;
        src82 <= 12'h85f;
        src83 <= 12'hb4b;
        src84 <= 12'h8e6;
        src85 <= 12'h502;
        src86 <= 12'heaa;
        src87 <= 12'h1a4;
        src88 <= 12'h9d6;
        src89 <= 12'ha69;
        src90 <= 12'hc1a;
        src91 <= 12'hc2d;
        src92 <= 12'h90b;
        src93 <= 12'hd2a;
        src94 <= 12'hc4b;
        src95 <= 12'h152;
        src96 <= 12'he16;
        src97 <= 12'h340;
        src98 <= 12'he54;
        src99 <= 12'h91;
        src100 <= 12'h5f1;
        src101 <= 12'hdd5;
        src102 <= 12'h9a8;
        src103 <= 12'hd96;
        src104 <= 12'h5ac;
        src105 <= 12'hb8a;
        src106 <= 12'hdbd;
        src107 <= 12'hb7e;
        src108 <= 12'hd8d;
        src109 <= 12'hb6;
        src110 <= 12'h9a3;
        src111 <= 12'h3fc;
        src112 <= 12'h21f;
        src113 <= 12'he22;
        src114 <= 12'h1b;
        src115 <= 12'h567;
        src116 <= 12'hd71;
        src117 <= 12'h716;
        src118 <= 12'heca;
        src119 <= 12'h14a;
        src120 <= 12'h524;
        src121 <= 12'hd96;
        src122 <= 12'h427;
        src123 <= 12'heaf;
        src124 <= 12'h1e9;
        src125 <= 12'h504;
        src126 <= 12'h512;
        src127 <= 12'h4f1;
        src128 <= 12'h657;
        src129 <= 12'h5e7;
        src130 <= 12'h9a4;
        src131 <= 12'hff2;
        src132 <= 12'hd77;
        src133 <= 12'hb59;
        src134 <= 12'h6dd;
        src135 <= 12'h4a8;
        src136 <= 12'hca7;
        src137 <= 12'h994;
        src138 <= 12'h1b2;
        src139 <= 12'he4b;
        src140 <= 12'h88d;
        src141 <= 12'hbe3;
        src142 <= 12'h6ff;
        src143 <= 12'hf84;
        src144 <= 12'h4c8;
        src145 <= 12'h3c7;
        src146 <= 12'ha90;
        src147 <= 12'h7c2;
        src148 <= 12'h6a1;
        src149 <= 12'hb76;
        src150 <= 12'hac8;
        src151 <= 12'hb5a;
        src152 <= 12'h8b;
        src153 <= 12'h5;
        src154 <= 12'h6a3;
        src155 <= 12'h3c4;
        src156 <= 12'h62e;
        src157 <= 12'h68e;
        src158 <= 12'hbb7;
        src159 <= 12'h1c5;
        src160 <= 12'h102;
        src161 <= 12'h383;
        src162 <= 12'h2da;
        src163 <= 12'hf39;
        src164 <= 12'h740;
        src165 <= 12'h47c;
        src166 <= 12'h29e;
        src167 <= 12'h798;
        src168 <= 12'he56;
        src169 <= 12'h17a;
        src170 <= 12'h6a6;
        src171 <= 12'haef;
        src172 <= 12'h7d;
        src173 <= 12'h876;
        src174 <= 12'h7a7;
        src175 <= 12'hda7;
        src176 <= 12'h2fd;
        src177 <= 12'hb6b;
        src178 <= 12'had5;
        src179 <= 12'h68a;
        src180 <= 12'h988;
        src181 <= 12'h416;
        src182 <= 12'h448;
        src183 <= 12'hcde;
        src184 <= 12'h66e;
        src185 <= 12'h5b1;
        src186 <= 12'h2d9;
        src187 <= 12'h45c;
        src188 <= 12'h2bd;
        exp <= 20'h5c64b;
        #1
        src0 <= 12'h44;
        src1 <= 12'h565;
        src2 <= 12'h452;
        src3 <= 12'h41e;
        src4 <= 12'h7bb;
        src5 <= 12'hde7;
        src6 <= 12'hda1;
        src7 <= 12'h14;
        src8 <= 12'ha00;
        src9 <= 12'h8eb;
        src10 <= 12'h3f3;
        src11 <= 12'h145;
        src12 <= 12'h1f3;
        src13 <= 12'hc71;
        src14 <= 12'he1c;
        src15 <= 12'h188;
        src16 <= 12'h584;
        src17 <= 12'h435;
        src18 <= 12'hc53;
        src19 <= 12'hd64;
        src20 <= 12'hc2b;
        src21 <= 12'h596;
        src22 <= 12'hf3c;
        src23 <= 12'ha74;
        src24 <= 12'h4b1;
        src25 <= 12'h1a0;
        src26 <= 12'h15d;
        src27 <= 12'he6b;
        src28 <= 12'hc4a;
        src29 <= 12'h85e;
        src30 <= 12'ha4b;
        src31 <= 12'h9af;
        src32 <= 12'hef9;
        src33 <= 12'hcdb;
        src34 <= 12'h473;
        src35 <= 12'h811;
        src36 <= 12'h5a8;
        src37 <= 12'h38;
        src38 <= 12'h886;
        src39 <= 12'haff;
        src40 <= 12'h76a;
        src41 <= 12'h906;
        src42 <= 12'he13;
        src43 <= 12'he1b;
        src44 <= 12'hc5b;
        src45 <= 12'he9b;
        src46 <= 12'h88f;
        src47 <= 12'h92c;
        src48 <= 12'h342;
        src49 <= 12'h901;
        src50 <= 12'h7c6;
        src51 <= 12'h6af;
        src52 <= 12'h4f5;
        src53 <= 12'h35f;
        src54 <= 12'h35;
        src55 <= 12'h3ae;
        src56 <= 12'hb16;
        src57 <= 12'h70f;
        src58 <= 12'hf55;
        src59 <= 12'he6e;
        src60 <= 12'hbca;
        src61 <= 12'h16d;
        src62 <= 12'h8d2;
        src63 <= 12'h628;
        src64 <= 12'hce2;
        src65 <= 12'hae5;
        src66 <= 12'h82f;
        src67 <= 12'hbb0;
        src68 <= 12'h501;
        src69 <= 12'h287;
        src70 <= 12'h358;
        src71 <= 12'hb10;
        src72 <= 12'he94;
        src73 <= 12'h968;
        src74 <= 12'hf5d;
        src75 <= 12'hc1c;
        src76 <= 12'hce0;
        src77 <= 12'hf8a;
        src78 <= 12'h5a6;
        src79 <= 12'h639;
        src80 <= 12'ha83;
        src81 <= 12'h472;
        src82 <= 12'hb9d;
        src83 <= 12'h940;
        src84 <= 12'h91e;
        src85 <= 12'hca;
        src86 <= 12'h229;
        src87 <= 12'h811;
        src88 <= 12'h678;
        src89 <= 12'h3f7;
        src90 <= 12'h72a;
        src91 <= 12'hbf0;
        src92 <= 12'hfa3;
        src93 <= 12'hc5c;
        src94 <= 12'hc4a;
        src95 <= 12'h83f;
        src96 <= 12'h471;
        src97 <= 12'h38c;
        src98 <= 12'hc4d;
        src99 <= 12'ha8e;
        src100 <= 12'h700;
        src101 <= 12'h322;
        src102 <= 12'ha1;
        src103 <= 12'hf59;
        src104 <= 12'hbc2;
        src105 <= 12'hac9;
        src106 <= 12'h834;
        src107 <= 12'h31;
        src108 <= 12'hb8e;
        src109 <= 12'h360;
        src110 <= 12'h15f;
        src111 <= 12'h5f8;
        src112 <= 12'h59;
        src113 <= 12'h654;
        src114 <= 12'hdff;
        src115 <= 12'hd06;
        src116 <= 12'h415;
        src117 <= 12'ha65;
        src118 <= 12'hb63;
        src119 <= 12'h626;
        src120 <= 12'h59f;
        src121 <= 12'h70c;
        src122 <= 12'h31a;
        src123 <= 12'h18d;
        src124 <= 12'hb0c;
        src125 <= 12'h8e3;
        src126 <= 12'h9ac;
        src127 <= 12'h9b8;
        src128 <= 12'h82e;
        src129 <= 12'h51d;
        src130 <= 12'hafe;
        src131 <= 12'hbe8;
        src132 <= 12'hea1;
        src133 <= 12'h43;
        src134 <= 12'h940;
        src135 <= 12'hb26;
        src136 <= 12'h3f7;
        src137 <= 12'h2eb;
        src138 <= 12'h673;
        src139 <= 12'h157;
        src140 <= 12'haea;
        src141 <= 12'hea7;
        src142 <= 12'h57;
        src143 <= 12'h2a8;
        src144 <= 12'h53;
        src145 <= 12'hb70;
        src146 <= 12'hc29;
        src147 <= 12'h8d7;
        src148 <= 12'h597;
        src149 <= 12'h32;
        src150 <= 12'hd25;
        src151 <= 12'h97d;
        src152 <= 12'h6d3;
        src153 <= 12'hb4f;
        src154 <= 12'h970;
        src155 <= 12'h77f;
        src156 <= 12'he85;
        src157 <= 12'h7ff;
        src158 <= 12'hdd9;
        src159 <= 12'hd19;
        src160 <= 12'hcea;
        src161 <= 12'hb3c;
        src162 <= 12'h455;
        src163 <= 12'h7ee;
        src164 <= 12'hfd0;
        src165 <= 12'hc4c;
        src166 <= 12'hcd3;
        src167 <= 12'h548;
        src168 <= 12'hb79;
        src169 <= 12'h301;
        src170 <= 12'h7c1;
        src171 <= 12'hf18;
        src172 <= 12'he26;
        src173 <= 12'h48f;
        src174 <= 12'ha7;
        src175 <= 12'hd85;
        src176 <= 12'h456;
        src177 <= 12'hdb9;
        src178 <= 12'h65;
        src179 <= 12'hd1;
        src180 <= 12'h7c;
        src181 <= 12'he44;
        src182 <= 12'h305;
        src183 <= 12'hbce;
        src184 <= 12'h4f0;
        src185 <= 12'h869;
        src186 <= 12'h820;
        src187 <= 12'hdc9;
        src188 <= 12'h2df;
        exp <= 20'h60360;
        #1
        src0 <= 12'he8c;
        src1 <= 12'h9cc;
        src2 <= 12'hd00;
        src3 <= 12'ha3c;
        src4 <= 12'h8bb;
        src5 <= 12'hc36;
        src6 <= 12'hcc4;
        src7 <= 12'he8f;
        src8 <= 12'hfd8;
        src9 <= 12'hca1;
        src10 <= 12'ha01;
        src11 <= 12'h926;
        src12 <= 12'hd8;
        src13 <= 12'h8bb;
        src14 <= 12'hb4d;
        src15 <= 12'hce5;
        src16 <= 12'h137;
        src17 <= 12'hf5c;
        src18 <= 12'h9a3;
        src19 <= 12'h3e3;
        src20 <= 12'h9e4;
        src21 <= 12'h73b;
        src22 <= 12'h94c;
        src23 <= 12'h6b3;
        src24 <= 12'hc71;
        src25 <= 12'hf61;
        src26 <= 12'hddc;
        src27 <= 12'hc8c;
        src28 <= 12'h29f;
        src29 <= 12'h5b2;
        src30 <= 12'h74c;
        src31 <= 12'ha96;
        src32 <= 12'he00;
        src33 <= 12'h785;
        src34 <= 12'hb1e;
        src35 <= 12'h345;
        src36 <= 12'hf9c;
        src37 <= 12'h93a;
        src38 <= 12'h16b;
        src39 <= 12'h19b;
        src40 <= 12'ha1b;
        src41 <= 12'hebd;
        src42 <= 12'hbdb;
        src43 <= 12'h668;
        src44 <= 12'h350;
        src45 <= 12'h154;
        src46 <= 12'h686;
        src47 <= 12'hab4;
        src48 <= 12'hfc8;
        src49 <= 12'hc1a;
        src50 <= 12'hc7;
        src51 <= 12'haee;
        src52 <= 12'hbc6;
        src53 <= 12'hf9e;
        src54 <= 12'hc58;
        src55 <= 12'h93f;
        src56 <= 12'h88d;
        src57 <= 12'h57d;
        src58 <= 12'hc0a;
        src59 <= 12'h143;
        src60 <= 12'hcff;
        src61 <= 12'hc86;
        src62 <= 12'h214;
        src63 <= 12'h1de;
        src64 <= 12'h94a;
        src65 <= 12'ha45;
        src66 <= 12'hb04;
        src67 <= 12'h450;
        src68 <= 12'hdec;
        src69 <= 12'hb46;
        src70 <= 12'h3d5;
        src71 <= 12'hc66;
        src72 <= 12'hf35;
        src73 <= 12'h1c;
        src74 <= 12'hd6f;
        src75 <= 12'h505;
        src76 <= 12'h5c;
        src77 <= 12'h4a;
        src78 <= 12'h5f0;
        src79 <= 12'h732;
        src80 <= 12'h92d;
        src81 <= 12'hbf4;
        src82 <= 12'hd95;
        src83 <= 12'h772;
        src84 <= 12'h951;
        src85 <= 12'h68e;
        src86 <= 12'hd78;
        src87 <= 12'ha5;
        src88 <= 12'h53c;
        src89 <= 12'hfd1;
        src90 <= 12'h5a;
        src91 <= 12'h97f;
        src92 <= 12'hed5;
        src93 <= 12'h8bb;
        src94 <= 12'h7eb;
        src95 <= 12'h7ac;
        src96 <= 12'hb1c;
        src97 <= 12'hfe;
        src98 <= 12'h4ff;
        src99 <= 12'hfcf;
        src100 <= 12'haaf;
        src101 <= 12'h8de;
        src102 <= 12'h971;
        src103 <= 12'h46a;
        src104 <= 12'hb2d;
        src105 <= 12'hc0a;
        src106 <= 12'h64a;
        src107 <= 12'h5cb;
        src108 <= 12'h9fd;
        src109 <= 12'h63d;
        src110 <= 12'hbcd;
        src111 <= 12'he98;
        src112 <= 12'hfe4;
        src113 <= 12'h426;
        src114 <= 12'h44f;
        src115 <= 12'h8e;
        src116 <= 12'hec6;
        src117 <= 12'hd35;
        src118 <= 12'h9d8;
        src119 <= 12'ha68;
        src120 <= 12'h66;
        src121 <= 12'heaa;
        src122 <= 12'h367;
        src123 <= 12'hbe5;
        src124 <= 12'h935;
        src125 <= 12'hf46;
        src126 <= 12'h9f8;
        src127 <= 12'h5d5;
        src128 <= 12'h1fb;
        src129 <= 12'hc31;
        src130 <= 12'h2cd;
        src131 <= 12'h3fc;
        src132 <= 12'hf20;
        src133 <= 12'h419;
        src134 <= 12'hfe7;
        src135 <= 12'h67;
        src136 <= 12'h9b6;
        src137 <= 12'hfb9;
        src138 <= 12'h4fc;
        src139 <= 12'h733;
        src140 <= 12'hcb6;
        src141 <= 12'h325;
        src142 <= 12'h79c;
        src143 <= 12'hada;
        src144 <= 12'h65a;
        src145 <= 12'he2f;
        src146 <= 12'h221;
        src147 <= 12'hbc1;
        src148 <= 12'h891;
        src149 <= 12'h99c;
        src150 <= 12'h6a8;
        src151 <= 12'hb71;
        src152 <= 12'h7c9;
        src153 <= 12'hed5;
        src154 <= 12'h2a5;
        src155 <= 12'hbef;
        src156 <= 12'hcbb;
        src157 <= 12'haca;
        src158 <= 12'hf83;
        src159 <= 12'h1b4;
        src160 <= 12'h8c;
        src161 <= 12'h183;
        src162 <= 12'h563;
        src163 <= 12'h47f;
        src164 <= 12'h7fc;
        src165 <= 12'h4b6;
        src166 <= 12'h853;
        src167 <= 12'h7ad;
        src168 <= 12'h990;
        src169 <= 12'hbf;
        src170 <= 12'ha1d;
        src171 <= 12'h33b;
        src172 <= 12'h983;
        src173 <= 12'ha94;
        src174 <= 12'h8dc;
        src175 <= 12'hff5;
        src176 <= 12'h2f3;
        src177 <= 12'h9f8;
        src178 <= 12'hb13;
        src179 <= 12'hd63;
        src180 <= 12'hd8b;
        src181 <= 12'hebd;
        src182 <= 12'ha16;
        src183 <= 12'h47;
        src184 <= 12'hbe6;
        src185 <= 12'h1ba;
        src186 <= 12'h814;
        src187 <= 12'hc51;
        src188 <= 12'hed;
        exp <= 20'h66e41;
        #1
        src0 <= 12'h38;
        src1 <= 12'hb42;
        src2 <= 12'hd91;
        src3 <= 12'h7cc;
        src4 <= 12'h305;
        src5 <= 12'h49b;
        src6 <= 12'h34;
        src7 <= 12'h42a;
        src8 <= 12'h67f;
        src9 <= 12'h1a1;
        src10 <= 12'hf24;
        src11 <= 12'h22c;
        src12 <= 12'hd68;
        src13 <= 12'h690;
        src14 <= 12'h20e;
        src15 <= 12'ha7d;
        src16 <= 12'h1d3;
        src17 <= 12'hdf0;
        src18 <= 12'hece;
        src19 <= 12'hc2d;
        src20 <= 12'h2cd;
        src21 <= 12'h176;
        src22 <= 12'ha83;
        src23 <= 12'h4b9;
        src24 <= 12'hc81;
        src25 <= 12'hb34;
        src26 <= 12'h6c2;
        src27 <= 12'h73d;
        src28 <= 12'h137;
        src29 <= 12'h2b5;
        src30 <= 12'h9a2;
        src31 <= 12'h53f;
        src32 <= 12'hf22;
        src33 <= 12'h744;
        src34 <= 12'h4ed;
        src35 <= 12'hb44;
        src36 <= 12'h41;
        src37 <= 12'h51;
        src38 <= 12'heda;
        src39 <= 12'hf4;
        src40 <= 12'ha10;
        src41 <= 12'h567;
        src42 <= 12'h4b5;
        src43 <= 12'h780;
        src44 <= 12'h61b;
        src45 <= 12'h219;
        src46 <= 12'h9bc;
        src47 <= 12'h2a7;
        src48 <= 12'h69c;
        src49 <= 12'hb8c;
        src50 <= 12'h6ab;
        src51 <= 12'hade;
        src52 <= 12'h893;
        src53 <= 12'he60;
        src54 <= 12'h572;
        src55 <= 12'h4d5;
        src56 <= 12'hb0a;
        src57 <= 12'h622;
        src58 <= 12'h90c;
        src59 <= 12'ha2f;
        src60 <= 12'h8bb;
        src61 <= 12'hea1;
        src62 <= 12'h339;
        src63 <= 12'h852;
        src64 <= 12'h319;
        src65 <= 12'h2d2;
        src66 <= 12'h13a;
        src67 <= 12'h3b9;
        src68 <= 12'hf25;
        src69 <= 12'h88;
        src70 <= 12'hf4c;
        src71 <= 12'hc11;
        src72 <= 12'h199;
        src73 <= 12'h892;
        src74 <= 12'hd23;
        src75 <= 12'h296;
        src76 <= 12'he9e;
        src77 <= 12'hff7;
        src78 <= 12'h73b;
        src79 <= 12'hdc8;
        src80 <= 12'h216;
        src81 <= 12'ha4a;
        src82 <= 12'h1e8;
        src83 <= 12'h2c9;
        src84 <= 12'hdc1;
        src85 <= 12'hbd8;
        src86 <= 12'h61e;
        src87 <= 12'h26a;
        src88 <= 12'h304;
        src89 <= 12'h213;
        src90 <= 12'haed;
        src91 <= 12'h140;
        src92 <= 12'hf9;
        src93 <= 12'hc74;
        src94 <= 12'h521;
        src95 <= 12'he50;
        src96 <= 12'he85;
        src97 <= 12'hdf3;
        src98 <= 12'h88b;
        src99 <= 12'h399;
        src100 <= 12'h55;
        src101 <= 12'h571;
        src102 <= 12'hab8;
        src103 <= 12'h2;
        src104 <= 12'hdf7;
        src105 <= 12'hfcf;
        src106 <= 12'ha34;
        src107 <= 12'h91c;
        src108 <= 12'h120;
        src109 <= 12'h79f;
        src110 <= 12'hc7c;
        src111 <= 12'h4f1;
        src112 <= 12'hace;
        src113 <= 12'h109;
        src114 <= 12'h4f;
        src115 <= 12'h3af;
        src116 <= 12'heb;
        src117 <= 12'h43b;
        src118 <= 12'hd44;
        src119 <= 12'hb7c;
        src120 <= 12'h433;
        src121 <= 12'h432;
        src122 <= 12'h244;
        src123 <= 12'hb16;
        src124 <= 12'h5b;
        src125 <= 12'hdea;
        src126 <= 12'h762;
        src127 <= 12'he43;
        src128 <= 12'hb84;
        src129 <= 12'h937;
        src130 <= 12'h1e1;
        src131 <= 12'h49c;
        src132 <= 12'hc99;
        src133 <= 12'hf88;
        src134 <= 12'hd1;
        src135 <= 12'hdfb;
        src136 <= 12'h576;
        src137 <= 12'h22a;
        src138 <= 12'he7e;
        src139 <= 12'hd7b;
        src140 <= 12'h288;
        src141 <= 12'h50d;
        src142 <= 12'hd71;
        src143 <= 12'hf7e;
        src144 <= 12'h263;
        src145 <= 12'h7d5;
        src146 <= 12'h7f8;
        src147 <= 12'h91d;
        src148 <= 12'hd47;
        src149 <= 12'h7c4;
        src150 <= 12'hec8;
        src151 <= 12'hd96;
        src152 <= 12'h1ea;
        src153 <= 12'h4cc;
        src154 <= 12'h5e3;
        src155 <= 12'h269;
        src156 <= 12'hf28;
        src157 <= 12'hebf;
        src158 <= 12'h263;
        src159 <= 12'hc0e;
        src160 <= 12'h327;
        src161 <= 12'hb67;
        src162 <= 12'h6a6;
        src163 <= 12'hc59;
        src164 <= 12'hbb6;
        src165 <= 12'h410;
        src166 <= 12'h7d0;
        src167 <= 12'h2aa;
        src168 <= 12'hb2d;
        src169 <= 12'h3d9;
        src170 <= 12'h8ad;
        src171 <= 12'h19f;
        src172 <= 12'hdbf;
        src173 <= 12'h626;
        src174 <= 12'h549;
        src175 <= 12'h29c;
        src176 <= 12'hc0f;
        src177 <= 12'hc5e;
        src178 <= 12'h220;
        src179 <= 12'hb5e;
        src180 <= 12'h614;
        src181 <= 12'h62e;
        src182 <= 12'hb0;
        src183 <= 12'h7f8;
        src184 <= 12'h793;
        src185 <= 12'h219;
        src186 <= 12'h857;
        src187 <= 12'h6c7;
        src188 <= 12'hdec;
        exp <= 20'h58e39;
        #1
        src0 <= 12'h6ff;
        src1 <= 12'he21;
        src2 <= 12'h332;
        src3 <= 12'hd3d;
        src4 <= 12'hc2d;
        src5 <= 12'h33c;
        src6 <= 12'h8e0;
        src7 <= 12'h814;
        src8 <= 12'h12f;
        src9 <= 12'hdbc;
        src10 <= 12'h9ee;
        src11 <= 12'h68a;
        src12 <= 12'h492;
        src13 <= 12'hd61;
        src14 <= 12'hf14;
        src15 <= 12'h299;
        src16 <= 12'h76a;
        src17 <= 12'hc32;
        src18 <= 12'heb9;
        src19 <= 12'h171;
        src20 <= 12'h7cf;
        src21 <= 12'hfb8;
        src22 <= 12'h799;
        src23 <= 12'h34d;
        src24 <= 12'h934;
        src25 <= 12'h88b;
        src26 <= 12'h4ae;
        src27 <= 12'hc4d;
        src28 <= 12'hf70;
        src29 <= 12'he19;
        src30 <= 12'h26e;
        src31 <= 12'hcc5;
        src32 <= 12'h188;
        src33 <= 12'h145;
        src34 <= 12'h24e;
        src35 <= 12'h2d3;
        src36 <= 12'h881;
        src37 <= 12'h435;
        src38 <= 12'h6a3;
        src39 <= 12'h6b1;
        src40 <= 12'ha5d;
        src41 <= 12'ha83;
        src42 <= 12'hf85;
        src43 <= 12'h800;
        src44 <= 12'h861;
        src45 <= 12'h435;
        src46 <= 12'h8ef;
        src47 <= 12'h8ef;
        src48 <= 12'h94f;
        src49 <= 12'hfb1;
        src50 <= 12'h761;
        src51 <= 12'hd10;
        src52 <= 12'h54;
        src53 <= 12'ha9a;
        src54 <= 12'h4c;
        src55 <= 12'h7b;
        src56 <= 12'h84c;
        src57 <= 12'hff8;
        src58 <= 12'hcb9;
        src59 <= 12'hce8;
        src60 <= 12'h88c;
        src61 <= 12'h16e;
        src62 <= 12'hbcc;
        src63 <= 12'hfd;
        src64 <= 12'h8a1;
        src65 <= 12'h1b0;
        src66 <= 12'h777;
        src67 <= 12'h1ce;
        src68 <= 12'h3dc;
        src69 <= 12'h6c2;
        src70 <= 12'h581;
        src71 <= 12'hf;
        src72 <= 12'h591;
        src73 <= 12'haef;
        src74 <= 12'hdb1;
        src75 <= 12'h85c;
        src76 <= 12'hf4b;
        src77 <= 12'hc31;
        src78 <= 12'hab;
        src79 <= 12'h597;
        src80 <= 12'he56;
        src81 <= 12'hdaa;
        src82 <= 12'hdf3;
        src83 <= 12'h296;
        src84 <= 12'hed7;
        src85 <= 12'hcc6;
        src86 <= 12'h8d6;
        src87 <= 12'h3ab;
        src88 <= 12'hdf1;
        src89 <= 12'he7e;
        src90 <= 12'h7a0;
        src91 <= 12'h141;
        src92 <= 12'h9dc;
        src93 <= 12'h56d;
        src94 <= 12'h3d3;
        src95 <= 12'h336;
        src96 <= 12'h66e;
        src97 <= 12'ha07;
        src98 <= 12'h992;
        src99 <= 12'h741;
        src100 <= 12'he6e;
        src101 <= 12'h5a0;
        src102 <= 12'h95c;
        src103 <= 12'he22;
        src104 <= 12'h810;
        src105 <= 12'ha7d;
        src106 <= 12'h484;
        src107 <= 12'h1c3;
        src108 <= 12'hf02;
        src109 <= 12'h7cf;
        src110 <= 12'h22;
        src111 <= 12'hdf1;
        src112 <= 12'hd2e;
        src113 <= 12'h1ed;
        src114 <= 12'hacf;
        src115 <= 12'h701;
        src116 <= 12'he49;
        src117 <= 12'hdb;
        src118 <= 12'h40d;
        src119 <= 12'h221;
        src120 <= 12'hc97;
        src121 <= 12'h2e5;
        src122 <= 12'h1e3;
        src123 <= 12'h553;
        src124 <= 12'h76b;
        src125 <= 12'he87;
        src126 <= 12'h412;
        src127 <= 12'hac4;
        src128 <= 12'hc8b;
        src129 <= 12'h883;
        src130 <= 12'h519;
        src131 <= 12'he64;
        src132 <= 12'h981;
        src133 <= 12'h1ac;
        src134 <= 12'h53e;
        src135 <= 12'h5d0;
        src136 <= 12'ha23;
        src137 <= 12'h3d0;
        src138 <= 12'h16f;
        src139 <= 12'h290;
        src140 <= 12'he9f;
        src141 <= 12'h9dc;
        src142 <= 12'hd2f;
        src143 <= 12'h7fc;
        src144 <= 12'h706;
        src145 <= 12'ha0c;
        src146 <= 12'hada;
        src147 <= 12'h63b;
        src148 <= 12'h716;
        src149 <= 12'hc9a;
        src150 <= 12'hae2;
        src151 <= 12'hddf;
        src152 <= 12'h305;
        src153 <= 12'he17;
        src154 <= 12'hd3c;
        src155 <= 12'h895;
        src156 <= 12'h967;
        src157 <= 12'h8aa;
        src158 <= 12'h291;
        src159 <= 12'h406;
        src160 <= 12'he71;
        src161 <= 12'h4a;
        src162 <= 12'h9b8;
        src163 <= 12'h6df;
        src164 <= 12'h484;
        src165 <= 12'hcad;
        src166 <= 12'h2cc;
        src167 <= 12'hc8c;
        src168 <= 12'h8ee;
        src169 <= 12'ha17;
        src170 <= 12'hbce;
        src171 <= 12'h97f;
        src172 <= 12'hd9;
        src173 <= 12'hca3;
        src174 <= 12'h14f;
        src175 <= 12'h366;
        src176 <= 12'hb33;
        src177 <= 12'h2c1;
        src178 <= 12'h8e2;
        src179 <= 12'hf6c;
        src180 <= 12'h9af;
        src181 <= 12'hda2;
        src182 <= 12'h542;
        src183 <= 12'h240;
        src184 <= 12'hc40;
        src185 <= 12'h6a;
        src186 <= 12'h3c1;
        src187 <= 12'h87f;
        src188 <= 12'he8f;
        exp <= 20'h5f949;
        #1
        src0 <= 12'hb9f;
        src1 <= 12'ha9d;
        src2 <= 12'ha40;
        src3 <= 12'ha6b;
        src4 <= 12'hf50;
        src5 <= 12'h10f;
        src6 <= 12'hd25;
        src7 <= 12'hef6;
        src8 <= 12'h400;
        src9 <= 12'h21a;
        src10 <= 12'h8b6;
        src11 <= 12'h740;
        src12 <= 12'h95;
        src13 <= 12'h1c9;
        src14 <= 12'h536;
        src15 <= 12'hf68;
        src16 <= 12'haba;
        src17 <= 12'hd2b;
        src18 <= 12'h229;
        src19 <= 12'hf69;
        src20 <= 12'h316;
        src21 <= 12'h723;
        src22 <= 12'hb0b;
        src23 <= 12'ha84;
        src24 <= 12'h740;
        src25 <= 12'h18d;
        src26 <= 12'h8;
        src27 <= 12'h6e9;
        src28 <= 12'h65;
        src29 <= 12'h4e4;
        src30 <= 12'h702;
        src31 <= 12'h372;
        src32 <= 12'h228;
        src33 <= 12'h8a7;
        src34 <= 12'hbae;
        src35 <= 12'hbf5;
        src36 <= 12'h4fb;
        src37 <= 12'h840;
        src38 <= 12'he21;
        src39 <= 12'h260;
        src40 <= 12'hd6a;
        src41 <= 12'h92e;
        src42 <= 12'h2c8;
        src43 <= 12'hd39;
        src44 <= 12'h4c1;
        src45 <= 12'h6d8;
        src46 <= 12'h0;
        src47 <= 12'h28d;
        src48 <= 12'h25f;
        src49 <= 12'h2c3;
        src50 <= 12'hc77;
        src51 <= 12'ha6;
        src52 <= 12'hfe1;
        src53 <= 12'hf55;
        src54 <= 12'hc49;
        src55 <= 12'h367;
        src56 <= 12'h505;
        src57 <= 12'h964;
        src58 <= 12'hf54;
        src59 <= 12'hb3f;
        src60 <= 12'hb1c;
        src61 <= 12'hbcd;
        src62 <= 12'hb5b;
        src63 <= 12'h33d;
        src64 <= 12'h5ba;
        src65 <= 12'h737;
        src66 <= 12'hc89;
        src67 <= 12'h824;
        src68 <= 12'h9fd;
        src69 <= 12'h4da;
        src70 <= 12'h2bb;
        src71 <= 12'h46d;
        src72 <= 12'ha05;
        src73 <= 12'h322;
        src74 <= 12'h352;
        src75 <= 12'hf83;
        src76 <= 12'h4ed;
        src77 <= 12'h467;
        src78 <= 12'h216;
        src79 <= 12'h6e1;
        src80 <= 12'h3db;
        src81 <= 12'h688;
        src82 <= 12'h2e5;
        src83 <= 12'h560;
        src84 <= 12'h50c;
        src85 <= 12'h5ba;
        src86 <= 12'hb3;
        src87 <= 12'h226;
        src88 <= 12'h245;
        src89 <= 12'had4;
        src90 <= 12'h5ad;
        src91 <= 12'h45d;
        src92 <= 12'h180;
        src93 <= 12'h80;
        src94 <= 12'h533;
        src95 <= 12'hed8;
        src96 <= 12'h3fc;
        src97 <= 12'h5d;
        src98 <= 12'h9e2;
        src99 <= 12'hf98;
        src100 <= 12'h914;
        src101 <= 12'hb35;
        src102 <= 12'hfd2;
        src103 <= 12'h942;
        src104 <= 12'h521;
        src105 <= 12'h7ee;
        src106 <= 12'hced;
        src107 <= 12'h31b;
        src108 <= 12'hbe1;
        src109 <= 12'h595;
        src110 <= 12'h89;
        src111 <= 12'hfbd;
        src112 <= 12'h189;
        src113 <= 12'h5f0;
        src114 <= 12'hb2;
        src115 <= 12'hbb;
        src116 <= 12'hdab;
        src117 <= 12'hfd6;
        src118 <= 12'h82;
        src119 <= 12'h93f;
        src120 <= 12'h6ee;
        src121 <= 12'h75c;
        src122 <= 12'h85;
        src123 <= 12'h326;
        src124 <= 12'hc61;
        src125 <= 12'hda2;
        src126 <= 12'h523;
        src127 <= 12'h15e;
        src128 <= 12'h462;
        src129 <= 12'h723;
        src130 <= 12'he84;
        src131 <= 12'hc19;
        src132 <= 12'h775;
        src133 <= 12'hf11;
        src134 <= 12'h2cd;
        src135 <= 12'hafe;
        src136 <= 12'he0f;
        src137 <= 12'h36a;
        src138 <= 12'hac5;
        src139 <= 12'h932;
        src140 <= 12'hf73;
        src141 <= 12'h3e1;
        src142 <= 12'h215;
        src143 <= 12'h798;
        src144 <= 12'hd1d;
        src145 <= 12'hda4;
        src146 <= 12'hc2e;
        src147 <= 12'he55;
        src148 <= 12'hc2a;
        src149 <= 12'hc58;
        src150 <= 12'h76a;
        src151 <= 12'hea3;
        src152 <= 12'h353;
        src153 <= 12'hc50;
        src154 <= 12'h67d;
        src155 <= 12'h567;
        src156 <= 12'hc39;
        src157 <= 12'h6c3;
        src158 <= 12'h525;
        src159 <= 12'h746;
        src160 <= 12'hdfc;
        src161 <= 12'hba3;
        src162 <= 12'h7f0;
        src163 <= 12'hc41;
        src164 <= 12'hb58;
        src165 <= 12'h7f;
        src166 <= 12'h856;
        src167 <= 12'hf13;
        src168 <= 12'h2d9;
        src169 <= 12'h366;
        src170 <= 12'h232;
        src171 <= 12'h2ce;
        src172 <= 12'ha36;
        src173 <= 12'h5fb;
        src174 <= 12'h7b5;
        src175 <= 12'h651;
        src176 <= 12'h5ed;
        src177 <= 12'h489;
        src178 <= 12'hef1;
        src179 <= 12'h93b;
        src180 <= 12'hf6;
        src181 <= 12'ha3e;
        src182 <= 12'h2d7;
        src183 <= 12'h1a2;
        src184 <= 12'h309;
        src185 <= 12'h486;
        src186 <= 12'h803;
        src187 <= 12'hea3;
        src188 <= 12'h5e7;
        exp <= 20'h59249;
        #1
        src0 <= 12'h699;
        src1 <= 12'hb8;
        src2 <= 12'h530;
        src3 <= 12'ha12;
        src4 <= 12'h2cf;
        src5 <= 12'hdf2;
        src6 <= 12'hef2;
        src7 <= 12'hdbf;
        src8 <= 12'h50b;
        src9 <= 12'h6ba;
        src10 <= 12'h687;
        src11 <= 12'h226;
        src12 <= 12'h81d;
        src13 <= 12'hb2d;
        src14 <= 12'hd3d;
        src15 <= 12'hbe8;
        src16 <= 12'ha58;
        src17 <= 12'h5d0;
        src18 <= 12'h4ec;
        src19 <= 12'hffe;
        src20 <= 12'h975;
        src21 <= 12'ha85;
        src22 <= 12'hf18;
        src23 <= 12'h40b;
        src24 <= 12'hd41;
        src25 <= 12'h128;
        src26 <= 12'h91f;
        src27 <= 12'h79b;
        src28 <= 12'h6de;
        src29 <= 12'h3de;
        src30 <= 12'h1e7;
        src31 <= 12'h56d;
        src32 <= 12'hb34;
        src33 <= 12'h7c9;
        src34 <= 12'h7fb;
        src35 <= 12'h831;
        src36 <= 12'h8ca;
        src37 <= 12'hde5;
        src38 <= 12'h4d3;
        src39 <= 12'ha6;
        src40 <= 12'ha8;
        src41 <= 12'hc76;
        src42 <= 12'hb2b;
        src43 <= 12'h188;
        src44 <= 12'he4d;
        src45 <= 12'h4dd;
        src46 <= 12'h5e7;
        src47 <= 12'ha00;
        src48 <= 12'h146;
        src49 <= 12'h19e;
        src50 <= 12'h989;
        src51 <= 12'hfec;
        src52 <= 12'hb6d;
        src53 <= 12'h2a0;
        src54 <= 12'hc76;
        src55 <= 12'h5a9;
        src56 <= 12'h97d;
        src57 <= 12'hb95;
        src58 <= 12'h987;
        src59 <= 12'h5bf;
        src60 <= 12'h297;
        src61 <= 12'h5ed;
        src62 <= 12'h29d;
        src63 <= 12'hff0;
        src64 <= 12'hc65;
        src65 <= 12'hab8;
        src66 <= 12'h715;
        src67 <= 12'h59;
        src68 <= 12'hfaa;
        src69 <= 12'hb3;
        src70 <= 12'h6bc;
        src71 <= 12'h4b;
        src72 <= 12'h9dc;
        src73 <= 12'hc72;
        src74 <= 12'h4a3;
        src75 <= 12'hf54;
        src76 <= 12'h558;
        src77 <= 12'h666;
        src78 <= 12'ha7;
        src79 <= 12'hdd3;
        src80 <= 12'h2cc;
        src81 <= 12'h710;
        src82 <= 12'h3ac;
        src83 <= 12'hca4;
        src84 <= 12'ha5a;
        src85 <= 12'hed5;
        src86 <= 12'h2ac;
        src87 <= 12'he80;
        src88 <= 12'h2be;
        src89 <= 12'h975;
        src90 <= 12'hdc8;
        src91 <= 12'h7f3;
        src92 <= 12'h38a;
        src93 <= 12'h6ce;
        src94 <= 12'hd71;
        src95 <= 12'h66f;
        src96 <= 12'h988;
        src97 <= 12'hb7b;
        src98 <= 12'he24;
        src99 <= 12'h2f0;
        src100 <= 12'hba1;
        src101 <= 12'h7a1;
        src102 <= 12'h51b;
        src103 <= 12'h114;
        src104 <= 12'hd64;
        src105 <= 12'h8c1;
        src106 <= 12'hff1;
        src107 <= 12'h5bc;
        src108 <= 12'hcc1;
        src109 <= 12'h6b4;
        src110 <= 12'h9b2;
        src111 <= 12'h2ab;
        src112 <= 12'habc;
        src113 <= 12'he95;
        src114 <= 12'ha0b;
        src115 <= 12'h4a5;
        src116 <= 12'h6c5;
        src117 <= 12'h5fc;
        src118 <= 12'h7d4;
        src119 <= 12'h6b8;
        src120 <= 12'h539;
        src121 <= 12'h68d;
        src122 <= 12'h116;
        src123 <= 12'h8d0;
        src124 <= 12'hb87;
        src125 <= 12'he42;
        src126 <= 12'h5d2;
        src127 <= 12'ha;
        src128 <= 12'h907;
        src129 <= 12'h54d;
        src130 <= 12'hb82;
        src131 <= 12'h865;
        src132 <= 12'h334;
        src133 <= 12'h93d;
        src134 <= 12'h841;
        src135 <= 12'hb13;
        src136 <= 12'h977;
        src137 <= 12'hfc;
        src138 <= 12'h666;
        src139 <= 12'h571;
        src140 <= 12'h199;
        src141 <= 12'h3fc;
        src142 <= 12'hb7a;
        src143 <= 12'hb3a;
        src144 <= 12'h3ae;
        src145 <= 12'hde7;
        src146 <= 12'h847;
        src147 <= 12'h7ec;
        src148 <= 12'h5d2;
        src149 <= 12'h854;
        src150 <= 12'ha5a;
        src151 <= 12'hcd2;
        src152 <= 12'haea;
        src153 <= 12'hb58;
        src154 <= 12'h4d2;
        src155 <= 12'h828;
        src156 <= 12'h7d4;
        src157 <= 12'hc7f;
        src158 <= 12'ha3c;
        src159 <= 12'h472;
        src160 <= 12'hb7a;
        src161 <= 12'h3c1;
        src162 <= 12'h769;
        src163 <= 12'h541;
        src164 <= 12'h23b;
        src165 <= 12'h2b7;
        src166 <= 12'h960;
        src167 <= 12'h7a2;
        src168 <= 12'h51e;
        src169 <= 12'h1c7;
        src170 <= 12'h4dd;
        src171 <= 12'h64b;
        src172 <= 12'h605;
        src173 <= 12'hb55;
        src174 <= 12'h5fb;
        src175 <= 12'h33;
        src176 <= 12'h2a5;
        src177 <= 12'ha75;
        src178 <= 12'h1c9;
        src179 <= 12'h5fc;
        src180 <= 12'h4ce;
        src181 <= 12'hac2;
        src182 <= 12'hc4c;
        src183 <= 12'h498;
        src184 <= 12'h68d;
        src185 <= 12'h405;
        src186 <= 12'h23f;
        src187 <= 12'hbe0;
        src188 <= 12'hd3c;
        exp <= 20'h5b5e5;
        #1
        src0 <= 12'hb7a;
        src1 <= 12'h1b0;
        src2 <= 12'h9b5;
        src3 <= 12'ha81;
        src4 <= 12'h6de;
        src5 <= 12'h57d;
        src6 <= 12'h559;
        src7 <= 12'h38a;
        src8 <= 12'h1f3;
        src9 <= 12'ha8f;
        src10 <= 12'hc89;
        src11 <= 12'h849;
        src12 <= 12'he0c;
        src13 <= 12'h688;
        src14 <= 12'hd3d;
        src15 <= 12'h8ae;
        src16 <= 12'h811;
        src17 <= 12'hff6;
        src18 <= 12'h241;
        src19 <= 12'hddb;
        src20 <= 12'h4ae;
        src21 <= 12'h163;
        src22 <= 12'h4c7;
        src23 <= 12'h5da;
        src24 <= 12'hbe6;
        src25 <= 12'h987;
        src26 <= 12'h579;
        src27 <= 12'h119;
        src28 <= 12'hb14;
        src29 <= 12'hfc4;
        src30 <= 12'h765;
        src31 <= 12'haf9;
        src32 <= 12'h510;
        src33 <= 12'h68f;
        src34 <= 12'hdd2;
        src35 <= 12'h91a;
        src36 <= 12'hfbf;
        src37 <= 12'hffc;
        src38 <= 12'hb6c;
        src39 <= 12'h846;
        src40 <= 12'hf5f;
        src41 <= 12'h60c;
        src42 <= 12'h894;
        src43 <= 12'haec;
        src44 <= 12'h40;
        src45 <= 12'hebc;
        src46 <= 12'h986;
        src47 <= 12'h19;
        src48 <= 12'h8f4;
        src49 <= 12'h617;
        src50 <= 12'h57d;
        src51 <= 12'hc1b;
        src52 <= 12'h2a9;
        src53 <= 12'hfcb;
        src54 <= 12'h800;
        src55 <= 12'h932;
        src56 <= 12'h45f;
        src57 <= 12'hb79;
        src58 <= 12'he52;
        src59 <= 12'h1e3;
        src60 <= 12'h3a7;
        src61 <= 12'hac6;
        src62 <= 12'h66a;
        src63 <= 12'hbf2;
        src64 <= 12'h440;
        src65 <= 12'ha37;
        src66 <= 12'hda7;
        src67 <= 12'hb0b;
        src68 <= 12'h106;
        src69 <= 12'hb07;
        src70 <= 12'h795;
        src71 <= 12'hb74;
        src72 <= 12'hc37;
        src73 <= 12'h897;
        src74 <= 12'h8d0;
        src75 <= 12'h944;
        src76 <= 12'h761;
        src77 <= 12'hc7b;
        src78 <= 12'hc77;
        src79 <= 12'h1b5;
        src80 <= 12'h1a9;
        src81 <= 12'h375;
        src82 <= 12'h334;
        src83 <= 12'hef1;
        src84 <= 12'h4d1;
        src85 <= 12'h640;
        src86 <= 12'h838;
        src87 <= 12'hea0;
        src88 <= 12'h55f;
        src89 <= 12'h286;
        src90 <= 12'h2b;
        src91 <= 12'h80a;
        src92 <= 12'h1fb;
        src93 <= 12'h116;
        src94 <= 12'h4dd;
        src95 <= 12'h6;
        src96 <= 12'h94d;
        src97 <= 12'h2da;
        src98 <= 12'h464;
        src99 <= 12'h29b;
        src100 <= 12'h51a;
        src101 <= 12'hc2c;
        src102 <= 12'hb35;
        src103 <= 12'hcdd;
        src104 <= 12'hebd;
        src105 <= 12'hc10;
        src106 <= 12'h6b2;
        src107 <= 12'h6ed;
        src108 <= 12'ha28;
        src109 <= 12'h99d;
        src110 <= 12'hc88;
        src111 <= 12'h45a;
        src112 <= 12'h118;
        src113 <= 12'h890;
        src114 <= 12'hdde;
        src115 <= 12'h9a;
        src116 <= 12'hf22;
        src117 <= 12'ha4f;
        src118 <= 12'h38c;
        src119 <= 12'h1f9;
        src120 <= 12'h244;
        src121 <= 12'h74;
        src122 <= 12'h3c0;
        src123 <= 12'hafc;
        src124 <= 12'h269;
        src125 <= 12'h4c1;
        src126 <= 12'h840;
        src127 <= 12'he69;
        src128 <= 12'h605;
        src129 <= 12'h784;
        src130 <= 12'hd61;
        src131 <= 12'haa6;
        src132 <= 12'ha25;
        src133 <= 12'h837;
        src134 <= 12'he08;
        src135 <= 12'h577;
        src136 <= 12'h55b;
        src137 <= 12'hfd1;
        src138 <= 12'he1c;
        src139 <= 12'h7d5;
        src140 <= 12'h96b;
        src141 <= 12'h873;
        src142 <= 12'h513;
        src143 <= 12'h95c;
        src144 <= 12'h9df;
        src145 <= 12'ha8b;
        src146 <= 12'h45f;
        src147 <= 12'h55c;
        src148 <= 12'h2af;
        src149 <= 12'ha3b;
        src150 <= 12'h4c5;
        src151 <= 12'h80f;
        src152 <= 12'hbc4;
        src153 <= 12'h275;
        src154 <= 12'h284;
        src155 <= 12'h420;
        src156 <= 12'h357;
        src157 <= 12'ha8;
        src158 <= 12'hee;
        src159 <= 12'he;
        src160 <= 12'hb0d;
        src161 <= 12'h7e9;
        src162 <= 12'h4f0;
        src163 <= 12'h186;
        src164 <= 12'hf17;
        src165 <= 12'hda6;
        src166 <= 12'hca9;
        src167 <= 12'h4a8;
        src168 <= 12'hdd8;
        src169 <= 12'h761;
        src170 <= 12'h36;
        src171 <= 12'h16;
        src172 <= 12'h53;
        src173 <= 12'he49;
        src174 <= 12'he1b;
        src175 <= 12'h247;
        src176 <= 12'hc06;
        src177 <= 12'hdc9;
        src178 <= 12'hbaf;
        src179 <= 12'ha6a;
        src180 <= 12'h2c;
        src181 <= 12'hf18;
        src182 <= 12'h797;
        src183 <= 12'hcb2;
        src184 <= 12'hcb7;
        src185 <= 12'haba;
        src186 <= 12'ha02;
        src187 <= 12'he48;
        src188 <= 12'h9fe;
        exp <= 20'h5e324;
        #1
        src0 <= 12'h3f2;
        src1 <= 12'h43c;
        src2 <= 12'hebc;
        src3 <= 12'h80e;
        src4 <= 12'haba;
        src5 <= 12'h1e7;
        src6 <= 12'he2;
        src7 <= 12'h1ec;
        src8 <= 12'h1ff;
        src9 <= 12'heb3;
        src10 <= 12'h884;
        src11 <= 12'h205;
        src12 <= 12'h4b4;
        src13 <= 12'h5bb;
        src14 <= 12'h834;
        src15 <= 12'h242;
        src16 <= 12'h867;
        src17 <= 12'h6a0;
        src18 <= 12'hba9;
        src19 <= 12'h740;
        src20 <= 12'h58b;
        src21 <= 12'h977;
        src22 <= 12'h405;
        src23 <= 12'hfd;
        src24 <= 12'h7b;
        src25 <= 12'he7;
        src26 <= 12'hf0f;
        src27 <= 12'he3e;
        src28 <= 12'h998;
        src29 <= 12'hf67;
        src30 <= 12'h8ed;
        src31 <= 12'h796;
        src32 <= 12'hcf9;
        src33 <= 12'h781;
        src34 <= 12'h705;
        src35 <= 12'hf4e;
        src36 <= 12'h36b;
        src37 <= 12'hf96;
        src38 <= 12'h3a4;
        src39 <= 12'h1eb;
        src40 <= 12'h237;
        src41 <= 12'h14b;
        src42 <= 12'hbe5;
        src43 <= 12'h818;
        src44 <= 12'h1bd;
        src45 <= 12'h5ca;
        src46 <= 12'h857;
        src47 <= 12'h4e8;
        src48 <= 12'h86b;
        src49 <= 12'he03;
        src50 <= 12'h632;
        src51 <= 12'hd90;
        src52 <= 12'hbe5;
        src53 <= 12'h91f;
        src54 <= 12'h595;
        src55 <= 12'ha42;
        src56 <= 12'h394;
        src57 <= 12'h186;
        src58 <= 12'h186;
        src59 <= 12'h23a;
        src60 <= 12'hc9e;
        src61 <= 12'h699;
        src62 <= 12'h931;
        src63 <= 12'hd5a;
        src64 <= 12'h352;
        src65 <= 12'h926;
        src66 <= 12'h10c;
        src67 <= 12'he77;
        src68 <= 12'hce0;
        src69 <= 12'heab;
        src70 <= 12'hbaf;
        src71 <= 12'hf6e;
        src72 <= 12'hd8a;
        src73 <= 12'h33;
        src74 <= 12'h313;
        src75 <= 12'h6be;
        src76 <= 12'h77b;
        src77 <= 12'hc0d;
        src78 <= 12'hb2e;
        src79 <= 12'hab2;
        src80 <= 12'hde8;
        src81 <= 12'h7e6;
        src82 <= 12'hc8;
        src83 <= 12'h6aa;
        src84 <= 12'hbb;
        src85 <= 12'h847;
        src86 <= 12'haf0;
        src87 <= 12'hc5;
        src88 <= 12'h2f1;
        src89 <= 12'hc70;
        src90 <= 12'h3aa;
        src91 <= 12'ha0c;
        src92 <= 12'h27b;
        src93 <= 12'hdce;
        src94 <= 12'h8d0;
        src95 <= 12'hfd1;
        src96 <= 12'h8c2;
        src97 <= 12'h233;
        src98 <= 12'hba3;
        src99 <= 12'h4fd;
        src100 <= 12'h88a;
        src101 <= 12'ha4d;
        src102 <= 12'h71e;
        src103 <= 12'he9c;
        src104 <= 12'hd;
        src105 <= 12'h7af;
        src106 <= 12'h561;
        src107 <= 12'hef1;
        src108 <= 12'hc50;
        src109 <= 12'h23a;
        src110 <= 12'h89f;
        src111 <= 12'hc1c;
        src112 <= 12'h2f;
        src113 <= 12'h236;
        src114 <= 12'h89e;
        src115 <= 12'hc45;
        src116 <= 12'h815;
        src117 <= 12'h66d;
        src118 <= 12'ha5;
        src119 <= 12'hf7;
        src120 <= 12'h7a9;
        src121 <= 12'ha17;
        src122 <= 12'h75b;
        src123 <= 12'h8ab;
        src124 <= 12'he5e;
        src125 <= 12'h932;
        src126 <= 12'hf73;
        src127 <= 12'hbb0;
        src128 <= 12'h8a5;
        src129 <= 12'he3f;
        src130 <= 12'h9b4;
        src131 <= 12'h6f2;
        src132 <= 12'hd32;
        src133 <= 12'haa0;
        src134 <= 12'h84f;
        src135 <= 12'h5f3;
        src136 <= 12'h4ee;
        src137 <= 12'hbdd;
        src138 <= 12'hf75;
        src139 <= 12'h1;
        src140 <= 12'h661;
        src141 <= 12'h6c3;
        src142 <= 12'h56b;
        src143 <= 12'hfab;
        src144 <= 12'hf9d;
        src145 <= 12'h8bf;
        src146 <= 12'hff;
        src147 <= 12'h24;
        src148 <= 12'hb0;
        src149 <= 12'h263;
        src150 <= 12'ha64;
        src151 <= 12'hb46;
        src152 <= 12'hb79;
        src153 <= 12'hfd9;
        src154 <= 12'hf0b;
        src155 <= 12'h90a;
        src156 <= 12'hed5;
        src157 <= 12'h227;
        src158 <= 12'h960;
        src159 <= 12'hebf;
        src160 <= 12'hfea;
        src161 <= 12'h504;
        src162 <= 12'h19a;
        src163 <= 12'he68;
        src164 <= 12'hd1d;
        src165 <= 12'h997;
        src166 <= 12'h35a;
        src167 <= 12'ha04;
        src168 <= 12'h89;
        src169 <= 12'h99d;
        src170 <= 12'h148;
        src171 <= 12'hff0;
        src172 <= 12'h1b5;
        src173 <= 12'h2d3;
        src174 <= 12'hb62;
        src175 <= 12'h1d8;
        src176 <= 12'h6c2;
        src177 <= 12'hd7b;
        src178 <= 12'h69d;
        src179 <= 12'h988;
        src180 <= 12'hda1;
        src181 <= 12'ha09;
        src182 <= 12'h986;
        src183 <= 12'h757;
        src184 <= 12'h9a1;
        src185 <= 12'h2be;
        src186 <= 12'ha4f;
        src187 <= 12'h33c;
        src188 <= 12'h9e5;
        exp <= 20'h5de8f;
        #1
        src0 <= 12'h762;
        src1 <= 12'h6e1;
        src2 <= 12'h752;
        src3 <= 12'h72d;
        src4 <= 12'h599;
        src5 <= 12'h316;
        src6 <= 12'h96f;
        src7 <= 12'h43b;
        src8 <= 12'hef1;
        src9 <= 12'h725;
        src10 <= 12'hc74;
        src11 <= 12'hbbc;
        src12 <= 12'h1db;
        src13 <= 12'h56f;
        src14 <= 12'hf5d;
        src15 <= 12'h37c;
        src16 <= 12'h982;
        src17 <= 12'h492;
        src18 <= 12'h4d4;
        src19 <= 12'h388;
        src20 <= 12'hb02;
        src21 <= 12'h65b;
        src22 <= 12'h1be;
        src23 <= 12'hfea;
        src24 <= 12'ha82;
        src25 <= 12'h903;
        src26 <= 12'h1c4;
        src27 <= 12'hd33;
        src28 <= 12'h9f;
        src29 <= 12'hfb;
        src30 <= 12'h89e;
        src31 <= 12'hd53;
        src32 <= 12'h629;
        src33 <= 12'h19a;
        src34 <= 12'hdd3;
        src35 <= 12'haf6;
        src36 <= 12'h8e8;
        src37 <= 12'h395;
        src38 <= 12'h499;
        src39 <= 12'hab9;
        src40 <= 12'h97a;
        src41 <= 12'h61b;
        src42 <= 12'h7e;
        src43 <= 12'h58e;
        src44 <= 12'hb1b;
        src45 <= 12'h7e4;
        src46 <= 12'h914;
        src47 <= 12'h4b;
        src48 <= 12'haeb;
        src49 <= 12'h307;
        src50 <= 12'h361;
        src51 <= 12'hc9a;
        src52 <= 12'hd3e;
        src53 <= 12'hc;
        src54 <= 12'h725;
        src55 <= 12'h41f;
        src56 <= 12'hd5;
        src57 <= 12'h321;
        src58 <= 12'heda;
        src59 <= 12'h50b;
        src60 <= 12'h120;
        src61 <= 12'h983;
        src62 <= 12'h2c3;
        src63 <= 12'h40f;
        src64 <= 12'hb61;
        src65 <= 12'h6b1;
        src66 <= 12'h51f;
        src67 <= 12'h6e3;
        src68 <= 12'h9a9;
        src69 <= 12'hc07;
        src70 <= 12'he06;
        src71 <= 12'h5fe;
        src72 <= 12'h9f8;
        src73 <= 12'h4fb;
        src74 <= 12'h80c;
        src75 <= 12'ha7a;
        src76 <= 12'h13c;
        src77 <= 12'h3d2;
        src78 <= 12'hb36;
        src79 <= 12'h8b7;
        src80 <= 12'hfce;
        src81 <= 12'h744;
        src82 <= 12'h69d;
        src83 <= 12'h5ea;
        src84 <= 12'h62a;
        src85 <= 12'h4b0;
        src86 <= 12'h235;
        src87 <= 12'h1e8;
        src88 <= 12'hbbd;
        src89 <= 12'he3;
        src90 <= 12'h2a6;
        src91 <= 12'haa9;
        src92 <= 12'hba8;
        src93 <= 12'h49a;
        src94 <= 12'hd7a;
        src95 <= 12'hf1c;
        src96 <= 12'he47;
        src97 <= 12'h84f;
        src98 <= 12'h7c7;
        src99 <= 12'h9b4;
        src100 <= 12'h4bc;
        src101 <= 12'h3a1;
        src102 <= 12'hf72;
        src103 <= 12'he87;
        src104 <= 12'hae0;
        src105 <= 12'h45d;
        src106 <= 12'h28;
        src107 <= 12'h363;
        src108 <= 12'hd93;
        src109 <= 12'h305;
        src110 <= 12'h935;
        src111 <= 12'h8eb;
        src112 <= 12'h48;
        src113 <= 12'h6f8;
        src114 <= 12'h5f2;
        src115 <= 12'h4f5;
        src116 <= 12'he2;
        src117 <= 12'ha7d;
        src118 <= 12'hdc7;
        src119 <= 12'hef6;
        src120 <= 12'he1f;
        src121 <= 12'h3aa;
        src122 <= 12'hf5c;
        src123 <= 12'h657;
        src124 <= 12'h651;
        src125 <= 12'hcc6;
        src126 <= 12'hedd;
        src127 <= 12'h278;
        src128 <= 12'hbfc;
        src129 <= 12'h47f;
        src130 <= 12'he18;
        src131 <= 12'he62;
        src132 <= 12'h19f;
        src133 <= 12'h15a;
        src134 <= 12'hd17;
        src135 <= 12'h15;
        src136 <= 12'hc94;
        src137 <= 12'hd6e;
        src138 <= 12'hcb1;
        src139 <= 12'hf91;
        src140 <= 12'ha69;
        src141 <= 12'hb24;
        src142 <= 12'haef;
        src143 <= 12'h767;
        src144 <= 12'hbf8;
        src145 <= 12'h116;
        src146 <= 12'hdbe;
        src147 <= 12'hd0e;
        src148 <= 12'hfd2;
        src149 <= 12'he44;
        src150 <= 12'ha85;
        src151 <= 12'h6ef;
        src152 <= 12'h4fa;
        src153 <= 12'hdb0;
        src154 <= 12'h29f;
        src155 <= 12'h351;
        src156 <= 12'hb8b;
        src157 <= 12'hf8c;
        src158 <= 12'hb8f;
        src159 <= 12'h713;
        src160 <= 12'h12f;
        src161 <= 12'h3e8;
        src162 <= 12'h374;
        src163 <= 12'hf47;
        src164 <= 12'h8fb;
        src165 <= 12'h96a;
        src166 <= 12'h9bc;
        src167 <= 12'hb1c;
        src168 <= 12'h369;
        src169 <= 12'h319;
        src170 <= 12'h7b;
        src171 <= 12'he9d;
        src172 <= 12'h633;
        src173 <= 12'h94b;
        src174 <= 12'h59b;
        src175 <= 12'h7a2;
        src176 <= 12'h6b;
        src177 <= 12'hbcb;
        src178 <= 12'h8d8;
        src179 <= 12'h910;
        src180 <= 12'hed1;
        src181 <= 12'h3f;
        src182 <= 12'hf6f;
        src183 <= 12'h42;
        src184 <= 12'h1b7;
        src185 <= 12'he47;
        src186 <= 12'h1e8;
        src187 <= 12'h4b3;
        src188 <= 12'h2f7;
        exp <= 20'h5c395;
        #1
        src0 <= 12'hae7;
        src1 <= 12'h52b;
        src2 <= 12'hcaa;
        src3 <= 12'hcde;
        src4 <= 12'hf3b;
        src5 <= 12'h148;
        src6 <= 12'h85a;
        src7 <= 12'hcba;
        src8 <= 12'h8df;
        src9 <= 12'h5f9;
        src10 <= 12'h377;
        src11 <= 12'hb34;
        src12 <= 12'h272;
        src13 <= 12'h18a;
        src14 <= 12'h449;
        src15 <= 12'h4db;
        src16 <= 12'h1a6;
        src17 <= 12'h579;
        src18 <= 12'h645;
        src19 <= 12'he92;
        src20 <= 12'h38d;
        src21 <= 12'h147;
        src22 <= 12'hc67;
        src23 <= 12'hf55;
        src24 <= 12'hd0e;
        src25 <= 12'h82b;
        src26 <= 12'h21c;
        src27 <= 12'h93b;
        src28 <= 12'h6ce;
        src29 <= 12'hbea;
        src30 <= 12'haf6;
        src31 <= 12'h8d8;
        src32 <= 12'hdd1;
        src33 <= 12'h87e;
        src34 <= 12'ha44;
        src35 <= 12'hb2e;
        src36 <= 12'h582;
        src37 <= 12'h68f;
        src38 <= 12'hae0;
        src39 <= 12'ha64;
        src40 <= 12'h15e;
        src41 <= 12'h7c9;
        src42 <= 12'h562;
        src43 <= 12'h40b;
        src44 <= 12'h488;
        src45 <= 12'h92e;
        src46 <= 12'h69f;
        src47 <= 12'hd43;
        src48 <= 12'h788;
        src49 <= 12'h2f6;
        src50 <= 12'h7ce;
        src51 <= 12'hd92;
        src52 <= 12'h924;
        src53 <= 12'h303;
        src54 <= 12'h117;
        src55 <= 12'h7d0;
        src56 <= 12'h6b3;
        src57 <= 12'h63e;
        src58 <= 12'h583;
        src59 <= 12'hf21;
        src60 <= 12'h270;
        src61 <= 12'hd4e;
        src62 <= 12'hd4c;
        src63 <= 12'h7d7;
        src64 <= 12'hf0;
        src65 <= 12'h8b;
        src66 <= 12'h6b9;
        src67 <= 12'hc10;
        src68 <= 12'h290;
        src69 <= 12'h5c2;
        src70 <= 12'he70;
        src71 <= 12'h9f8;
        src72 <= 12'hd53;
        src73 <= 12'h9c1;
        src74 <= 12'hf14;
        src75 <= 12'h5ce;
        src76 <= 12'h276;
        src77 <= 12'h973;
        src78 <= 12'h522;
        src79 <= 12'hf39;
        src80 <= 12'h38f;
        src81 <= 12'hd11;
        src82 <= 12'h6f8;
        src83 <= 12'hebd;
        src84 <= 12'h6ba;
        src85 <= 12'h5b;
        src86 <= 12'hd02;
        src87 <= 12'h29;
        src88 <= 12'h1b1;
        src89 <= 12'hcb5;
        src90 <= 12'hb75;
        src91 <= 12'hca0;
        src92 <= 12'hff9;
        src93 <= 12'hb7a;
        src94 <= 12'hcc7;
        src95 <= 12'h488;
        src96 <= 12'ha05;
        src97 <= 12'h4ce;
        src98 <= 12'hdfe;
        src99 <= 12'h1c1;
        src100 <= 12'h177;
        src101 <= 12'he65;
        src102 <= 12'h151;
        src103 <= 12'hbd;
        src104 <= 12'hbfb;
        src105 <= 12'h1f6;
        src106 <= 12'h989;
        src107 <= 12'hb8b;
        src108 <= 12'h3e6;
        src109 <= 12'h7ed;
        src110 <= 12'h4e6;
        src111 <= 12'h581;
        src112 <= 12'hf32;
        src113 <= 12'h682;
        src114 <= 12'hf75;
        src115 <= 12'ha80;
        src116 <= 12'hc1;
        src117 <= 12'h900;
        src118 <= 12'hcea;
        src119 <= 12'hf;
        src120 <= 12'h922;
        src121 <= 12'hee6;
        src122 <= 12'he6c;
        src123 <= 12'hdd9;
        src124 <= 12'h645;
        src125 <= 12'hea5;
        src126 <= 12'he1;
        src127 <= 12'h967;
        src128 <= 12'ha5f;
        src129 <= 12'he5e;
        src130 <= 12'h1eb;
        src131 <= 12'hb7c;
        src132 <= 12'h8a2;
        src133 <= 12'ha99;
        src134 <= 12'h453;
        src135 <= 12'h970;
        src136 <= 12'he72;
        src137 <= 12'hd4d;
        src138 <= 12'hfec;
        src139 <= 12'hac8;
        src140 <= 12'heec;
        src141 <= 12'h62c;
        src142 <= 12'h59c;
        src143 <= 12'h759;
        src144 <= 12'hb6a;
        src145 <= 12'h795;
        src146 <= 12'h44f;
        src147 <= 12'h421;
        src148 <= 12'hf24;
        src149 <= 12'h3ee;
        src150 <= 12'he5a;
        src151 <= 12'he91;
        src152 <= 12'hf11;
        src153 <= 12'ha49;
        src154 <= 12'haf7;
        src155 <= 12'h1e3;
        src156 <= 12'hfd5;
        src157 <= 12'h2ed;
        src158 <= 12'h6d2;
        src159 <= 12'h58e;
        src160 <= 12'hd2f;
        src161 <= 12'h9f8;
        src162 <= 12'h28b;
        src163 <= 12'h629;
        src164 <= 12'hfc0;
        src165 <= 12'hbec;
        src166 <= 12'h9f2;
        src167 <= 12'hf0a;
        src168 <= 12'hfef;
        src169 <= 12'h2f3;
        src170 <= 12'he08;
        src171 <= 12'he5c;
        src172 <= 12'h82c;
        src173 <= 12'h31c;
        src174 <= 12'h152;
        src175 <= 12'h87;
        src176 <= 12'ha03;
        src177 <= 12'hdb5;
        src178 <= 12'hea5;
        src179 <= 12'hde5;
        src180 <= 12'hfbe;
        src181 <= 12'h16d;
        src182 <= 12'h39b;
        src183 <= 12'ha99;
        src184 <= 12'he2c;
        src185 <= 12'hcfb;
        src186 <= 12'hddd;
        src187 <= 12'hec6;
        src188 <= 12'h342;
        exp <= 20'h65cb6;
        #1
        src0 <= 12'hb5f;
        src1 <= 12'h9d5;
        src2 <= 12'h117;
        src3 <= 12'h32e;
        src4 <= 12'he8e;
        src5 <= 12'h43b;
        src6 <= 12'h12f;
        src7 <= 12'hc50;
        src8 <= 12'hab1;
        src9 <= 12'h1f6;
        src10 <= 12'hcc6;
        src11 <= 12'hfd2;
        src12 <= 12'haa3;
        src13 <= 12'h5d7;
        src14 <= 12'h49d;
        src15 <= 12'h6b5;
        src16 <= 12'hf0a;
        src17 <= 12'h144;
        src18 <= 12'h2aa;
        src19 <= 12'h34f;
        src20 <= 12'h81e;
        src21 <= 12'hab;
        src22 <= 12'hc22;
        src23 <= 12'h386;
        src24 <= 12'h3c1;
        src25 <= 12'h947;
        src26 <= 12'hd54;
        src27 <= 12'hdb0;
        src28 <= 12'hf97;
        src29 <= 12'h850;
        src30 <= 12'he64;
        src31 <= 12'h43e;
        src32 <= 12'h870;
        src33 <= 12'h5a6;
        src34 <= 12'h291;
        src35 <= 12'h164;
        src36 <= 12'hc7a;
        src37 <= 12'h5e8;
        src38 <= 12'h2ef;
        src39 <= 12'hf7d;
        src40 <= 12'hfe3;
        src41 <= 12'h323;
        src42 <= 12'hdea;
        src43 <= 12'he51;
        src44 <= 12'h27e;
        src45 <= 12'h2b3;
        src46 <= 12'h890;
        src47 <= 12'hf6c;
        src48 <= 12'h1bf;
        src49 <= 12'hc96;
        src50 <= 12'h45a;
        src51 <= 12'h953;
        src52 <= 12'h81a;
        src53 <= 12'h458;
        src54 <= 12'hb76;
        src55 <= 12'h89e;
        src56 <= 12'h325;
        src57 <= 12'h2a5;
        src58 <= 12'h60c;
        src59 <= 12'hfa2;
        src60 <= 12'he49;
        src61 <= 12'h57d;
        src62 <= 12'h46b;
        src63 <= 12'h3e3;
        src64 <= 12'h131;
        src65 <= 12'h2cc;
        src66 <= 12'h6ef;
        src67 <= 12'h7a3;
        src68 <= 12'h5f;
        src69 <= 12'hcdc;
        src70 <= 12'hf41;
        src71 <= 12'h5a7;
        src72 <= 12'hb7a;
        src73 <= 12'h23a;
        src74 <= 12'h83f;
        src75 <= 12'hffe;
        src76 <= 12'hc2a;
        src77 <= 12'hc2;
        src78 <= 12'hcc6;
        src79 <= 12'h646;
        src80 <= 12'h9d8;
        src81 <= 12'h3a8;
        src82 <= 12'h1c5;
        src83 <= 12'hced;
        src84 <= 12'hbb;
        src85 <= 12'h67a;
        src86 <= 12'hbe7;
        src87 <= 12'h826;
        src88 <= 12'h418;
        src89 <= 12'hb87;
        src90 <= 12'hb65;
        src91 <= 12'hb5f;
        src92 <= 12'hd57;
        src93 <= 12'ha38;
        src94 <= 12'hc93;
        src95 <= 12'h64a;
        src96 <= 12'h64a;
        src97 <= 12'hf66;
        src98 <= 12'he53;
        src99 <= 12'hbd2;
        src100 <= 12'h171;
        src101 <= 12'h5e3;
        src102 <= 12'h82b;
        src103 <= 12'h15a;
        src104 <= 12'h462;
        src105 <= 12'he31;
        src106 <= 12'h452;
        src107 <= 12'hd1a;
        src108 <= 12'he76;
        src109 <= 12'h992;
        src110 <= 12'h4b1;
        src111 <= 12'h8b5;
        src112 <= 12'h47b;
        src113 <= 12'ha44;
        src114 <= 12'hcb5;
        src115 <= 12'hbd5;
        src116 <= 12'h885;
        src117 <= 12'h706;
        src118 <= 12'hd76;
        src119 <= 12'h23e;
        src120 <= 12'h7fa;
        src121 <= 12'h7b6;
        src122 <= 12'ha30;
        src123 <= 12'h198;
        src124 <= 12'hf16;
        src125 <= 12'he60;
        src126 <= 12'h615;
        src127 <= 12'hd30;
        src128 <= 12'h277;
        src129 <= 12'h36c;
        src130 <= 12'h1ac;
        src131 <= 12'hdf1;
        src132 <= 12'h42d;
        src133 <= 12'h821;
        src134 <= 12'hf66;
        src135 <= 12'h14e;
        src136 <= 12'h4d2;
        src137 <= 12'hf17;
        src138 <= 12'hf72;
        src139 <= 12'h150;
        src140 <= 12'hbf3;
        src141 <= 12'h9ea;
        src142 <= 12'h18e;
        src143 <= 12'h5b3;
        src144 <= 12'h31d;
        src145 <= 12'h190;
        src146 <= 12'hda2;
        src147 <= 12'hff1;
        src148 <= 12'h8bf;
        src149 <= 12'h5c3;
        src150 <= 12'h190;
        src151 <= 12'ha65;
        src152 <= 12'h108;
        src153 <= 12'hc7c;
        src154 <= 12'hff0;
        src155 <= 12'h407;
        src156 <= 12'hcc0;
        src157 <= 12'hbf6;
        src158 <= 12'hf22;
        src159 <= 12'hb79;
        src160 <= 12'h329;
        src161 <= 12'h21f;
        src162 <= 12'h5e5;
        src163 <= 12'hae5;
        src164 <= 12'h355;
        src165 <= 12'h436;
        src166 <= 12'h1a;
        src167 <= 12'hc9d;
        src168 <= 12'h330;
        src169 <= 12'h47e;
        src170 <= 12'h3fc;
        src171 <= 12'hbc5;
        src172 <= 12'h59d;
        src173 <= 12'hbb9;
        src174 <= 12'h839;
        src175 <= 12'h4ef;
        src176 <= 12'hced;
        src177 <= 12'h57f;
        src178 <= 12'h4cc;
        src179 <= 12'hd43;
        src180 <= 12'h7f5;
        src181 <= 12'hdfd;
        src182 <= 12'h549;
        src183 <= 12'hb51;
        src184 <= 12'h41a;
        src185 <= 12'h4b2;
        src186 <= 12'hdae;
        src187 <= 12'h95a;
        src188 <= 12'h9bd;
        exp <= 20'h5f1cf;
        #1
        src0 <= 12'hba2;
        src1 <= 12'h5f8;
        src2 <= 12'h7ad;
        src3 <= 12'hf9c;
        src4 <= 12'he2e;
        src5 <= 12'h3db;
        src6 <= 12'h77c;
        src7 <= 12'he0a;
        src8 <= 12'h518;
        src9 <= 12'hc17;
        src10 <= 12'h467;
        src11 <= 12'h67a;
        src12 <= 12'hf14;
        src13 <= 12'hac3;
        src14 <= 12'h4c6;
        src15 <= 12'h48f;
        src16 <= 12'he12;
        src17 <= 12'h137;
        src18 <= 12'h82f;
        src19 <= 12'h8f9;
        src20 <= 12'he86;
        src21 <= 12'h589;
        src22 <= 12'h1fd;
        src23 <= 12'h231;
        src24 <= 12'h983;
        src25 <= 12'hdfa;
        src26 <= 12'h6fb;
        src27 <= 12'h990;
        src28 <= 12'h3e9;
        src29 <= 12'h49c;
        src30 <= 12'h843;
        src31 <= 12'hf39;
        src32 <= 12'h8b;
        src33 <= 12'h55f;
        src34 <= 12'h8c3;
        src35 <= 12'h64f;
        src36 <= 12'hfb5;
        src37 <= 12'hde0;
        src38 <= 12'ha2f;
        src39 <= 12'h2b3;
        src40 <= 12'hec0;
        src41 <= 12'ha21;
        src42 <= 12'hfb5;
        src43 <= 12'h94e;
        src44 <= 12'hbf6;
        src45 <= 12'he9;
        src46 <= 12'h14c;
        src47 <= 12'hcd1;
        src48 <= 12'h691;
        src49 <= 12'had5;
        src50 <= 12'h1f3;
        src51 <= 12'h2d7;
        src52 <= 12'h9dd;
        src53 <= 12'h428;
        src54 <= 12'hda5;
        src55 <= 12'h1cf;
        src56 <= 12'he74;
        src57 <= 12'h9cf;
        src58 <= 12'hdb3;
        src59 <= 12'hf12;
        src60 <= 12'hb80;
        src61 <= 12'h9ae;
        src62 <= 12'hb23;
        src63 <= 12'he54;
        src64 <= 12'h95b;
        src65 <= 12'h193;
        src66 <= 12'h7e2;
        src67 <= 12'h383;
        src68 <= 12'h184;
        src69 <= 12'h70c;
        src70 <= 12'h292;
        src71 <= 12'h1ff;
        src72 <= 12'h1ca;
        src73 <= 12'h7e5;
        src74 <= 12'hb39;
        src75 <= 12'h783;
        src76 <= 12'h690;
        src77 <= 12'h88b;
        src78 <= 12'habd;
        src79 <= 12'he33;
        src80 <= 12'ha82;
        src81 <= 12'hb3;
        src82 <= 12'hfb2;
        src83 <= 12'h734;
        src84 <= 12'hb4d;
        src85 <= 12'h57e;
        src86 <= 12'ha39;
        src87 <= 12'h802;
        src88 <= 12'h704;
        src89 <= 12'h658;
        src90 <= 12'hc15;
        src91 <= 12'h9df;
        src92 <= 12'hc45;
        src93 <= 12'h9b1;
        src94 <= 12'h25f;
        src95 <= 12'ha38;
        src96 <= 12'hcf5;
        src97 <= 12'he5d;
        src98 <= 12'ha0;
        src99 <= 12'h1c;
        src100 <= 12'hf6a;
        src101 <= 12'h8ac;
        src102 <= 12'he63;
        src103 <= 12'h507;
        src104 <= 12'h509;
        src105 <= 12'had5;
        src106 <= 12'hc53;
        src107 <= 12'hf23;
        src108 <= 12'h825;
        src109 <= 12'h3e1;
        src110 <= 12'h64d;
        src111 <= 12'hfed;
        src112 <= 12'h3a;
        src113 <= 12'hb25;
        src114 <= 12'h20c;
        src115 <= 12'he1b;
        src116 <= 12'he30;
        src117 <= 12'h4;
        src118 <= 12'hb86;
        src119 <= 12'haa0;
        src120 <= 12'h657;
        src121 <= 12'h182;
        src122 <= 12'h19c;
        src123 <= 12'hb06;
        src124 <= 12'h89b;
        src125 <= 12'hfd9;
        src126 <= 12'h82d;
        src127 <= 12'h93a;
        src128 <= 12'hd57;
        src129 <= 12'h67a;
        src130 <= 12'h6dc;
        src131 <= 12'he;
        src132 <= 12'h1ac;
        src133 <= 12'heb9;
        src134 <= 12'hf5f;
        src135 <= 12'h803;
        src136 <= 12'h3ec;
        src137 <= 12'h7ba;
        src138 <= 12'h51a;
        src139 <= 12'h9af;
        src140 <= 12'h5b6;
        src141 <= 12'h34;
        src142 <= 12'h22f;
        src143 <= 12'h4a7;
        src144 <= 12'h2d7;
        src145 <= 12'hfec;
        src146 <= 12'hd21;
        src147 <= 12'h135;
        src148 <= 12'h24a;
        src149 <= 12'he0c;
        src150 <= 12'h76;
        src151 <= 12'h4f3;
        src152 <= 12'h9fd;
        src153 <= 12'hd1b;
        src154 <= 12'h8d4;
        src155 <= 12'he19;
        src156 <= 12'hd36;
        src157 <= 12'hd27;
        src158 <= 12'h346;
        src159 <= 12'h5d7;
        src160 <= 12'h200;
        src161 <= 12'ha5d;
        src162 <= 12'h66a;
        src163 <= 12'h24e;
        src164 <= 12'h2e2;
        src165 <= 12'hce3;
        src166 <= 12'h57e;
        src167 <= 12'hbbf;
        src168 <= 12'h521;
        src169 <= 12'h52b;
        src170 <= 12'h390;
        src171 <= 12'hf1;
        src172 <= 12'hbfd;
        src173 <= 12'hc53;
        src174 <= 12'h5c3;
        src175 <= 12'hf41;
        src176 <= 12'h706;
        src177 <= 12'ha42;
        src178 <= 12'h2fd;
        src179 <= 12'he74;
        src180 <= 12'h879;
        src181 <= 12'ha6;
        src182 <= 12'h4fd;
        src183 <= 12'h8b4;
        src184 <= 12'hd6b;
        src185 <= 12'h695;
        src186 <= 12'h2a0;
        src187 <= 12'h24d;
        src188 <= 12'hc7f;
        exp <= 20'h5fd83;
        #1
        src0 <= 12'h5cd;
        src1 <= 12'hddc;
        src2 <= 12'h4bd;
        src3 <= 12'h70d;
        src4 <= 12'h7f9;
        src5 <= 12'h724;
        src6 <= 12'he9c;
        src7 <= 12'hde2;
        src8 <= 12'h1ca;
        src9 <= 12'hf8c;
        src10 <= 12'he67;
        src11 <= 12'h57a;
        src12 <= 12'h963;
        src13 <= 12'ha3d;
        src14 <= 12'hfde;
        src15 <= 12'hfe1;
        src16 <= 12'h212;
        src17 <= 12'h25e;
        src18 <= 12'h9df;
        src19 <= 12'hcaf;
        src20 <= 12'hc81;
        src21 <= 12'h82c;
        src22 <= 12'h48d;
        src23 <= 12'h4b2;
        src24 <= 12'hc5d;
        src25 <= 12'ha2f;
        src26 <= 12'h195;
        src27 <= 12'hdee;
        src28 <= 12'h2cb;
        src29 <= 12'ha9c;
        src30 <= 12'h22f;
        src31 <= 12'h7ef;
        src32 <= 12'ha3b;
        src33 <= 12'h81b;
        src34 <= 12'h5b7;
        src35 <= 12'hca5;
        src36 <= 12'he49;
        src37 <= 12'hc43;
        src38 <= 12'h66a;
        src39 <= 12'h5f0;
        src40 <= 12'hf4c;
        src41 <= 12'hd3a;
        src42 <= 12'h4bc;
        src43 <= 12'h711;
        src44 <= 12'h84a;
        src45 <= 12'h4dd;
        src46 <= 12'h3a1;
        src47 <= 12'hb28;
        src48 <= 12'he3e;
        src49 <= 12'h95d;
        src50 <= 12'h3ca;
        src51 <= 12'h273;
        src52 <= 12'h857;
        src53 <= 12'h8ba;
        src54 <= 12'h161;
        src55 <= 12'hf9c;
        src56 <= 12'h1de;
        src57 <= 12'hff9;
        src58 <= 12'hc32;
        src59 <= 12'hcd0;
        src60 <= 12'h9e1;
        src61 <= 12'h85a;
        src62 <= 12'h3d9;
        src63 <= 12'ha9c;
        src64 <= 12'ha35;
        src65 <= 12'hd0d;
        src66 <= 12'hfd3;
        src67 <= 12'hda5;
        src68 <= 12'h8b9;
        src69 <= 12'h95f;
        src70 <= 12'hd0c;
        src71 <= 12'h7bd;
        src72 <= 12'h802;
        src73 <= 12'hb1e;
        src74 <= 12'hdd4;
        src75 <= 12'h5a5;
        src76 <= 12'hbd;
        src77 <= 12'hf78;
        src78 <= 12'h1c3;
        src79 <= 12'h967;
        src80 <= 12'he46;
        src81 <= 12'h16e;
        src82 <= 12'hea7;
        src83 <= 12'hce3;
        src84 <= 12'he9;
        src85 <= 12'h4a0;
        src86 <= 12'h1ed;
        src87 <= 12'h749;
        src88 <= 12'h70c;
        src89 <= 12'hcca;
        src90 <= 12'h17d;
        src91 <= 12'h8df;
        src92 <= 12'h523;
        src93 <= 12'h7df;
        src94 <= 12'h1d3;
        src95 <= 12'h41;
        src96 <= 12'h235;
        src97 <= 12'h86b;
        src98 <= 12'h16b;
        src99 <= 12'hee8;
        src100 <= 12'h439;
        src101 <= 12'h5e4;
        src102 <= 12'hab;
        src103 <= 12'h84;
        src104 <= 12'hfc;
        src105 <= 12'h965;
        src106 <= 12'hffd;
        src107 <= 12'hda6;
        src108 <= 12'h247;
        src109 <= 12'hfaa;
        src110 <= 12'h8f9;
        src111 <= 12'h5ed;
        src112 <= 12'h799;
        src113 <= 12'h4aa;
        src114 <= 12'h94a;
        src115 <= 12'h871;
        src116 <= 12'h919;
        src117 <= 12'h6e0;
        src118 <= 12'hb1f;
        src119 <= 12'he31;
        src120 <= 12'h618;
        src121 <= 12'h909;
        src122 <= 12'h352;
        src123 <= 12'h3f7;
        src124 <= 12'h957;
        src125 <= 12'h1d1;
        src126 <= 12'h163;
        src127 <= 12'hb52;
        src128 <= 12'h4e4;
        src129 <= 12'had1;
        src130 <= 12'hbc9;
        src131 <= 12'h570;
        src132 <= 12'hb01;
        src133 <= 12'hf0c;
        src134 <= 12'h714;
        src135 <= 12'hf76;
        src136 <= 12'hc46;
        src137 <= 12'h523;
        src138 <= 12'h913;
        src139 <= 12'h59a;
        src140 <= 12'he1;
        src141 <= 12'ha10;
        src142 <= 12'h8d1;
        src143 <= 12'hf0b;
        src144 <= 12'hffc;
        src145 <= 12'hf5b;
        src146 <= 12'h459;
        src147 <= 12'h5bd;
        src148 <= 12'hdb4;
        src149 <= 12'hccd;
        src150 <= 12'hba4;
        src151 <= 12'h33f;
        src152 <= 12'h38f;
        src153 <= 12'ha2f;
        src154 <= 12'hacf;
        src155 <= 12'hf9f;
        src156 <= 12'hf30;
        src157 <= 12'h6f3;
        src158 <= 12'h5b4;
        src159 <= 12'h582;
        src160 <= 12'h22b;
        src161 <= 12'hfb6;
        src162 <= 12'hd23;
        src163 <= 12'h880;
        src164 <= 12'h96d;
        src165 <= 12'h4a7;
        src166 <= 12'h83d;
        src167 <= 12'h672;
        src168 <= 12'hfb2;
        src169 <= 12'h35e;
        src170 <= 12'h32d;
        src171 <= 12'h271;
        src172 <= 12'ha6f;
        src173 <= 12'hf23;
        src174 <= 12'ha37;
        src175 <= 12'hfa9;
        src176 <= 12'h690;
        src177 <= 12'h4b4;
        src178 <= 12'h3c9;
        src179 <= 12'hd9f;
        src180 <= 12'hfa5;
        src181 <= 12'hdd3;
        src182 <= 12'hcd9;
        src183 <= 12'h88b;
        src184 <= 12'he46;
        src185 <= 12'h211;
        src186 <= 12'heb5;
        src187 <= 12'h99c;
        src188 <= 12'h7c4;
        exp <= 20'h66005;
        #1
        src0 <= 12'h1f6;
        src1 <= 12'h664;
        src2 <= 12'hba0;
        src3 <= 12'he50;
        src4 <= 12'ha47;
        src5 <= 12'hed0;
        src6 <= 12'h8f0;
        src7 <= 12'h6ce;
        src8 <= 12'h30d;
        src9 <= 12'hcde;
        src10 <= 12'h117;
        src11 <= 12'h4fb;
        src12 <= 12'hb00;
        src13 <= 12'h9a2;
        src14 <= 12'h9aa;
        src15 <= 12'hebb;
        src16 <= 12'hc15;
        src17 <= 12'h5d0;
        src18 <= 12'hf0b;
        src19 <= 12'hbf9;
        src20 <= 12'h65b;
        src21 <= 12'h205;
        src22 <= 12'hbb3;
        src23 <= 12'hfb;
        src24 <= 12'h11a;
        src25 <= 12'h6b1;
        src26 <= 12'h73a;
        src27 <= 12'hf5d;
        src28 <= 12'hed1;
        src29 <= 12'h385;
        src30 <= 12'h4fd;
        src31 <= 12'h70f;
        src32 <= 12'h92b;
        src33 <= 12'h5a6;
        src34 <= 12'h50a;
        src35 <= 12'h9d5;
        src36 <= 12'h649;
        src37 <= 12'h263;
        src38 <= 12'h169;
        src39 <= 12'h510;
        src40 <= 12'h67d;
        src41 <= 12'h8a1;
        src42 <= 12'hfa9;
        src43 <= 12'hbf7;
        src44 <= 12'h8de;
        src45 <= 12'h129;
        src46 <= 12'h53e;
        src47 <= 12'ha4e;
        src48 <= 12'h995;
        src49 <= 12'h7a9;
        src50 <= 12'h69e;
        src51 <= 12'h23e;
        src52 <= 12'hec1;
        src53 <= 12'h2c2;
        src54 <= 12'h318;
        src55 <= 12'h140;
        src56 <= 12'h17a;
        src57 <= 12'h89f;
        src58 <= 12'hf7f;
        src59 <= 12'hd48;
        src60 <= 12'hde9;
        src61 <= 12'hfcf;
        src62 <= 12'hc1b;
        src63 <= 12'h1a4;
        src64 <= 12'h103;
        src65 <= 12'hc53;
        src66 <= 12'hf2d;
        src67 <= 12'hd30;
        src68 <= 12'h45c;
        src69 <= 12'h52e;
        src70 <= 12'h200;
        src71 <= 12'hd2a;
        src72 <= 12'h632;
        src73 <= 12'h9cb;
        src74 <= 12'hddb;
        src75 <= 12'h138;
        src76 <= 12'h1e;
        src77 <= 12'h6d6;
        src78 <= 12'h579;
        src79 <= 12'had9;
        src80 <= 12'h105;
        src81 <= 12'h9c9;
        src82 <= 12'h33;
        src83 <= 12'h70f;
        src84 <= 12'h950;
        src85 <= 12'h5f7;
        src86 <= 12'h648;
        src87 <= 12'h90c;
        src88 <= 12'h935;
        src89 <= 12'haaf;
        src90 <= 12'he20;
        src91 <= 12'hca3;
        src92 <= 12'ha5b;
        src93 <= 12'h65f;
        src94 <= 12'h946;
        src95 <= 12'hade;
        src96 <= 12'hd17;
        src97 <= 12'hb7e;
        src98 <= 12'hc83;
        src99 <= 12'h201;
        src100 <= 12'h784;
        src101 <= 12'h33c;
        src102 <= 12'hc9d;
        src103 <= 12'h8e1;
        src104 <= 12'h2c6;
        src105 <= 12'hc3;
        src106 <= 12'hf0a;
        src107 <= 12'hada;
        src108 <= 12'h33b;
        src109 <= 12'hf77;
        src110 <= 12'he69;
        src111 <= 12'h2d0;
        src112 <= 12'hfe0;
        src113 <= 12'h6c6;
        src114 <= 12'h9e5;
        src115 <= 12'h475;
        src116 <= 12'hffe;
        src117 <= 12'hcb1;
        src118 <= 12'h8cb;
        src119 <= 12'hbea;
        src120 <= 12'hc6d;
        src121 <= 12'habe;
        src122 <= 12'heb4;
        src123 <= 12'h150;
        src124 <= 12'h42f;
        src125 <= 12'hd39;
        src126 <= 12'hdb8;
        src127 <= 12'h89f;
        src128 <= 12'h4d3;
        src129 <= 12'hcd;
        src130 <= 12'h890;
        src131 <= 12'hde4;
        src132 <= 12'hdba;
        src133 <= 12'h831;
        src134 <= 12'he6a;
        src135 <= 12'hf32;
        src136 <= 12'h7ea;
        src137 <= 12'h86e;
        src138 <= 12'h953;
        src139 <= 12'h57c;
        src140 <= 12'h8e9;
        src141 <= 12'h8ba;
        src142 <= 12'he13;
        src143 <= 12'h58f;
        src144 <= 12'hb6c;
        src145 <= 12'hef1;
        src146 <= 12'h5b2;
        src147 <= 12'h432;
        src148 <= 12'h3bf;
        src149 <= 12'h3d9;
        src150 <= 12'h657;
        src151 <= 12'h653;
        src152 <= 12'hd84;
        src153 <= 12'h4;
        src154 <= 12'h32f;
        src155 <= 12'h553;
        src156 <= 12'h3ff;
        src157 <= 12'ha3a;
        src158 <= 12'h5df;
        src159 <= 12'h3f5;
        src160 <= 12'h14a;
        src161 <= 12'hdec;
        src162 <= 12'h8e4;
        src163 <= 12'h901;
        src164 <= 12'h558;
        src165 <= 12'hf0d;
        src166 <= 12'h3bd;
        src167 <= 12'he74;
        src168 <= 12'h989;
        src169 <= 12'hb86;
        src170 <= 12'h77a;
        src171 <= 12'h415;
        src172 <= 12'h879;
        src173 <= 12'hd4a;
        src174 <= 12'h79f;
        src175 <= 12'hf0e;
        src176 <= 12'hc8b;
        src177 <= 12'h236;
        src178 <= 12'hb4e;
        src179 <= 12'h3f2;
        src180 <= 12'hfca;
        src181 <= 12'h89;
        src182 <= 12'hc9c;
        src183 <= 12'h709;
        src184 <= 12'h9fb;
        src185 <= 12'h5dd;
        src186 <= 12'h6f2;
        src187 <= 12'hbde;
        src188 <= 12'ha9;
        exp <= 20'h61fe8;
        #1
        src0 <= 12'h3ce;
        src1 <= 12'hd5c;
        src2 <= 12'h88b;
        src3 <= 12'hbb1;
        src4 <= 12'h24c;
        src5 <= 12'had2;
        src6 <= 12'h100;
        src7 <= 12'h2e8;
        src8 <= 12'hab4;
        src9 <= 12'hffd;
        src10 <= 12'h435;
        src11 <= 12'ha19;
        src12 <= 12'h1fb;
        src13 <= 12'ha82;
        src14 <= 12'hf4b;
        src15 <= 12'hd44;
        src16 <= 12'hae6;
        src17 <= 12'hbfd;
        src18 <= 12'h2e5;
        src19 <= 12'h35e;
        src20 <= 12'hf35;
        src21 <= 12'hc84;
        src22 <= 12'h9b4;
        src23 <= 12'h8d2;
        src24 <= 12'hbfd;
        src25 <= 12'h4c;
        src26 <= 12'h4b0;
        src27 <= 12'h6b6;
        src28 <= 12'h290;
        src29 <= 12'hb4;
        src30 <= 12'h39c;
        src31 <= 12'h693;
        src32 <= 12'he84;
        src33 <= 12'hcb8;
        src34 <= 12'hc2e;
        src35 <= 12'ha15;
        src36 <= 12'hf12;
        src37 <= 12'h949;
        src38 <= 12'he82;
        src39 <= 12'hb60;
        src40 <= 12'h3fc;
        src41 <= 12'h31;
        src42 <= 12'h20a;
        src43 <= 12'h751;
        src44 <= 12'hc60;
        src45 <= 12'h891;
        src46 <= 12'h18c;
        src47 <= 12'h2e9;
        src48 <= 12'hbb8;
        src49 <= 12'hcb;
        src50 <= 12'h662;
        src51 <= 12'h5cc;
        src52 <= 12'h579;
        src53 <= 12'h75e;
        src54 <= 12'hbea;
        src55 <= 12'h97;
        src56 <= 12'h471;
        src57 <= 12'ha2e;
        src58 <= 12'h870;
        src59 <= 12'hb84;
        src60 <= 12'h88a;
        src61 <= 12'h94;
        src62 <= 12'h89f;
        src63 <= 12'h92f;
        src64 <= 12'hfb2;
        src65 <= 12'h5e4;
        src66 <= 12'h8f5;
        src67 <= 12'h8b4;
        src68 <= 12'he4a;
        src69 <= 12'h863;
        src70 <= 12'h7e8;
        src71 <= 12'h912;
        src72 <= 12'h172;
        src73 <= 12'h8b0;
        src74 <= 12'h1b4;
        src75 <= 12'hdb4;
        src76 <= 12'h9fd;
        src77 <= 12'he75;
        src78 <= 12'h521;
        src79 <= 12'h6ac;
        src80 <= 12'h5bf;
        src81 <= 12'h5ef;
        src82 <= 12'h165;
        src83 <= 12'h15e;
        src84 <= 12'hcb6;
        src85 <= 12'h301;
        src86 <= 12'hc10;
        src87 <= 12'hac7;
        src88 <= 12'h580;
        src89 <= 12'h1b0;
        src90 <= 12'hf13;
        src91 <= 12'h59d;
        src92 <= 12'hfe7;
        src93 <= 12'h43a;
        src94 <= 12'h278;
        src95 <= 12'h6c0;
        src96 <= 12'h9ec;
        src97 <= 12'h6c6;
        src98 <= 12'hd2f;
        src99 <= 12'hc9a;
        src100 <= 12'hefd;
        src101 <= 12'hc8c;
        src102 <= 12'hc1e;
        src103 <= 12'h457;
        src104 <= 12'ha17;
        src105 <= 12'h5c4;
        src106 <= 12'h7c6;
        src107 <= 12'h1d4;
        src108 <= 12'h86a;
        src109 <= 12'h2b2;
        src110 <= 12'hdb9;
        src111 <= 12'hc2f;
        src112 <= 12'ha07;
        src113 <= 12'hba4;
        src114 <= 12'h6cc;
        src115 <= 12'h716;
        src116 <= 12'h4e7;
        src117 <= 12'hc9a;
        src118 <= 12'h136;
        src119 <= 12'hbb8;
        src120 <= 12'h46b;
        src121 <= 12'he9f;
        src122 <= 12'hf55;
        src123 <= 12'he38;
        src124 <= 12'h148;
        src125 <= 12'hac6;
        src126 <= 12'hb4b;
        src127 <= 12'h3c7;
        src128 <= 12'h827;
        src129 <= 12'h5f8;
        src130 <= 12'h563;
        src131 <= 12'hd46;
        src132 <= 12'hf3b;
        src133 <= 12'hbf2;
        src134 <= 12'h474;
        src135 <= 12'h722;
        src136 <= 12'he40;
        src137 <= 12'h9ab;
        src138 <= 12'hf30;
        src139 <= 12'h867;
        src140 <= 12'h568;
        src141 <= 12'hbae;
        src142 <= 12'haf4;
        src143 <= 12'hf2a;
        src144 <= 12'h664;
        src145 <= 12'hea0;
        src146 <= 12'hd9f;
        src147 <= 12'hfca;
        src148 <= 12'h904;
        src149 <= 12'hc6;
        src150 <= 12'h29f;
        src151 <= 12'hf46;
        src152 <= 12'hfe0;
        src153 <= 12'h197;
        src154 <= 12'h306;
        src155 <= 12'h9a8;
        src156 <= 12'he1;
        src157 <= 12'h461;
        src158 <= 12'he46;
        src159 <= 12'h64d;
        src160 <= 12'h230;
        src161 <= 12'h16e;
        src162 <= 12'h77f;
        src163 <= 12'h408;
        src164 <= 12'h3a6;
        src165 <= 12'hae7;
        src166 <= 12'h436;
        src167 <= 12'he4;
        src168 <= 12'h528;
        src169 <= 12'h2c3;
        src170 <= 12'h2de;
        src171 <= 12'h8c2;
        src172 <= 12'h4c9;
        src173 <= 12'h291;
        src174 <= 12'hcc4;
        src175 <= 12'h81b;
        src176 <= 12'hcff;
        src177 <= 12'hb0c;
        src178 <= 12'h26b;
        src179 <= 12'hc2b;
        src180 <= 12'h45a;
        src181 <= 12'h632;
        src182 <= 12'hc52;
        src183 <= 12'hbf;
        src184 <= 12'hf1b;
        src185 <= 12'hfd8;
        src186 <= 12'h8b0;
        src187 <= 12'h4bb;
        src188 <= 12'h682;
        exp <= 20'h5fcc1;
        #1
        src0 <= 12'h572;
        src1 <= 12'hbc2;
        src2 <= 12'h971;
        src3 <= 12'hdb1;
        src4 <= 12'h860;
        src5 <= 12'he67;
        src6 <= 12'h119;
        src7 <= 12'ha59;
        src8 <= 12'hd78;
        src9 <= 12'h683;
        src10 <= 12'he9b;
        src11 <= 12'h5fb;
        src12 <= 12'h342;
        src13 <= 12'hd53;
        src14 <= 12'h156;
        src15 <= 12'h7c6;
        src16 <= 12'h7a1;
        src17 <= 12'h4b3;
        src18 <= 12'hb6a;
        src19 <= 12'hd88;
        src20 <= 12'hafc;
        src21 <= 12'hafa;
        src22 <= 12'hd99;
        src23 <= 12'h81a;
        src24 <= 12'h3c6;
        src25 <= 12'ha68;
        src26 <= 12'h7f5;
        src27 <= 12'h750;
        src28 <= 12'h675;
        src29 <= 12'h497;
        src30 <= 12'hceb;
        src31 <= 12'hf2c;
        src32 <= 12'h8fb;
        src33 <= 12'h57c;
        src34 <= 12'hcab;
        src35 <= 12'h754;
        src36 <= 12'hba0;
        src37 <= 12'h1fa;
        src38 <= 12'h1b3;
        src39 <= 12'hd84;
        src40 <= 12'h6b2;
        src41 <= 12'h732;
        src42 <= 12'hf87;
        src43 <= 12'h7fc;
        src44 <= 12'h14;
        src45 <= 12'hff3;
        src46 <= 12'h23f;
        src47 <= 12'he5c;
        src48 <= 12'h55b;
        src49 <= 12'hd41;
        src50 <= 12'h367;
        src51 <= 12'hdcc;
        src52 <= 12'h4c3;
        src53 <= 12'ha90;
        src54 <= 12'h960;
        src55 <= 12'h237;
        src56 <= 12'h34;
        src57 <= 12'hf6;
        src58 <= 12'h834;
        src59 <= 12'h194;
        src60 <= 12'hdf5;
        src61 <= 12'hc6e;
        src62 <= 12'hfb5;
        src63 <= 12'h1f;
        src64 <= 12'h9a;
        src65 <= 12'h1bd;
        src66 <= 12'hd7e;
        src67 <= 12'h2d5;
        src68 <= 12'hf69;
        src69 <= 12'h395;
        src70 <= 12'h2dc;
        src71 <= 12'ha95;
        src72 <= 12'h578;
        src73 <= 12'hb69;
        src74 <= 12'h52d;
        src75 <= 12'h875;
        src76 <= 12'h476;
        src77 <= 12'h103;
        src78 <= 12'hba;
        src79 <= 12'h7e4;
        src80 <= 12'hb0f;
        src81 <= 12'h27b;
        src82 <= 12'ha6c;
        src83 <= 12'hbd5;
        src84 <= 12'ha14;
        src85 <= 12'h58d;
        src86 <= 12'h16c;
        src87 <= 12'h2bc;
        src88 <= 12'hd43;
        src89 <= 12'h5af;
        src90 <= 12'heb0;
        src91 <= 12'hb6b;
        src92 <= 12'ha68;
        src93 <= 12'h6d6;
        src94 <= 12'h6ee;
        src95 <= 12'hf1e;
        src96 <= 12'h1f9;
        src97 <= 12'h62;
        src98 <= 12'h37d;
        src99 <= 12'h4;
        src100 <= 12'hde5;
        src101 <= 12'h678;
        src102 <= 12'h867;
        src103 <= 12'hc52;
        src104 <= 12'hbee;
        src105 <= 12'h7c4;
        src106 <= 12'h753;
        src107 <= 12'h114;
        src108 <= 12'h5fb;
        src109 <= 12'h974;
        src110 <= 12'hc0b;
        src111 <= 12'h75e;
        src112 <= 12'hc06;
        src113 <= 12'hc4b;
        src114 <= 12'hb8e;
        src115 <= 12'h8a2;
        src116 <= 12'h334;
        src117 <= 12'h914;
        src118 <= 12'h7e2;
        src119 <= 12'hfb6;
        src120 <= 12'he46;
        src121 <= 12'heb3;
        src122 <= 12'h1a6;
        src123 <= 12'hf42;
        src124 <= 12'h152;
        src125 <= 12'h329;
        src126 <= 12'hbe6;
        src127 <= 12'hb9f;
        src128 <= 12'h499;
        src129 <= 12'ha4;
        src130 <= 12'he2d;
        src131 <= 12'h6c8;
        src132 <= 12'h95c;
        src133 <= 12'h274;
        src134 <= 12'hc27;
        src135 <= 12'h28d;
        src136 <= 12'h89f;
        src137 <= 12'hbf;
        src138 <= 12'h42b;
        src139 <= 12'h8e1;
        src140 <= 12'h5b9;
        src141 <= 12'h954;
        src142 <= 12'hf39;
        src143 <= 12'h866;
        src144 <= 12'h550;
        src145 <= 12'h21c;
        src146 <= 12'hb1;
        src147 <= 12'h1a2;
        src148 <= 12'h621;
        src149 <= 12'h712;
        src150 <= 12'h7cc;
        src151 <= 12'h914;
        src152 <= 12'h7f0;
        src153 <= 12'h10e;
        src154 <= 12'haa7;
        src155 <= 12'hd3;
        src156 <= 12'h817;
        src157 <= 12'ha9c;
        src158 <= 12'h7f;
        src159 <= 12'h5cf;
        src160 <= 12'he11;
        src161 <= 12'hd39;
        src162 <= 12'hee;
        src163 <= 12'h1f7;
        src164 <= 12'h96d;
        src165 <= 12'h1fe;
        src166 <= 12'h5f0;
        src167 <= 12'ha22;
        src168 <= 12'heab;
        src169 <= 12'h1cd;
        src170 <= 12'hfa1;
        src171 <= 12'he20;
        src172 <= 12'h702;
        src173 <= 12'h6f0;
        src174 <= 12'hd5e;
        src175 <= 12'h4ab;
        src176 <= 12'h4c9;
        src177 <= 12'hdd5;
        src178 <= 12'h335;
        src179 <= 12'heea;
        src180 <= 12'h6e3;
        src181 <= 12'h5;
        src182 <= 12'h604;
        src183 <= 12'he64;
        src184 <= 12'h78d;
        src185 <= 12'h9;
        src186 <= 12'h581;
        src187 <= 12'h512;
        src188 <= 12'h846;
        exp <= 20'h5b8be;
        #1
        src0 <= 12'haed;
        src1 <= 12'hc39;
        src2 <= 12'h9cc;
        src3 <= 12'hc14;
        src4 <= 12'h469;
        src5 <= 12'had1;
        src6 <= 12'he1;
        src7 <= 12'h505;
        src8 <= 12'h3a8;
        src9 <= 12'hbf8;
        src10 <= 12'h3de;
        src11 <= 12'hfb3;
        src12 <= 12'h8a5;
        src13 <= 12'h4da;
        src14 <= 12'h85d;
        src15 <= 12'hea7;
        src16 <= 12'hfa2;
        src17 <= 12'heac;
        src18 <= 12'he47;
        src19 <= 12'hdf3;
        src20 <= 12'ha17;
        src21 <= 12'h8e;
        src22 <= 12'he25;
        src23 <= 12'h701;
        src24 <= 12'h75b;
        src25 <= 12'hbb3;
        src26 <= 12'h4cc;
        src27 <= 12'h9f1;
        src28 <= 12'h51a;
        src29 <= 12'hfb6;
        src30 <= 12'h295;
        src31 <= 12'h70b;
        src32 <= 12'hdcc;
        src33 <= 12'h9be;
        src34 <= 12'h2c6;
        src35 <= 12'ha4e;
        src36 <= 12'h80;
        src37 <= 12'h8cc;
        src38 <= 12'hd5b;
        src39 <= 12'hbfc;
        src40 <= 12'hd5f;
        src41 <= 12'hc60;
        src42 <= 12'h11;
        src43 <= 12'h49a;
        src44 <= 12'ha62;
        src45 <= 12'h795;
        src46 <= 12'h130;
        src47 <= 12'h497;
        src48 <= 12'hcd1;
        src49 <= 12'h107;
        src50 <= 12'h833;
        src51 <= 12'hd52;
        src52 <= 12'h2da;
        src53 <= 12'h1d4;
        src54 <= 12'hbf3;
        src55 <= 12'h676;
        src56 <= 12'h998;
        src57 <= 12'haf0;
        src58 <= 12'hcd;
        src59 <= 12'h812;
        src60 <= 12'h261;
        src61 <= 12'hd36;
        src62 <= 12'h259;
        src63 <= 12'h906;
        src64 <= 12'hca2;
        src65 <= 12'h688;
        src66 <= 12'h95c;
        src67 <= 12'h1e;
        src68 <= 12'h8c2;
        src69 <= 12'hf47;
        src70 <= 12'h19f;
        src71 <= 12'hb96;
        src72 <= 12'h4dc;
        src73 <= 12'hf8b;
        src74 <= 12'ha74;
        src75 <= 12'hb72;
        src76 <= 12'h49;
        src77 <= 12'h5ff;
        src78 <= 12'h83e;
        src79 <= 12'h160;
        src80 <= 12'h933;
        src81 <= 12'h25c;
        src82 <= 12'hcf3;
        src83 <= 12'h4d4;
        src84 <= 12'h5cc;
        src85 <= 12'h64f;
        src86 <= 12'h436;
        src87 <= 12'hf0c;
        src88 <= 12'h82;
        src89 <= 12'h97a;
        src90 <= 12'hbc5;
        src91 <= 12'hb0c;
        src92 <= 12'hc9d;
        src93 <= 12'h590;
        src94 <= 12'h24d;
        src95 <= 12'h5eb;
        src96 <= 12'h4ad;
        src97 <= 12'h8e8;
        src98 <= 12'hf5e;
        src99 <= 12'h345;
        src100 <= 12'h5e;
        src101 <= 12'h7a1;
        src102 <= 12'ha63;
        src103 <= 12'hae9;
        src104 <= 12'h3cb;
        src105 <= 12'haf5;
        src106 <= 12'h175;
        src107 <= 12'h7ab;
        src108 <= 12'h48b;
        src109 <= 12'hdbd;
        src110 <= 12'h67d;
        src111 <= 12'he2f;
        src112 <= 12'h5f;
        src113 <= 12'h680;
        src114 <= 12'h98b;
        src115 <= 12'h8a6;
        src116 <= 12'hd84;
        src117 <= 12'hf10;
        src118 <= 12'hfa9;
        src119 <= 12'h381;
        src120 <= 12'hcc3;
        src121 <= 12'hd2e;
        src122 <= 12'h8b;
        src123 <= 12'h672;
        src124 <= 12'h66e;
        src125 <= 12'he0c;
        src126 <= 12'hcdd;
        src127 <= 12'h846;
        src128 <= 12'hae2;
        src129 <= 12'h702;
        src130 <= 12'h593;
        src131 <= 12'hb5e;
        src132 <= 12'hc44;
        src133 <= 12'hc81;
        src134 <= 12'hee5;
        src135 <= 12'hd79;
        src136 <= 12'h621;
        src137 <= 12'h1db;
        src138 <= 12'h1e9;
        src139 <= 12'h227;
        src140 <= 12'h5f4;
        src141 <= 12'h754;
        src142 <= 12'ha82;
        src143 <= 12'hde2;
        src144 <= 12'hd72;
        src145 <= 12'h1da;
        src146 <= 12'hb3d;
        src147 <= 12'hd1d;
        src148 <= 12'hcc7;
        src149 <= 12'h34a;
        src150 <= 12'hcb5;
        src151 <= 12'hf4b;
        src152 <= 12'h1a3;
        src153 <= 12'hc9f;
        src154 <= 12'h73c;
        src155 <= 12'h903;
        src156 <= 12'hb7e;
        src157 <= 12'h3c4;
        src158 <= 12'h21e;
        src159 <= 12'hc99;
        src160 <= 12'he8e;
        src161 <= 12'hd52;
        src162 <= 12'h3d5;
        src163 <= 12'hff2;
        src164 <= 12'h2c5;
        src165 <= 12'h606;
        src166 <= 12'hb30;
        src167 <= 12'hf86;
        src168 <= 12'hb7b;
        src169 <= 12'h39c;
        src170 <= 12'h903;
        src171 <= 12'h517;
        src172 <= 12'h501;
        src173 <= 12'h9c7;
        src174 <= 12'h522;
        src175 <= 12'ha2c;
        src176 <= 12'h213;
        src177 <= 12'hb4;
        src178 <= 12'hc4e;
        src179 <= 12'h9dc;
        src180 <= 12'h4bc;
        src181 <= 12'h609;
        src182 <= 12'hde4;
        src183 <= 12'hf5b;
        src184 <= 12'h874;
        src185 <= 12'hb99;
        src186 <= 12'ha84;
        src187 <= 12'hddd;
        src188 <= 12'h74e;
        exp <= 20'h6354d;
        #1
        src0 <= 12'hfe6;
        src1 <= 12'h445;
        src2 <= 12'h620;
        src3 <= 12'h44b;
        src4 <= 12'hdd1;
        src5 <= 12'h937;
        src6 <= 12'h7c7;
        src7 <= 12'h93d;
        src8 <= 12'h216;
        src9 <= 12'h7a9;
        src10 <= 12'h55a;
        src11 <= 12'h1d4;
        src12 <= 12'haac;
        src13 <= 12'hee2;
        src14 <= 12'h11a;
        src15 <= 12'h6bb;
        src16 <= 12'h627;
        src17 <= 12'h1d4;
        src18 <= 12'h246;
        src19 <= 12'h4d1;
        src20 <= 12'hca0;
        src21 <= 12'h11c;
        src22 <= 12'h809;
        src23 <= 12'h4b;
        src24 <= 12'hf35;
        src25 <= 12'h626;
        src26 <= 12'hbae;
        src27 <= 12'h8c9;
        src28 <= 12'h75;
        src29 <= 12'hb9c;
        src30 <= 12'h138;
        src31 <= 12'hba6;
        src32 <= 12'he84;
        src33 <= 12'h3;
        src34 <= 12'hab5;
        src35 <= 12'hc42;
        src36 <= 12'h989;
        src37 <= 12'h920;
        src38 <= 12'h198;
        src39 <= 12'h38;
        src40 <= 12'h1cb;
        src41 <= 12'he2f;
        src42 <= 12'hf0d;
        src43 <= 12'hf29;
        src44 <= 12'hf01;
        src45 <= 12'hd80;
        src46 <= 12'h6e;
        src47 <= 12'h827;
        src48 <= 12'h57f;
        src49 <= 12'he79;
        src50 <= 12'h519;
        src51 <= 12'hfbc;
        src52 <= 12'h43a;
        src53 <= 12'h9c9;
        src54 <= 12'hf54;
        src55 <= 12'hcdc;
        src56 <= 12'h8c5;
        src57 <= 12'h5c5;
        src58 <= 12'h170;
        src59 <= 12'h4af;
        src60 <= 12'h20f;
        src61 <= 12'h6c7;
        src62 <= 12'hd99;
        src63 <= 12'h3f5;
        src64 <= 12'h9bb;
        src65 <= 12'h1b8;
        src66 <= 12'h558;
        src67 <= 12'h440;
        src68 <= 12'h344;
        src69 <= 12'hbf2;
        src70 <= 12'h51b;
        src71 <= 12'hcc5;
        src72 <= 12'hf23;
        src73 <= 12'hd2e;
        src74 <= 12'h72e;
        src75 <= 12'hf57;
        src76 <= 12'hf93;
        src77 <= 12'h924;
        src78 <= 12'h433;
        src79 <= 12'hf51;
        src80 <= 12'h38b;
        src81 <= 12'hc1c;
        src82 <= 12'hd2;
        src83 <= 12'h7d7;
        src84 <= 12'h5df;
        src85 <= 12'ha0f;
        src86 <= 12'hc97;
        src87 <= 12'h421;
        src88 <= 12'hb92;
        src89 <= 12'h9a2;
        src90 <= 12'h30;
        src91 <= 12'hc0;
        src92 <= 12'h831;
        src93 <= 12'hc46;
        src94 <= 12'hf73;
        src95 <= 12'h6a6;
        src96 <= 12'hfa0;
        src97 <= 12'h75c;
        src98 <= 12'h142;
        src99 <= 12'h8ea;
        src100 <= 12'h9fb;
        src101 <= 12'he3a;
        src102 <= 12'h3b9;
        src103 <= 12'h27a;
        src104 <= 12'h3fc;
        src105 <= 12'h604;
        src106 <= 12'h892;
        src107 <= 12'he8f;
        src108 <= 12'h58d;
        src109 <= 12'h2aa;
        src110 <= 12'h709;
        src111 <= 12'h706;
        src112 <= 12'hf65;
        src113 <= 12'ha9a;
        src114 <= 12'hc73;
        src115 <= 12'h8f4;
        src116 <= 12'hab5;
        src117 <= 12'h6b6;
        src118 <= 12'hc5f;
        src119 <= 12'h6ad;
        src120 <= 12'h7c2;
        src121 <= 12'h188;
        src122 <= 12'hadb;
        src123 <= 12'h650;
        src124 <= 12'h3e8;
        src125 <= 12'h667;
        src126 <= 12'hf66;
        src127 <= 12'hc0b;
        src128 <= 12'h443;
        src129 <= 12'hdb1;
        src130 <= 12'h7e8;
        src131 <= 12'ha6b;
        src132 <= 12'h15;
        src133 <= 12'haf1;
        src134 <= 12'ha74;
        src135 <= 12'he2a;
        src136 <= 12'hd93;
        src137 <= 12'h177;
        src138 <= 12'h29e;
        src139 <= 12'hddf;
        src140 <= 12'hb73;
        src141 <= 12'h5c6;
        src142 <= 12'h742;
        src143 <= 12'ha5b;
        src144 <= 12'hd3e;
        src145 <= 12'hac;
        src146 <= 12'ha6e;
        src147 <= 12'hc5;
        src148 <= 12'h180;
        src149 <= 12'h4a9;
        src150 <= 12'ha70;
        src151 <= 12'hbf8;
        src152 <= 12'h25c;
        src153 <= 12'h8c2;
        src154 <= 12'h39c;
        src155 <= 12'hff7;
        src156 <= 12'ha2a;
        src157 <= 12'hf35;
        src158 <= 12'hb4e;
        src159 <= 12'he19;
        src160 <= 12'hb1d;
        src161 <= 12'h6c4;
        src162 <= 12'hb39;
        src163 <= 12'hcb3;
        src164 <= 12'hb69;
        src165 <= 12'hd76;
        src166 <= 12'h2b7;
        src167 <= 12'hb3e;
        src168 <= 12'hd6c;
        src169 <= 12'h782;
        src170 <= 12'h1fd;
        src171 <= 12'h3b3;
        src172 <= 12'h820;
        src173 <= 12'ha0e;
        src174 <= 12'h367;
        src175 <= 12'h433;
        src176 <= 12'h40;
        src177 <= 12'h86d;
        src178 <= 12'h9fb;
        src179 <= 12'h522;
        src180 <= 12'hea6;
        src181 <= 12'h9d;
        src182 <= 12'h26;
        src183 <= 12'h642;
        src184 <= 12'hd8f;
        src185 <= 12'h176;
        src186 <= 12'h1da;
        src187 <= 12'h808;
        src188 <= 12'hfd6;
        exp <= 20'h5f6aa;
        #1
        src0 <= 12'h850;
        src1 <= 12'h78;
        src2 <= 12'h391;
        src3 <= 12'h9a9;
        src4 <= 12'h3df;
        src5 <= 12'h377;
        src6 <= 12'h33e;
        src7 <= 12'h6f9;
        src8 <= 12'h6bf;
        src9 <= 12'hfcc;
        src10 <= 12'h677;
        src11 <= 12'h2e;
        src12 <= 12'h77a;
        src13 <= 12'hdf6;
        src14 <= 12'hb62;
        src15 <= 12'he50;
        src16 <= 12'h94b;
        src17 <= 12'h3a3;
        src18 <= 12'h8ef;
        src19 <= 12'h1f;
        src20 <= 12'h988;
        src21 <= 12'h948;
        src22 <= 12'hf4;
        src23 <= 12'h444;
        src24 <= 12'h657;
        src25 <= 12'hb1d;
        src26 <= 12'hab8;
        src27 <= 12'hd29;
        src28 <= 12'h9b0;
        src29 <= 12'hf68;
        src30 <= 12'h15d;
        src31 <= 12'hfdf;
        src32 <= 12'h2bf;
        src33 <= 12'h22;
        src34 <= 12'h4ec;
        src35 <= 12'h79d;
        src36 <= 12'hc73;
        src37 <= 12'h4e;
        src38 <= 12'h6a0;
        src39 <= 12'h633;
        src40 <= 12'h53;
        src41 <= 12'h247;
        src42 <= 12'h335;
        src43 <= 12'hc41;
        src44 <= 12'hd1d;
        src45 <= 12'h82a;
        src46 <= 12'h686;
        src47 <= 12'h55a;
        src48 <= 12'h240;
        src49 <= 12'hba4;
        src50 <= 12'hb49;
        src51 <= 12'he2f;
        src52 <= 12'he5d;
        src53 <= 12'h214;
        src54 <= 12'h18c;
        src55 <= 12'h2b8;
        src56 <= 12'h4a2;
        src57 <= 12'h1;
        src58 <= 12'h1c2;
        src59 <= 12'h44b;
        src60 <= 12'he6a;
        src61 <= 12'h501;
        src62 <= 12'h3ce;
        src63 <= 12'h785;
        src64 <= 12'h59b;
        src65 <= 12'ha3c;
        src66 <= 12'h9c;
        src67 <= 12'had8;
        src68 <= 12'h3cc;
        src69 <= 12'h681;
        src70 <= 12'h838;
        src71 <= 12'h65e;
        src72 <= 12'hd7f;
        src73 <= 12'h5d6;
        src74 <= 12'h447;
        src75 <= 12'h7e0;
        src76 <= 12'h384;
        src77 <= 12'h331;
        src78 <= 12'h1fc;
        src79 <= 12'h6d5;
        src80 <= 12'hc3;
        src81 <= 12'h5c0;
        src82 <= 12'h9b5;
        src83 <= 12'h107;
        src84 <= 12'hb57;
        src85 <= 12'h4f3;
        src86 <= 12'hba9;
        src87 <= 12'h9dd;
        src88 <= 12'h942;
        src89 <= 12'h758;
        src90 <= 12'h47c;
        src91 <= 12'h35f;
        src92 <= 12'hfc;
        src93 <= 12'h6d4;
        src94 <= 12'hdd8;
        src95 <= 12'hd36;
        src96 <= 12'h8ca;
        src97 <= 12'h5;
        src98 <= 12'h340;
        src99 <= 12'hd04;
        src100 <= 12'hcff;
        src101 <= 12'h720;
        src102 <= 12'h39a;
        src103 <= 12'h60c;
        src104 <= 12'h954;
        src105 <= 12'h1c4;
        src106 <= 12'h5c3;
        src107 <= 12'h8ca;
        src108 <= 12'ha2a;
        src109 <= 12'h3ef;
        src110 <= 12'h1e0;
        src111 <= 12'hd3c;
        src112 <= 12'h296;
        src113 <= 12'hb63;
        src114 <= 12'hc85;
        src115 <= 12'hbbd;
        src116 <= 12'h83c;
        src117 <= 12'h4f6;
        src118 <= 12'he7f;
        src119 <= 12'h4c8;
        src120 <= 12'h8c1;
        src121 <= 12'hb51;
        src122 <= 12'hf96;
        src123 <= 12'h76a;
        src124 <= 12'h970;
        src125 <= 12'hd18;
        src126 <= 12'hddc;
        src127 <= 12'h548;
        src128 <= 12'hb46;
        src129 <= 12'hf0e;
        src130 <= 12'h284;
        src131 <= 12'h25f;
        src132 <= 12'he17;
        src133 <= 12'he15;
        src134 <= 12'h32;
        src135 <= 12'h753;
        src136 <= 12'h8fc;
        src137 <= 12'h448;
        src138 <= 12'h144;
        src139 <= 12'hf36;
        src140 <= 12'h654;
        src141 <= 12'h187;
        src142 <= 12'h288;
        src143 <= 12'h313;
        src144 <= 12'h58d;
        src145 <= 12'hd9b;
        src146 <= 12'h2b;
        src147 <= 12'hf86;
        src148 <= 12'hd20;
        src149 <= 12'hd48;
        src150 <= 12'h8c7;
        src151 <= 12'h718;
        src152 <= 12'h24f;
        src153 <= 12'h926;
        src154 <= 12'h250;
        src155 <= 12'h45e;
        src156 <= 12'haac;
        src157 <= 12'h61;
        src158 <= 12'h8a3;
        src159 <= 12'h5aa;
        src160 <= 12'he91;
        src161 <= 12'h8c0;
        src162 <= 12'h83a;
        src163 <= 12'hc3b;
        src164 <= 12'h96e;
        src165 <= 12'he5f;
        src166 <= 12'ha93;
        src167 <= 12'h6b9;
        src168 <= 12'hab6;
        src169 <= 12'h268;
        src170 <= 12'he5e;
        src171 <= 12'h2d2;
        src172 <= 12'hf40;
        src173 <= 12'hf95;
        src174 <= 12'haf0;
        src175 <= 12'he1;
        src176 <= 12'hcf7;
        src177 <= 12'h2e9;
        src178 <= 12'h861;
        src179 <= 12'hfd5;
        src180 <= 12'hbd6;
        src181 <= 12'hd75;
        src182 <= 12'h34e;
        src183 <= 12'h4de;
        src184 <= 12'h64c;
        src185 <= 12'h512;
        src186 <= 12'h738;
        src187 <= 12'hffd;
        src188 <= 12'h193;
        exp <= 20'h58837;
        #1
        src0 <= 12'hf35;
        src1 <= 12'h573;
        src2 <= 12'h418;
        src3 <= 12'hd98;
        src4 <= 12'h42b;
        src5 <= 12'h80c;
        src6 <= 12'ha09;
        src7 <= 12'he2c;
        src8 <= 12'heff;
        src9 <= 12'ha18;
        src10 <= 12'hc4e;
        src11 <= 12'hb01;
        src12 <= 12'hc64;
        src13 <= 12'h22e;
        src14 <= 12'he49;
        src15 <= 12'hd24;
        src16 <= 12'hd2b;
        src17 <= 12'had;
        src18 <= 12'h26b;
        src19 <= 12'ha7;
        src20 <= 12'h716;
        src21 <= 12'h400;
        src22 <= 12'hef;
        src23 <= 12'h10;
        src24 <= 12'he26;
        src25 <= 12'h692;
        src26 <= 12'h6a8;
        src27 <= 12'hf5c;
        src28 <= 12'h3b8;
        src29 <= 12'ha3d;
        src30 <= 12'hcdc;
        src31 <= 12'h32a;
        src32 <= 12'h23f;
        src33 <= 12'h364;
        src34 <= 12'habd;
        src35 <= 12'hd28;
        src36 <= 12'hfdf;
        src37 <= 12'h484;
        src38 <= 12'hf85;
        src39 <= 12'hef5;
        src40 <= 12'h23a;
        src41 <= 12'h2b7;
        src42 <= 12'h36b;
        src43 <= 12'hb5a;
        src44 <= 12'h27a;
        src45 <= 12'hd95;
        src46 <= 12'hb87;
        src47 <= 12'had9;
        src48 <= 12'h58b;
        src49 <= 12'hfda;
        src50 <= 12'h117;
        src51 <= 12'ha8e;
        src52 <= 12'hdbc;
        src53 <= 12'h5cd;
        src54 <= 12'h950;
        src55 <= 12'h3fc;
        src56 <= 12'h97e;
        src57 <= 12'h190;
        src58 <= 12'h75;
        src59 <= 12'h558;
        src60 <= 12'h41e;
        src61 <= 12'h1a3;
        src62 <= 12'h3cf;
        src63 <= 12'hb34;
        src64 <= 12'h451;
        src65 <= 12'h53;
        src66 <= 12'hc55;
        src67 <= 12'h76f;
        src68 <= 12'h894;
        src69 <= 12'ha56;
        src70 <= 12'hd01;
        src71 <= 12'hb9a;
        src72 <= 12'he24;
        src73 <= 12'he18;
        src74 <= 12'h811;
        src75 <= 12'h323;
        src76 <= 12'hd6;
        src77 <= 12'h90d;
        src78 <= 12'ha6d;
        src79 <= 12'hddc;
        src80 <= 12'h8d;
        src81 <= 12'h5d;
        src82 <= 12'hf32;
        src83 <= 12'hd02;
        src84 <= 12'heac;
        src85 <= 12'h183;
        src86 <= 12'h539;
        src87 <= 12'hd54;
        src88 <= 12'h33a;
        src89 <= 12'ha59;
        src90 <= 12'h79c;
        src91 <= 12'hc80;
        src92 <= 12'h61;
        src93 <= 12'hef7;
        src94 <= 12'hbb3;
        src95 <= 12'h8da;
        src96 <= 12'h316;
        src97 <= 12'h634;
        src98 <= 12'h604;
        src99 <= 12'hf3a;
        src100 <= 12'hec5;
        src101 <= 12'ha39;
        src102 <= 12'hcfa;
        src103 <= 12'hf16;
        src104 <= 12'haf0;
        src105 <= 12'h3bf;
        src106 <= 12'hc4b;
        src107 <= 12'h11d;
        src108 <= 12'h295;
        src109 <= 12'h208;
        src110 <= 12'hd3f;
        src111 <= 12'hea5;
        src112 <= 12'hcd1;
        src113 <= 12'h6;
        src114 <= 12'hbb;
        src115 <= 12'h403;
        src116 <= 12'h4bf;
        src117 <= 12'h6e6;
        src118 <= 12'hf55;
        src119 <= 12'hbd3;
        src120 <= 12'h191;
        src121 <= 12'hc8e;
        src122 <= 12'h9aa;
        src123 <= 12'h897;
        src124 <= 12'h3d7;
        src125 <= 12'ha7b;
        src126 <= 12'hc51;
        src127 <= 12'h2f0;
        src128 <= 12'ha8f;
        src129 <= 12'hab0;
        src130 <= 12'hf4c;
        src131 <= 12'h732;
        src132 <= 12'h758;
        src133 <= 12'hdef;
        src134 <= 12'haf6;
        src135 <= 12'haf7;
        src136 <= 12'h774;
        src137 <= 12'hf21;
        src138 <= 12'ha1;
        src139 <= 12'hc1f;
        src140 <= 12'h23b;
        src141 <= 12'h4bd;
        src142 <= 12'hd2f;
        src143 <= 12'h250;
        src144 <= 12'h45d;
        src145 <= 12'h63;
        src146 <= 12'h6e0;
        src147 <= 12'hd82;
        src148 <= 12'h7b3;
        src149 <= 12'ha76;
        src150 <= 12'h388;
        src151 <= 12'ha61;
        src152 <= 12'hc44;
        src153 <= 12'h4fa;
        src154 <= 12'hbeb;
        src155 <= 12'hbd6;
        src156 <= 12'hb61;
        src157 <= 12'hee1;
        src158 <= 12'hdef;
        src159 <= 12'hf65;
        src160 <= 12'hb6d;
        src161 <= 12'h93e;
        src162 <= 12'h1c3;
        src163 <= 12'h409;
        src164 <= 12'h19a;
        src165 <= 12'h3e3;
        src166 <= 12'h406;
        src167 <= 12'h318;
        src168 <= 12'hf01;
        src169 <= 12'hb76;
        src170 <= 12'hc4a;
        src171 <= 12'h567;
        src172 <= 12'hca4;
        src173 <= 12'hc37;
        src174 <= 12'hfd;
        src175 <= 12'h245;
        src176 <= 12'h2fa;
        src177 <= 12'h1fa;
        src178 <= 12'hfd8;
        src179 <= 12'h2b6;
        src180 <= 12'h633;
        src181 <= 12'h24e;
        src182 <= 12'h327;
        src183 <= 12'h247;
        src184 <= 12'hb71;
        src185 <= 12'h62d;
        src186 <= 12'h9ee;
        src187 <= 12'ha28;
        src188 <= 12'hb39;
        exp <= 20'h6069c;
        #1
        src0 <= 12'h5bf;
        src1 <= 12'h87a;
        src2 <= 12'h93f;
        src3 <= 12'h7d6;
        src4 <= 12'h37b;
        src5 <= 12'hf01;
        src6 <= 12'ha78;
        src7 <= 12'hfc4;
        src8 <= 12'h1ec;
        src9 <= 12'h223;
        src10 <= 12'hc88;
        src11 <= 12'hbf0;
        src12 <= 12'h42e;
        src13 <= 12'hd88;
        src14 <= 12'h89b;
        src15 <= 12'h78b;
        src16 <= 12'h9da;
        src17 <= 12'h9d0;
        src18 <= 12'h2ca;
        src19 <= 12'hb25;
        src20 <= 12'h2d8;
        src21 <= 12'h821;
        src22 <= 12'ha7b;
        src23 <= 12'h12b;
        src24 <= 12'hfd3;
        src25 <= 12'h709;
        src26 <= 12'hf71;
        src27 <= 12'h62a;
        src28 <= 12'h2d6;
        src29 <= 12'h2ce;
        src30 <= 12'h494;
        src31 <= 12'ha4e;
        src32 <= 12'he2c;
        src33 <= 12'hf8e;
        src34 <= 12'h87d;
        src35 <= 12'h6cd;
        src36 <= 12'h48;
        src37 <= 12'h4b3;
        src38 <= 12'hbc1;
        src39 <= 12'h5d2;
        src40 <= 12'hc99;
        src41 <= 12'h7d5;
        src42 <= 12'hfea;
        src43 <= 12'hfd1;
        src44 <= 12'hfec;
        src45 <= 12'hcfc;
        src46 <= 12'h207;
        src47 <= 12'h650;
        src48 <= 12'hf97;
        src49 <= 12'h250;
        src50 <= 12'h796;
        src51 <= 12'h91b;
        src52 <= 12'h352;
        src53 <= 12'h9e3;
        src54 <= 12'ha47;
        src55 <= 12'hecd;
        src56 <= 12'h9eb;
        src57 <= 12'h301;
        src58 <= 12'h828;
        src59 <= 12'h2cd;
        src60 <= 12'h90;
        src61 <= 12'h6d5;
        src62 <= 12'hcc4;
        src63 <= 12'hab2;
        src64 <= 12'h124;
        src65 <= 12'h135;
        src66 <= 12'h29;
        src67 <= 12'h21;
        src68 <= 12'h735;
        src69 <= 12'hfa6;
        src70 <= 12'hd71;
        src71 <= 12'h764;
        src72 <= 12'h344;
        src73 <= 12'heea;
        src74 <= 12'h90e;
        src75 <= 12'h863;
        src76 <= 12'h52a;
        src77 <= 12'he12;
        src78 <= 12'hf96;
        src79 <= 12'hb91;
        src80 <= 12'h7fc;
        src81 <= 12'hf45;
        src82 <= 12'he73;
        src83 <= 12'h3ec;
        src84 <= 12'h7b7;
        src85 <= 12'hb24;
        src86 <= 12'ha50;
        src87 <= 12'hc01;
        src88 <= 12'h773;
        src89 <= 12'h957;
        src90 <= 12'h61e;
        src91 <= 12'hc68;
        src92 <= 12'hcb0;
        src93 <= 12'h7ff;
        src94 <= 12'h9ff;
        src95 <= 12'hb24;
        src96 <= 12'hc38;
        src97 <= 12'hd36;
        src98 <= 12'hc23;
        src99 <= 12'h755;
        src100 <= 12'h50;
        src101 <= 12'hfa0;
        src102 <= 12'hbb;
        src103 <= 12'h6cc;
        src104 <= 12'hb3d;
        src105 <= 12'ha34;
        src106 <= 12'h218;
        src107 <= 12'h7df;
        src108 <= 12'h3e4;
        src109 <= 12'h128;
        src110 <= 12'he36;
        src111 <= 12'h2ed;
        src112 <= 12'hda1;
        src113 <= 12'ha0f;
        src114 <= 12'h49e;
        src115 <= 12'haac;
        src116 <= 12'h68f;
        src117 <= 12'hb45;
        src118 <= 12'h358;
        src119 <= 12'h80f;
        src120 <= 12'h993;
        src121 <= 12'h624;
        src122 <= 12'h336;
        src123 <= 12'h719;
        src124 <= 12'hefa;
        src125 <= 12'ha46;
        src126 <= 12'hb39;
        src127 <= 12'h5d4;
        src128 <= 12'haf8;
        src129 <= 12'h827;
        src130 <= 12'hd4f;
        src131 <= 12'hd24;
        src132 <= 12'h732;
        src133 <= 12'h4fd;
        src134 <= 12'h64b;
        src135 <= 12'h412;
        src136 <= 12'hdcc;
        src137 <= 12'h68;
        src138 <= 12'hd0c;
        src139 <= 12'h474;
        src140 <= 12'hc58;
        src141 <= 12'hb2;
        src142 <= 12'h5c3;
        src143 <= 12'hce6;
        src144 <= 12'hbf3;
        src145 <= 12'h424;
        src146 <= 12'h51d;
        src147 <= 12'hfff;
        src148 <= 12'hace;
        src149 <= 12'hd1b;
        src150 <= 12'h6e2;
        src151 <= 12'hcc4;
        src152 <= 12'h767;
        src153 <= 12'h874;
        src154 <= 12'h5;
        src155 <= 12'h748;
        src156 <= 12'hf60;
        src157 <= 12'hc4a;
        src158 <= 12'h236;
        src159 <= 12'h1ab;
        src160 <= 12'h56d;
        src161 <= 12'h381;
        src162 <= 12'hbd9;
        src163 <= 12'h976;
        src164 <= 12'hbda;
        src165 <= 12'h3da;
        src166 <= 12'hec3;
        src167 <= 12'h89;
        src168 <= 12'h657;
        src169 <= 12'he83;
        src170 <= 12'hf37;
        src171 <= 12'h91c;
        src172 <= 12'h42b;
        src173 <= 12'h250;
        src174 <= 12'h40f;
        src175 <= 12'h339;
        src176 <= 12'h796;
        src177 <= 12'h61;
        src178 <= 12'h257;
        src179 <= 12'hdc5;
        src180 <= 12'h467;
        src181 <= 12'h961;
        src182 <= 12'heaa;
        src183 <= 12'h724;
        src184 <= 12'he4a;
        src185 <= 12'hadd;
        src186 <= 12'h806;
        src187 <= 12'hf5b;
        src188 <= 12'h18f;
        exp <= 20'h633db;
        #1
        src0 <= 12'hc2d;
        src1 <= 12'h1f2;
        src2 <= 12'h51a;
        src3 <= 12'hb7d;
        src4 <= 12'h190;
        src5 <= 12'h4d6;
        src6 <= 12'h44f;
        src7 <= 12'he66;
        src8 <= 12'h328;
        src9 <= 12'h31a;
        src10 <= 12'hfc0;
        src11 <= 12'ha07;
        src12 <= 12'hdb6;
        src13 <= 12'h804;
        src14 <= 12'h7b9;
        src15 <= 12'h887;
        src16 <= 12'he24;
        src17 <= 12'h442;
        src18 <= 12'h744;
        src19 <= 12'h652;
        src20 <= 12'h919;
        src21 <= 12'hdda;
        src22 <= 12'hcf1;
        src23 <= 12'h4b8;
        src24 <= 12'he8e;
        src25 <= 12'h543;
        src26 <= 12'hc75;
        src27 <= 12'he73;
        src28 <= 12'ha84;
        src29 <= 12'h1d7;
        src30 <= 12'h48c;
        src31 <= 12'haf0;
        src32 <= 12'hf98;
        src33 <= 12'h5d3;
        src34 <= 12'hf1f;
        src35 <= 12'h85c;
        src36 <= 12'h5f0;
        src37 <= 12'h731;
        src38 <= 12'h2a2;
        src39 <= 12'he91;
        src40 <= 12'h78a;
        src41 <= 12'hed1;
        src42 <= 12'hee1;
        src43 <= 12'h3e8;
        src44 <= 12'he2;
        src45 <= 12'h9d0;
        src46 <= 12'h1c6;
        src47 <= 12'h8ce;
        src48 <= 12'h8d;
        src49 <= 12'hec5;
        src50 <= 12'h94c;
        src51 <= 12'h20;
        src52 <= 12'h678;
        src53 <= 12'h8e7;
        src54 <= 12'h376;
        src55 <= 12'hbc2;
        src56 <= 12'h5c2;
        src57 <= 12'hda4;
        src58 <= 12'he75;
        src59 <= 12'h8d1;
        src60 <= 12'hff8;
        src61 <= 12'h4e;
        src62 <= 12'h6cc;
        src63 <= 12'heb4;
        src64 <= 12'he7;
        src65 <= 12'hf0;
        src66 <= 12'hb9;
        src67 <= 12'h83;
        src68 <= 12'h707;
        src69 <= 12'had4;
        src70 <= 12'hb65;
        src71 <= 12'h6d4;
        src72 <= 12'h523;
        src73 <= 12'hfc9;
        src74 <= 12'hf80;
        src75 <= 12'hec8;
        src76 <= 12'hf53;
        src77 <= 12'h89;
        src78 <= 12'hce2;
        src79 <= 12'h479;
        src80 <= 12'hbf4;
        src81 <= 12'h99e;
        src82 <= 12'hb9d;
        src83 <= 12'hef6;
        src84 <= 12'h358;
        src85 <= 12'h2b;
        src86 <= 12'h96b;
        src87 <= 12'h93d;
        src88 <= 12'he13;
        src89 <= 12'hf62;
        src90 <= 12'h32e;
        src91 <= 12'h199;
        src92 <= 12'he8d;
        src93 <= 12'ha1f;
        src94 <= 12'ha45;
        src95 <= 12'h196;
        src96 <= 12'hd2b;
        src97 <= 12'h93c;
        src98 <= 12'h4e6;
        src99 <= 12'h971;
        src100 <= 12'h58b;
        src101 <= 12'h3fe;
        src102 <= 12'hef7;
        src103 <= 12'h439;
        src104 <= 12'ha78;
        src105 <= 12'hb20;
        src106 <= 12'h2ce;
        src107 <= 12'h2eb;
        src108 <= 12'h14d;
        src109 <= 12'h3a4;
        src110 <= 12'hc0e;
        src111 <= 12'h6fd;
        src112 <= 12'h49b;
        src113 <= 12'h3b5;
        src114 <= 12'ha6b;
        src115 <= 12'h9f5;
        src116 <= 12'he6c;
        src117 <= 12'hcbb;
        src118 <= 12'h4fc;
        src119 <= 12'h281;
        src120 <= 12'h131;
        src121 <= 12'h3e9;
        src122 <= 12'hcf4;
        src123 <= 12'h45c;
        src124 <= 12'hff4;
        src125 <= 12'hc50;
        src126 <= 12'h73;
        src127 <= 12'he3d;
        src128 <= 12'h918;
        src129 <= 12'hb89;
        src130 <= 12'h7aa;
        src131 <= 12'hd46;
        src132 <= 12'h65c;
        src133 <= 12'h331;
        src134 <= 12'hb31;
        src135 <= 12'hfcb;
        src136 <= 12'hc0b;
        src137 <= 12'hf43;
        src138 <= 12'h69c;
        src139 <= 12'h676;
        src140 <= 12'hbef;
        src141 <= 12'hc27;
        src142 <= 12'h1cf;
        src143 <= 12'h2be;
        src144 <= 12'hd7f;
        src145 <= 12'ha4c;
        src146 <= 12'h736;
        src147 <= 12'hf01;
        src148 <= 12'h89;
        src149 <= 12'h10b;
        src150 <= 12'h7c2;
        src151 <= 12'h5de;
        src152 <= 12'hfda;
        src153 <= 12'h10e;
        src154 <= 12'h7e2;
        src155 <= 12'hf63;
        src156 <= 12'hb68;
        src157 <= 12'h431;
        src158 <= 12'h44c;
        src159 <= 12'h96e;
        src160 <= 12'he2e;
        src161 <= 12'h9fa;
        src162 <= 12'h958;
        src163 <= 12'heb7;
        src164 <= 12'h9da;
        src165 <= 12'h452;
        src166 <= 12'hfb3;
        src167 <= 12'hebe;
        src168 <= 12'ha67;
        src169 <= 12'hdee;
        src170 <= 12'h584;
        src171 <= 12'h477;
        src172 <= 12'h1f0;
        src173 <= 12'ha0d;
        src174 <= 12'h899;
        src175 <= 12'hbcc;
        src176 <= 12'hc56;
        src177 <= 12'hb39;
        src178 <= 12'hfcc;
        src179 <= 12'h5ed;
        src180 <= 12'he53;
        src181 <= 12'h79f;
        src182 <= 12'h7c8;
        src183 <= 12'hdf4;
        src184 <= 12'he00;
        src185 <= 12'h5aa;
        src186 <= 12'h26c;
        src187 <= 12'h2ad;
        src188 <= 12'hd70;
        exp <= 20'h65504;
        #1
        src0 <= 12'h1b6;
        src1 <= 12'hbb1;
        src2 <= 12'hd5f;
        src3 <= 12'h5ef;
        src4 <= 12'h592;
        src5 <= 12'hd80;
        src6 <= 12'h34e;
        src7 <= 12'hc1a;
        src8 <= 12'h333;
        src9 <= 12'h658;
        src10 <= 12'h6ea;
        src11 <= 12'hadb;
        src12 <= 12'h736;
        src13 <= 12'h8c6;
        src14 <= 12'h83d;
        src15 <= 12'h186;
        src16 <= 12'h577;
        src17 <= 12'h99b;
        src18 <= 12'h140;
        src19 <= 12'h858;
        src20 <= 12'h5e1;
        src21 <= 12'hd56;
        src22 <= 12'h67c;
        src23 <= 12'h544;
        src24 <= 12'h619;
        src25 <= 12'hfb3;
        src26 <= 12'hed6;
        src27 <= 12'hcd2;
        src28 <= 12'hdbc;
        src29 <= 12'h443;
        src30 <= 12'hf05;
        src31 <= 12'h9bb;
        src32 <= 12'h7a2;
        src33 <= 12'he09;
        src34 <= 12'he6e;
        src35 <= 12'h4ac;
        src36 <= 12'ha74;
        src37 <= 12'h1af;
        src38 <= 12'he42;
        src39 <= 12'h752;
        src40 <= 12'ha61;
        src41 <= 12'hed0;
        src42 <= 12'h4d7;
        src43 <= 12'h469;
        src44 <= 12'h5c3;
        src45 <= 12'hf55;
        src46 <= 12'h14;
        src47 <= 12'heb8;
        src48 <= 12'h151;
        src49 <= 12'h331;
        src50 <= 12'h89f;
        src51 <= 12'h503;
        src52 <= 12'h719;
        src53 <= 12'h868;
        src54 <= 12'h538;
        src55 <= 12'hce5;
        src56 <= 12'h21e;
        src57 <= 12'h780;
        src58 <= 12'hf30;
        src59 <= 12'h18;
        src60 <= 12'hff4;
        src61 <= 12'h137;
        src62 <= 12'h28a;
        src63 <= 12'hed7;
        src64 <= 12'h851;
        src65 <= 12'h858;
        src66 <= 12'h45f;
        src67 <= 12'ha64;
        src68 <= 12'hf7f;
        src69 <= 12'hc59;
        src70 <= 12'h1b4;
        src71 <= 12'h4cb;
        src72 <= 12'heb0;
        src73 <= 12'h729;
        src74 <= 12'h946;
        src75 <= 12'haa7;
        src76 <= 12'h5d0;
        src77 <= 12'h19b;
        src78 <= 12'h385;
        src79 <= 12'hee0;
        src80 <= 12'hce8;
        src81 <= 12'h975;
        src82 <= 12'h17f;
        src83 <= 12'h457;
        src84 <= 12'hbb;
        src85 <= 12'hf18;
        src86 <= 12'h6e1;
        src87 <= 12'h6fc;
        src88 <= 12'h9ea;
        src89 <= 12'h889;
        src90 <= 12'hef4;
        src91 <= 12'he77;
        src92 <= 12'h2ce;
        src93 <= 12'hd15;
        src94 <= 12'he84;
        src95 <= 12'had7;
        src96 <= 12'h1c7;
        src97 <= 12'h487;
        src98 <= 12'h902;
        src99 <= 12'h54e;
        src100 <= 12'h962;
        src101 <= 12'haa6;
        src102 <= 12'hea2;
        src103 <= 12'h1c9;
        src104 <= 12'hd1d;
        src105 <= 12'hdab;
        src106 <= 12'he7;
        src107 <= 12'h513;
        src108 <= 12'hfcf;
        src109 <= 12'he59;
        src110 <= 12'h98f;
        src111 <= 12'h17e;
        src112 <= 12'h6bc;
        src113 <= 12'h370;
        src114 <= 12'h259;
        src115 <= 12'h786;
        src116 <= 12'he28;
        src117 <= 12'hea9;
        src118 <= 12'h509;
        src119 <= 12'h5da;
        src120 <= 12'h39;
        src121 <= 12'h89f;
        src122 <= 12'h63b;
        src123 <= 12'hf06;
        src124 <= 12'h5f;
        src125 <= 12'hc2a;
        src126 <= 12'ha8d;
        src127 <= 12'h31b;
        src128 <= 12'h9b5;
        src129 <= 12'h48d;
        src130 <= 12'h1a9;
        src131 <= 12'h322;
        src132 <= 12'hc7;
        src133 <= 12'h5fc;
        src134 <= 12'h488;
        src135 <= 12'had3;
        src136 <= 12'h392;
        src137 <= 12'h387;
        src138 <= 12'heca;
        src139 <= 12'h77b;
        src140 <= 12'h90c;
        src141 <= 12'hdac;
        src142 <= 12'h465;
        src143 <= 12'hfe6;
        src144 <= 12'hcfb;
        src145 <= 12'he1f;
        src146 <= 12'hb4d;
        src147 <= 12'haa2;
        src148 <= 12'hcb6;
        src149 <= 12'h3f6;
        src150 <= 12'h21b;
        src151 <= 12'hab8;
        src152 <= 12'h9c2;
        src153 <= 12'hb6b;
        src154 <= 12'h690;
        src155 <= 12'h810;
        src156 <= 12'h6a7;
        src157 <= 12'he16;
        src158 <= 12'h524;
        src159 <= 12'h6c7;
        src160 <= 12'h396;
        src161 <= 12'hecd;
        src162 <= 12'h541;
        src163 <= 12'h450;
        src164 <= 12'ha06;
        src165 <= 12'hd82;
        src166 <= 12'h8e8;
        src167 <= 12'h1cb;
        src168 <= 12'hd6;
        src169 <= 12'h9ef;
        src170 <= 12'h22f;
        src171 <= 12'hf3b;
        src172 <= 12'h71b;
        src173 <= 12'h546;
        src174 <= 12'h4dd;
        src175 <= 12'h266;
        src176 <= 12'hc02;
        src177 <= 12'hafe;
        src178 <= 12'hec1;
        src179 <= 12'h43d;
        src180 <= 12'h125;
        src181 <= 12'h7df;
        src182 <= 12'h1f6;
        src183 <= 12'h45a;
        src184 <= 12'h9bb;
        src185 <= 12'hca;
        src186 <= 12'h1b9;
        src187 <= 12'h1af;
        src188 <= 12'h19f;
        exp <= 20'h5d6e9;
        #1
        src0 <= 12'h6f4;
        src1 <= 12'hf68;
        src2 <= 12'hf3f;
        src3 <= 12'h215;
        src4 <= 12'h303;
        src5 <= 12'hb1b;
        src6 <= 12'h304;
        src7 <= 12'hc1a;
        src8 <= 12'hecd;
        src9 <= 12'h112;
        src10 <= 12'h68a;
        src11 <= 12'h539;
        src12 <= 12'h3f8;
        src13 <= 12'h112;
        src14 <= 12'ha8d;
        src15 <= 12'hfb7;
        src16 <= 12'had6;
        src17 <= 12'hcc3;
        src18 <= 12'h6d;
        src19 <= 12'hac7;
        src20 <= 12'h5bc;
        src21 <= 12'h1b5;
        src22 <= 12'hf53;
        src23 <= 12'h7f6;
        src24 <= 12'hbbd;
        src25 <= 12'h983;
        src26 <= 12'h3a0;
        src27 <= 12'h183;
        src28 <= 12'h9d;
        src29 <= 12'hce0;
        src30 <= 12'h5a;
        src31 <= 12'h65c;
        src32 <= 12'h5e1;
        src33 <= 12'h66e;
        src34 <= 12'h784;
        src35 <= 12'hfbf;
        src36 <= 12'hbf0;
        src37 <= 12'hd1;
        src38 <= 12'hf56;
        src39 <= 12'hd72;
        src40 <= 12'h25a;
        src41 <= 12'h9a2;
        src42 <= 12'h915;
        src43 <= 12'h36f;
        src44 <= 12'h174;
        src45 <= 12'hd12;
        src46 <= 12'h4a5;
        src47 <= 12'h5c0;
        src48 <= 12'hd2f;
        src49 <= 12'hb55;
        src50 <= 12'hff8;
        src51 <= 12'h87a;
        src52 <= 12'h289;
        src53 <= 12'h8c6;
        src54 <= 12'h415;
        src55 <= 12'h9f2;
        src56 <= 12'h49f;
        src57 <= 12'h65a;
        src58 <= 12'h144;
        src59 <= 12'h76e;
        src60 <= 12'h7b3;
        src61 <= 12'hc9e;
        src62 <= 12'hf5e;
        src63 <= 12'h1b3;
        src64 <= 12'h5cf;
        src65 <= 12'h556;
        src66 <= 12'h6c7;
        src67 <= 12'h30c;
        src68 <= 12'h5fc;
        src69 <= 12'hb09;
        src70 <= 12'h9c2;
        src71 <= 12'h303;
        src72 <= 12'h7ee;
        src73 <= 12'hf82;
        src74 <= 12'h35e;
        src75 <= 12'he1c;
        src76 <= 12'hea4;
        src77 <= 12'hd97;
        src78 <= 12'h5fd;
        src79 <= 12'h299;
        src80 <= 12'ha72;
        src81 <= 12'h9bf;
        src82 <= 12'h482;
        src83 <= 12'hb56;
        src84 <= 12'h6de;
        src85 <= 12'hc5d;
        src86 <= 12'h908;
        src87 <= 12'haab;
        src88 <= 12'h706;
        src89 <= 12'h4a3;
        src90 <= 12'ha45;
        src91 <= 12'h581;
        src92 <= 12'h392;
        src93 <= 12'hc9;
        src94 <= 12'haae;
        src95 <= 12'h8cf;
        src96 <= 12'hb66;
        src97 <= 12'h89b;
        src98 <= 12'hb04;
        src99 <= 12'h92c;
        src100 <= 12'hbe9;
        src101 <= 12'h822;
        src102 <= 12'h850;
        src103 <= 12'hd2;
        src104 <= 12'h990;
        src105 <= 12'hd86;
        src106 <= 12'h668;
        src107 <= 12'hfcb;
        src108 <= 12'h2e6;
        src109 <= 12'h3a8;
        src110 <= 12'h88a;
        src111 <= 12'h17e;
        src112 <= 12'h5ba;
        src113 <= 12'hfe6;
        src114 <= 12'h84a;
        src115 <= 12'h52d;
        src116 <= 12'hc2e;
        src117 <= 12'hbd5;
        src118 <= 12'h3e0;
        src119 <= 12'h21c;
        src120 <= 12'h6fa;
        src121 <= 12'haa2;
        src122 <= 12'h1b1;
        src123 <= 12'h71;
        src124 <= 12'h38f;
        src125 <= 12'hfac;
        src126 <= 12'h34d;
        src127 <= 12'h212;
        src128 <= 12'h777;
        src129 <= 12'he99;
        src130 <= 12'h981;
        src131 <= 12'h9de;
        src132 <= 12'hcab;
        src133 <= 12'h740;
        src134 <= 12'h823;
        src135 <= 12'ha15;
        src136 <= 12'h37a;
        src137 <= 12'h36f;
        src138 <= 12'hb62;
        src139 <= 12'hbea;
        src140 <= 12'h20a;
        src141 <= 12'h554;
        src142 <= 12'hdc8;
        src143 <= 12'h4bb;
        src144 <= 12'h5bc;
        src145 <= 12'h7e6;
        src146 <= 12'hd47;
        src147 <= 12'h6c2;
        src148 <= 12'h449;
        src149 <= 12'h5ee;
        src150 <= 12'ha2f;
        src151 <= 12'h4f2;
        src152 <= 12'h947;
        src153 <= 12'h671;
        src154 <= 12'h72d;
        src155 <= 12'h24a;
        src156 <= 12'h9dc;
        src157 <= 12'hf7;
        src158 <= 12'h25;
        src159 <= 12'h645;
        src160 <= 12'h769;
        src161 <= 12'he7e;
        src162 <= 12'hdbc;
        src163 <= 12'hd0b;
        src164 <= 12'h363;
        src165 <= 12'hc2a;
        src166 <= 12'he26;
        src167 <= 12'h49f;
        src168 <= 12'hcf9;
        src169 <= 12'hcb;
        src170 <= 12'h2c1;
        src171 <= 12'hc31;
        src172 <= 12'h805;
        src173 <= 12'h32f;
        src174 <= 12'h32d;
        src175 <= 12'h623;
        src176 <= 12'ha53;
        src177 <= 12'ha9f;
        src178 <= 12'hee9;
        src179 <= 12'hbf;
        src180 <= 12'h8b2;
        src181 <= 12'h79c;
        src182 <= 12'h1e7;
        src183 <= 12'h48;
        src184 <= 12'hd2b;
        src185 <= 12'hf0;
        src186 <= 12'hab0;
        src187 <= 12'hc38;
        src188 <= 12'hbd3;
        exp <= 20'h5ba7c;
        #1
        src0 <= 12'h5ae;
        src1 <= 12'h843;
        src2 <= 12'hdbc;
        src3 <= 12'h24a;
        src4 <= 12'h6db;
        src5 <= 12'h9e;
        src6 <= 12'h33a;
        src7 <= 12'h289;
        src8 <= 12'hc0e;
        src9 <= 12'he98;
        src10 <= 12'hdc1;
        src11 <= 12'h5ec;
        src12 <= 12'h618;
        src13 <= 12'hdaa;
        src14 <= 12'h939;
        src15 <= 12'hc35;
        src16 <= 12'h80a;
        src17 <= 12'h43b;
        src18 <= 12'h674;
        src19 <= 12'h752;
        src20 <= 12'h9b6;
        src21 <= 12'hc9f;
        src22 <= 12'h9cd;
        src23 <= 12'h27a;
        src24 <= 12'ha6a;
        src25 <= 12'hb9c;
        src26 <= 12'h57;
        src27 <= 12'he0e;
        src28 <= 12'hbc0;
        src29 <= 12'hf42;
        src30 <= 12'h5b2;
        src31 <= 12'hab1;
        src32 <= 12'h18f;
        src33 <= 12'hc6e;
        src34 <= 12'h20a;
        src35 <= 12'h738;
        src36 <= 12'hd36;
        src37 <= 12'hc88;
        src38 <= 12'h7ac;
        src39 <= 12'he3d;
        src40 <= 12'h3cd;
        src41 <= 12'h7b2;
        src42 <= 12'h8a0;
        src43 <= 12'h542;
        src44 <= 12'hb2c;
        src45 <= 12'hb45;
        src46 <= 12'h850;
        src47 <= 12'he7a;
        src48 <= 12'he9c;
        src49 <= 12'h53d;
        src50 <= 12'h24a;
        src51 <= 12'h8a2;
        src52 <= 12'he40;
        src53 <= 12'hecd;
        src54 <= 12'h937;
        src55 <= 12'hdd4;
        src56 <= 12'hea1;
        src57 <= 12'h394;
        src58 <= 12'hb49;
        src59 <= 12'hf6;
        src60 <= 12'h9d0;
        src61 <= 12'hdb;
        src62 <= 12'h512;
        src63 <= 12'h4e4;
        src64 <= 12'h730;
        src65 <= 12'h980;
        src66 <= 12'h524;
        src67 <= 12'h569;
        src68 <= 12'h6c6;
        src69 <= 12'h8f1;
        src70 <= 12'h4cd;
        src71 <= 12'hce0;
        src72 <= 12'hfde;
        src73 <= 12'h882;
        src74 <= 12'hf95;
        src75 <= 12'hfa5;
        src76 <= 12'ha3a;
        src77 <= 12'h642;
        src78 <= 12'h55c;
        src79 <= 12'h443;
        src80 <= 12'h71a;
        src81 <= 12'h4f9;
        src82 <= 12'h973;
        src83 <= 12'h897;
        src84 <= 12'h75;
        src85 <= 12'h713;
        src86 <= 12'ha32;
        src87 <= 12'hb1a;
        src88 <= 12'h989;
        src89 <= 12'h17f;
        src90 <= 12'hb8;
        src91 <= 12'h2a7;
        src92 <= 12'hfc2;
        src93 <= 12'h1e8;
        src94 <= 12'h56a;
        src95 <= 12'h82;
        src96 <= 12'hb1d;
        src97 <= 12'h665;
        src98 <= 12'h16e;
        src99 <= 12'he0d;
        src100 <= 12'h6b2;
        src101 <= 12'h1e7;
        src102 <= 12'h167;
        src103 <= 12'hf71;
        src104 <= 12'h29e;
        src105 <= 12'h318;
        src106 <= 12'h41e;
        src107 <= 12'hc6c;
        src108 <= 12'h623;
        src109 <= 12'hfbf;
        src110 <= 12'hab6;
        src111 <= 12'hb90;
        src112 <= 12'hfb;
        src113 <= 12'h75;
        src114 <= 12'h71c;
        src115 <= 12'hfef;
        src116 <= 12'hdd7;
        src117 <= 12'h314;
        src118 <= 12'h461;
        src119 <= 12'he4c;
        src120 <= 12'had1;
        src121 <= 12'hdb5;
        src122 <= 12'h8f6;
        src123 <= 12'hb58;
        src124 <= 12'h6a6;
        src125 <= 12'h186;
        src126 <= 12'h84;
        src127 <= 12'h144;
        src128 <= 12'h6ce;
        src129 <= 12'hc97;
        src130 <= 12'hefe;
        src131 <= 12'h93e;
        src132 <= 12'h364;
        src133 <= 12'haa2;
        src134 <= 12'h87;
        src135 <= 12'h978;
        src136 <= 12'hc8c;
        src137 <= 12'h6a6;
        src138 <= 12'h196;
        src139 <= 12'h1ef;
        src140 <= 12'h933;
        src141 <= 12'hc1c;
        src142 <= 12'hc4d;
        src143 <= 12'h48d;
        src144 <= 12'hf40;
        src145 <= 12'hbf2;
        src146 <= 12'hf80;
        src147 <= 12'hee7;
        src148 <= 12'hb32;
        src149 <= 12'h736;
        src150 <= 12'h767;
        src151 <= 12'hcaf;
        src152 <= 12'hdd8;
        src153 <= 12'hded;
        src154 <= 12'h4e7;
        src155 <= 12'h3ec;
        src156 <= 12'hd21;
        src157 <= 12'h353;
        src158 <= 12'h984;
        src159 <= 12'h826;
        src160 <= 12'h81e;
        src161 <= 12'hc1d;
        src162 <= 12'hb9;
        src163 <= 12'hfbe;
        src164 <= 12'hc6b;
        src165 <= 12'hd77;
        src166 <= 12'hce1;
        src167 <= 12'h198;
        src168 <= 12'he9;
        src169 <= 12'h4;
        src170 <= 12'h6b7;
        src171 <= 12'h2e4;
        src172 <= 12'h977;
        src173 <= 12'hce1;
        src174 <= 12'h7a2;
        src175 <= 12'hc85;
        src176 <= 12'h312;
        src177 <= 12'hde6;
        src178 <= 12'h40d;
        src179 <= 12'hd81;
        src180 <= 12'hf50;
        src181 <= 12'h1a8;
        src182 <= 12'hdcd;
        src183 <= 12'h94;
        src184 <= 12'h640;
        src185 <= 12'h8c0;
        src186 <= 12'h92a;
        src187 <= 12'h79;
        src188 <= 12'hc44;
        exp <= 20'h611c3;
        #1
        src0 <= 12'h3d2;
        src1 <= 12'he1c;
        src2 <= 12'h472;
        src3 <= 12'h9c5;
        src4 <= 12'h5c4;
        src5 <= 12'h229;
        src6 <= 12'hee9;
        src7 <= 12'hd72;
        src8 <= 12'h6d;
        src9 <= 12'h35b;
        src10 <= 12'h798;
        src11 <= 12'hac8;
        src12 <= 12'heab;
        src13 <= 12'hce9;
        src14 <= 12'h19a;
        src15 <= 12'ha96;
        src16 <= 12'hc78;
        src17 <= 12'h579;
        src18 <= 12'ha6;
        src19 <= 12'hc0b;
        src20 <= 12'h289;
        src21 <= 12'h742;
        src22 <= 12'hb84;
        src23 <= 12'hf18;
        src24 <= 12'h1b8;
        src25 <= 12'h558;
        src26 <= 12'h892;
        src27 <= 12'h164;
        src28 <= 12'h4d;
        src29 <= 12'h720;
        src30 <= 12'hce8;
        src31 <= 12'h72c;
        src32 <= 12'hd95;
        src33 <= 12'he4d;
        src34 <= 12'h119;
        src35 <= 12'hffb;
        src36 <= 12'hbf7;
        src37 <= 12'h4eb;
        src38 <= 12'hbab;
        src39 <= 12'he03;
        src40 <= 12'h8af;
        src41 <= 12'hbf0;
        src42 <= 12'h749;
        src43 <= 12'h3b6;
        src44 <= 12'h51;
        src45 <= 12'h2cd;
        src46 <= 12'ha2b;
        src47 <= 12'hdad;
        src48 <= 12'ha5c;
        src49 <= 12'hf81;
        src50 <= 12'h3e4;
        src51 <= 12'hfd8;
        src52 <= 12'h8c6;
        src53 <= 12'h438;
        src54 <= 12'h3ef;
        src55 <= 12'hbf6;
        src56 <= 12'hd49;
        src57 <= 12'hc9f;
        src58 <= 12'hd20;
        src59 <= 12'hb1;
        src60 <= 12'hcf;
        src61 <= 12'h7f0;
        src62 <= 12'hf25;
        src63 <= 12'h9a1;
        src64 <= 12'hc5;
        src65 <= 12'h4a3;
        src66 <= 12'h927;
        src67 <= 12'hae1;
        src68 <= 12'h977;
        src69 <= 12'hbab;
        src70 <= 12'ha7f;
        src71 <= 12'hb13;
        src72 <= 12'hecf;
        src73 <= 12'h174;
        src74 <= 12'h59c;
        src75 <= 12'hdbc;
        src76 <= 12'h140;
        src77 <= 12'he9c;
        src78 <= 12'h3de;
        src79 <= 12'h7ef;
        src80 <= 12'h80f;
        src81 <= 12'hd3e;
        src82 <= 12'h87f;
        src83 <= 12'h715;
        src84 <= 12'ha8f;
        src85 <= 12'h678;
        src86 <= 12'h5be;
        src87 <= 12'h58e;
        src88 <= 12'hbb9;
        src89 <= 12'h4f2;
        src90 <= 12'h266;
        src91 <= 12'h4cf;
        src92 <= 12'h788;
        src93 <= 12'h50d;
        src94 <= 12'haef;
        src95 <= 12'h416;
        src96 <= 12'h17e;
        src97 <= 12'h29c;
        src98 <= 12'h3e3;
        src99 <= 12'ha79;
        src100 <= 12'he0d;
        src101 <= 12'hf71;
        src102 <= 12'hbdc;
        src103 <= 12'h9ef;
        src104 <= 12'h848;
        src105 <= 12'h3eb;
        src106 <= 12'hd4d;
        src107 <= 12'h6eb;
        src108 <= 12'h1f4;
        src109 <= 12'hc6;
        src110 <= 12'hf41;
        src111 <= 12'h502;
        src112 <= 12'h26d;
        src113 <= 12'h188;
        src114 <= 12'h937;
        src115 <= 12'hee1;
        src116 <= 12'h226;
        src117 <= 12'h4db;
        src118 <= 12'h8f1;
        src119 <= 12'h873;
        src120 <= 12'h742;
        src121 <= 12'h931;
        src122 <= 12'h35a;
        src123 <= 12'h301;
        src124 <= 12'ha14;
        src125 <= 12'hb48;
        src126 <= 12'h68a;
        src127 <= 12'ha3d;
        src128 <= 12'he24;
        src129 <= 12'h8f3;
        src130 <= 12'h4f4;
        src131 <= 12'h4de;
        src132 <= 12'hd51;
        src133 <= 12'hfbe;
        src134 <= 12'hd13;
        src135 <= 12'h453;
        src136 <= 12'h93d;
        src137 <= 12'hbf9;
        src138 <= 12'h3c2;
        src139 <= 12'hf91;
        src140 <= 12'hc71;
        src141 <= 12'he2f;
        src142 <= 12'hf62;
        src143 <= 12'h2dd;
        src144 <= 12'h351;
        src145 <= 12'hf5c;
        src146 <= 12'he75;
        src147 <= 12'h262;
        src148 <= 12'hbc5;
        src149 <= 12'h937;
        src150 <= 12'h712;
        src151 <= 12'hb7c;
        src152 <= 12'hb4e;
        src153 <= 12'hed6;
        src154 <= 12'h4e7;
        src155 <= 12'h3c8;
        src156 <= 12'hbb9;
        src157 <= 12'h12f;
        src158 <= 12'h1e4;
        src159 <= 12'h2a4;
        src160 <= 12'hdf8;
        src161 <= 12'h1bd;
        src162 <= 12'h64a;
        src163 <= 12'h935;
        src164 <= 12'h1a2;
        src165 <= 12'h7b8;
        src166 <= 12'h4f6;
        src167 <= 12'h3c3;
        src168 <= 12'h232;
        src169 <= 12'hc9b;
        src170 <= 12'hda;
        src171 <= 12'hc00;
        src172 <= 12'hc18;
        src173 <= 12'hccb;
        src174 <= 12'h687;
        src175 <= 12'h397;
        src176 <= 12'h7fb;
        src177 <= 12'h38c;
        src178 <= 12'h1cc;
        src179 <= 12'hddd;
        src180 <= 12'h584;
        src181 <= 12'hab6;
        src182 <= 12'h243;
        src183 <= 12'hc3b;
        src184 <= 12'hd75;
        src185 <= 12'he05;
        src186 <= 12'h6a9;
        src187 <= 12'h911;
        src188 <= 12'h602;
        exp <= 20'h5fd81;
        #1
        src0 <= 12'ha19;
        src1 <= 12'had9;
        src2 <= 12'h1db;
        src3 <= 12'h6c9;
        src4 <= 12'h29e;
        src5 <= 12'hac2;
        src6 <= 12'ha0f;
        src7 <= 12'hd05;
        src8 <= 12'h14f;
        src9 <= 12'h132;
        src10 <= 12'hf9b;
        src11 <= 12'hc82;
        src12 <= 12'h1c2;
        src13 <= 12'hfbe;
        src14 <= 12'hc7d;
        src15 <= 12'hfc4;
        src16 <= 12'hb00;
        src17 <= 12'ha6e;
        src18 <= 12'hf90;
        src19 <= 12'h7cc;
        src20 <= 12'haa1;
        src21 <= 12'he28;
        src22 <= 12'h8ce;
        src23 <= 12'h300;
        src24 <= 12'h6dd;
        src25 <= 12'h68;
        src26 <= 12'h3e1;
        src27 <= 12'h101;
        src28 <= 12'h744;
        src29 <= 12'hcec;
        src30 <= 12'h590;
        src31 <= 12'h759;
        src32 <= 12'h820;
        src33 <= 12'he76;
        src34 <= 12'he3c;
        src35 <= 12'he02;
        src36 <= 12'h440;
        src37 <= 12'hf8b;
        src38 <= 12'he5;
        src39 <= 12'h453;
        src40 <= 12'hc24;
        src41 <= 12'h83a;
        src42 <= 12'hd9;
        src43 <= 12'hf8e;
        src44 <= 12'hd24;
        src45 <= 12'hce9;
        src46 <= 12'h9d5;
        src47 <= 12'h27b;
        src48 <= 12'h2a7;
        src49 <= 12'hf7e;
        src50 <= 12'h279;
        src51 <= 12'ha0c;
        src52 <= 12'hdc9;
        src53 <= 12'h65a;
        src54 <= 12'ha20;
        src55 <= 12'h157;
        src56 <= 12'hf8b;
        src57 <= 12'h2f1;
        src58 <= 12'hd9d;
        src59 <= 12'h65f;
        src60 <= 12'h7ff;
        src61 <= 12'h1f2;
        src62 <= 12'hd58;
        src63 <= 12'h2af;
        src64 <= 12'hf26;
        src65 <= 12'hd54;
        src66 <= 12'h6f0;
        src67 <= 12'h7ed;
        src68 <= 12'hf6a;
        src69 <= 12'h673;
        src70 <= 12'h2cf;
        src71 <= 12'h9a0;
        src72 <= 12'h2e;
        src73 <= 12'h2af;
        src74 <= 12'he8d;
        src75 <= 12'heb0;
        src76 <= 12'h1c8;
        src77 <= 12'h38e;
        src78 <= 12'h104;
        src79 <= 12'ha68;
        src80 <= 12'hcd7;
        src81 <= 12'h95d;
        src82 <= 12'h762;
        src83 <= 12'h3e6;
        src84 <= 12'hb8a;
        src85 <= 12'hdc5;
        src86 <= 12'hf58;
        src87 <= 12'h5d8;
        src88 <= 12'h4f3;
        src89 <= 12'h777;
        src90 <= 12'had0;
        src91 <= 12'ha93;
        src92 <= 12'h67a;
        src93 <= 12'hba;
        src94 <= 12'h8c8;
        src95 <= 12'h83e;
        src96 <= 12'h4f;
        src97 <= 12'hc54;
        src98 <= 12'h494;
        src99 <= 12'hcc1;
        src100 <= 12'h834;
        src101 <= 12'hf40;
        src102 <= 12'h86f;
        src103 <= 12'hbfa;
        src104 <= 12'h358;
        src105 <= 12'h3f4;
        src106 <= 12'ha04;
        src107 <= 12'h3a3;
        src108 <= 12'h2be;
        src109 <= 12'hce2;
        src110 <= 12'h38a;
        src111 <= 12'hb0a;
        src112 <= 12'h709;
        src113 <= 12'h14b;
        src114 <= 12'h22a;
        src115 <= 12'h231;
        src116 <= 12'h657;
        src117 <= 12'h554;
        src118 <= 12'h2cd;
        src119 <= 12'hd66;
        src120 <= 12'hd2c;
        src121 <= 12'ha7a;
        src122 <= 12'hdb;
        src123 <= 12'h972;
        src124 <= 12'h55e;
        src125 <= 12'hc8a;
        src126 <= 12'h653;
        src127 <= 12'h7f2;
        src128 <= 12'h29a;
        src129 <= 12'h962;
        src130 <= 12'h3bb;
        src131 <= 12'h6dc;
        src132 <= 12'h48b;
        src133 <= 12'h602;
        src134 <= 12'h9e4;
        src135 <= 12'hb2b;
        src136 <= 12'h3f4;
        src137 <= 12'hf49;
        src138 <= 12'hd9;
        src139 <= 12'h22a;
        src140 <= 12'h8de;
        src141 <= 12'hd23;
        src142 <= 12'he75;
        src143 <= 12'h13e;
        src144 <= 12'hf0;
        src145 <= 12'he1;
        src146 <= 12'hb28;
        src147 <= 12'hd03;
        src148 <= 12'h4c4;
        src149 <= 12'h80d;
        src150 <= 12'hd7d;
        src151 <= 12'h6ac;
        src152 <= 12'h18d;
        src153 <= 12'h6d4;
        src154 <= 12'ha50;
        src155 <= 12'h1f4;
        src156 <= 12'h2c7;
        src157 <= 12'habd;
        src158 <= 12'hf2;
        src159 <= 12'h196;
        src160 <= 12'hdcd;
        src161 <= 12'hade;
        src162 <= 12'ha50;
        src163 <= 12'h851;
        src164 <= 12'h92c;
        src165 <= 12'h496;
        src166 <= 12'h11c;
        src167 <= 12'hbf6;
        src168 <= 12'hbed;
        src169 <= 12'hed9;
        src170 <= 12'h6cc;
        src171 <= 12'h3de;
        src172 <= 12'h711;
        src173 <= 12'h4eb;
        src174 <= 12'hd09;
        src175 <= 12'ha84;
        src176 <= 12'h164;
        src177 <= 12'hd52;
        src178 <= 12'h9ce;
        src179 <= 12'ha9c;
        src180 <= 12'hc88;
        src181 <= 12'ha67;
        src182 <= 12'hdef;
        src183 <= 12'he64;
        src184 <= 12'h540;
        src185 <= 12'h2c6;
        src186 <= 12'h96a;
        src187 <= 12'hdec;
        src188 <= 12'h121;
        exp <= 20'h5eaa3;
        #1
        src0 <= 12'hec9;
        src1 <= 12'h526;
        src2 <= 12'h830;
        src3 <= 12'hd2c;
        src4 <= 12'hc1d;
        src5 <= 12'h3a7;
        src6 <= 12'ha7c;
        src7 <= 12'hea9;
        src8 <= 12'h351;
        src9 <= 12'h5de;
        src10 <= 12'hc32;
        src11 <= 12'h629;
        src12 <= 12'h6d7;
        src13 <= 12'hdb6;
        src14 <= 12'hc6f;
        src15 <= 12'h524;
        src16 <= 12'h71d;
        src17 <= 12'h7ba;
        src18 <= 12'ha5f;
        src19 <= 12'haee;
        src20 <= 12'haa5;
        src21 <= 12'ha46;
        src22 <= 12'hc02;
        src23 <= 12'hcd1;
        src24 <= 12'h7c3;
        src25 <= 12'h8c1;
        src26 <= 12'h108;
        src27 <= 12'h38b;
        src28 <= 12'h595;
        src29 <= 12'h659;
        src30 <= 12'h598;
        src31 <= 12'h6ea;
        src32 <= 12'hb91;
        src33 <= 12'hef0;
        src34 <= 12'h45a;
        src35 <= 12'h38;
        src36 <= 12'h253;
        src37 <= 12'hfdd;
        src38 <= 12'hb02;
        src39 <= 12'hed5;
        src40 <= 12'hdb6;
        src41 <= 12'h6d6;
        src42 <= 12'h8da;
        src43 <= 12'hb16;
        src44 <= 12'h530;
        src45 <= 12'h6df;
        src46 <= 12'hb0a;
        src47 <= 12'h7e1;
        src48 <= 12'h1f3;
        src49 <= 12'h8b3;
        src50 <= 12'hfb2;
        src51 <= 12'h9b0;
        src52 <= 12'h401;
        src53 <= 12'ha17;
        src54 <= 12'ha8a;
        src55 <= 12'ha23;
        src56 <= 12'hb5b;
        src57 <= 12'h7a0;
        src58 <= 12'h9e3;
        src59 <= 12'hebc;
        src60 <= 12'h51b;
        src61 <= 12'h1b8;
        src62 <= 12'h11;
        src63 <= 12'h9ab;
        src64 <= 12'h957;
        src65 <= 12'h6df;
        src66 <= 12'h9d8;
        src67 <= 12'h1a6;
        src68 <= 12'ha38;
        src69 <= 12'h3a5;
        src70 <= 12'h69e;
        src71 <= 12'hc69;
        src72 <= 12'hbfd;
        src73 <= 12'hf0f;
        src74 <= 12'hec9;
        src75 <= 12'h68c;
        src76 <= 12'h3e0;
        src77 <= 12'h755;
        src78 <= 12'h1af;
        src79 <= 12'h8be;
        src80 <= 12'hbfc;
        src81 <= 12'h68;
        src82 <= 12'hd41;
        src83 <= 12'hb9b;
        src84 <= 12'h5aa;
        src85 <= 12'h5a8;
        src86 <= 12'h19b;
        src87 <= 12'h53;
        src88 <= 12'h4bb;
        src89 <= 12'h343;
        src90 <= 12'ha97;
        src91 <= 12'haae;
        src92 <= 12'h7fd;
        src93 <= 12'hf09;
        src94 <= 12'he4b;
        src95 <= 12'haae;
        src96 <= 12'h3e7;
        src97 <= 12'h1ae;
        src98 <= 12'h1ce;
        src99 <= 12'hbb0;
        src100 <= 12'h79c;
        src101 <= 12'h5d2;
        src102 <= 12'h909;
        src103 <= 12'hcb5;
        src104 <= 12'hd0e;
        src105 <= 12'h12a;
        src106 <= 12'hec1;
        src107 <= 12'h356;
        src108 <= 12'h2;
        src109 <= 12'h432;
        src110 <= 12'h649;
        src111 <= 12'h3d7;
        src112 <= 12'h166;
        src113 <= 12'h2c9;
        src114 <= 12'h110;
        src115 <= 12'h8f2;
        src116 <= 12'h39b;
        src117 <= 12'hf39;
        src118 <= 12'h44e;
        src119 <= 12'hfaf;
        src120 <= 12'h1cd;
        src121 <= 12'hff2;
        src122 <= 12'hc0f;
        src123 <= 12'h238;
        src124 <= 12'hb74;
        src125 <= 12'h439;
        src126 <= 12'he5f;
        src127 <= 12'h8d2;
        src128 <= 12'hb06;
        src129 <= 12'hfa6;
        src130 <= 12'hfdc;
        src131 <= 12'h2ac;
        src132 <= 12'h590;
        src133 <= 12'h9f3;
        src134 <= 12'h960;
        src135 <= 12'hf30;
        src136 <= 12'hd23;
        src137 <= 12'h904;
        src138 <= 12'h29;
        src139 <= 12'h24f;
        src140 <= 12'h622;
        src141 <= 12'h470;
        src142 <= 12'h5fc;
        src143 <= 12'h9fd;
        src144 <= 12'hf15;
        src145 <= 12'h9cd;
        src146 <= 12'h922;
        src147 <= 12'h6a3;
        src148 <= 12'h8c;
        src149 <= 12'hf27;
        src150 <= 12'h34;
        src151 <= 12'ha17;
        src152 <= 12'h6ed;
        src153 <= 12'hda1;
        src154 <= 12'hd98;
        src155 <= 12'h71d;
        src156 <= 12'h1d0;
        src157 <= 12'h771;
        src158 <= 12'h585;
        src159 <= 12'h739;
        src160 <= 12'he46;
        src161 <= 12'hbe2;
        src162 <= 12'h533;
        src163 <= 12'hd58;
        src164 <= 12'hef6;
        src165 <= 12'h17f;
        src166 <= 12'h120;
        src167 <= 12'hd8e;
        src168 <= 12'h671;
        src169 <= 12'h809;
        src170 <= 12'h5b4;
        src171 <= 12'h8f;
        src172 <= 12'hab9;
        src173 <= 12'h3e7;
        src174 <= 12'h859;
        src175 <= 12'h7e;
        src176 <= 12'hcf2;
        src177 <= 12'hd3c;
        src178 <= 12'h5ce;
        src179 <= 12'hc8b;
        src180 <= 12'h3b6;
        src181 <= 12'h1f4;
        src182 <= 12'hc39;
        src183 <= 12'h442;
        src184 <= 12'h674;
        src185 <= 12'hc76;
        src186 <= 12'hed9;
        src187 <= 12'h5e7;
        src188 <= 12'hcf4;
        exp <= 20'h6059e;
        #1
        src0 <= 12'h980;
        src1 <= 12'hedd;
        src2 <= 12'hca2;
        src3 <= 12'h7a5;
        src4 <= 12'h8c2;
        src5 <= 12'h18b;
        src6 <= 12'h7e8;
        src7 <= 12'h852;
        src8 <= 12'hcb7;
        src9 <= 12'h50f;
        src10 <= 12'h9a8;
        src11 <= 12'h899;
        src12 <= 12'hd68;
        src13 <= 12'h44d;
        src14 <= 12'h46d;
        src15 <= 12'h92b;
        src16 <= 12'hc51;
        src17 <= 12'hb55;
        src18 <= 12'h307;
        src19 <= 12'h718;
        src20 <= 12'he3d;
        src21 <= 12'h918;
        src22 <= 12'he66;
        src23 <= 12'hb31;
        src24 <= 12'h5f5;
        src25 <= 12'h6d5;
        src26 <= 12'hb45;
        src27 <= 12'he32;
        src28 <= 12'h89;
        src29 <= 12'ha73;
        src30 <= 12'h76b;
        src31 <= 12'hd47;
        src32 <= 12'hd1f;
        src33 <= 12'h3d0;
        src34 <= 12'he8d;
        src35 <= 12'h5f9;
        src36 <= 12'h3de;
        src37 <= 12'hb34;
        src38 <= 12'h8e6;
        src39 <= 12'he8d;
        src40 <= 12'h956;
        src41 <= 12'h169;
        src42 <= 12'hf87;
        src43 <= 12'hc65;
        src44 <= 12'h3b7;
        src45 <= 12'h964;
        src46 <= 12'h94d;
        src47 <= 12'hb33;
        src48 <= 12'hc5f;
        src49 <= 12'h804;
        src50 <= 12'h83a;
        src51 <= 12'h5c6;
        src52 <= 12'h1a3;
        src53 <= 12'hac2;
        src54 <= 12'hfb7;
        src55 <= 12'h75d;
        src56 <= 12'h40e;
        src57 <= 12'h8f4;
        src58 <= 12'hf1c;
        src59 <= 12'h3e2;
        src60 <= 12'h468;
        src61 <= 12'h12e;
        src62 <= 12'h47a;
        src63 <= 12'h9;
        src64 <= 12'h9ca;
        src65 <= 12'h6dd;
        src66 <= 12'hd0c;
        src67 <= 12'had0;
        src68 <= 12'hc51;
        src69 <= 12'h922;
        src70 <= 12'h556;
        src71 <= 12'he90;
        src72 <= 12'h8ce;
        src73 <= 12'ha9a;
        src74 <= 12'ha40;
        src75 <= 12'h272;
        src76 <= 12'he5;
        src77 <= 12'h156;
        src78 <= 12'h875;
        src79 <= 12'h336;
        src80 <= 12'h945;
        src81 <= 12'h8ce;
        src82 <= 12'h86c;
        src83 <= 12'h9ab;
        src84 <= 12'hd92;
        src85 <= 12'hf49;
        src86 <= 12'h33a;
        src87 <= 12'h33a;
        src88 <= 12'h8df;
        src89 <= 12'ha83;
        src90 <= 12'he30;
        src91 <= 12'h580;
        src92 <= 12'hda9;
        src93 <= 12'h46a;
        src94 <= 12'h442;
        src95 <= 12'h5a7;
        src96 <= 12'hebe;
        src97 <= 12'hf86;
        src98 <= 12'hfce;
        src99 <= 12'h7f5;
        src100 <= 12'h2ee;
        src101 <= 12'hf8b;
        src102 <= 12'he64;
        src103 <= 12'h7f6;
        src104 <= 12'h463;
        src105 <= 12'hb93;
        src106 <= 12'hcb0;
        src107 <= 12'h53e;
        src108 <= 12'hac0;
        src109 <= 12'h6e;
        src110 <= 12'hfe3;
        src111 <= 12'h13f;
        src112 <= 12'h2d3;
        src113 <= 12'h6c3;
        src114 <= 12'hbf;
        src115 <= 12'hb72;
        src116 <= 12'h943;
        src117 <= 12'h4ad;
        src118 <= 12'h148;
        src119 <= 12'h642;
        src120 <= 12'h98c;
        src121 <= 12'h369;
        src122 <= 12'hc38;
        src123 <= 12'he3;
        src124 <= 12'h6bd;
        src125 <= 12'he7;
        src126 <= 12'h423;
        src127 <= 12'h2f5;
        src128 <= 12'h94e;
        src129 <= 12'h57f;
        src130 <= 12'hde6;
        src131 <= 12'h241;
        src132 <= 12'h4c3;
        src133 <= 12'ha14;
        src134 <= 12'hbf4;
        src135 <= 12'hd6a;
        src136 <= 12'h192;
        src137 <= 12'h474;
        src138 <= 12'hb05;
        src139 <= 12'h118;
        src140 <= 12'h4cc;
        src141 <= 12'h476;
        src142 <= 12'h59c;
        src143 <= 12'h7c0;
        src144 <= 12'h369;
        src145 <= 12'hb06;
        src146 <= 12'h910;
        src147 <= 12'hc4c;
        src148 <= 12'h2e9;
        src149 <= 12'h139;
        src150 <= 12'hd2;
        src151 <= 12'h5;
        src152 <= 12'h2ce;
        src153 <= 12'hbbb;
        src154 <= 12'he80;
        src155 <= 12'h949;
        src156 <= 12'h39e;
        src157 <= 12'h7e6;
        src158 <= 12'ha39;
        src159 <= 12'h261;
        src160 <= 12'hf44;
        src161 <= 12'h16b;
        src162 <= 12'he18;
        src163 <= 12'h93;
        src164 <= 12'hd21;
        src165 <= 12'h45e;
        src166 <= 12'h7ff;
        src167 <= 12'hf5c;
        src168 <= 12'hda2;
        src169 <= 12'h67a;
        src170 <= 12'h649;
        src171 <= 12'hb50;
        src172 <= 12'hd63;
        src173 <= 12'hc6e;
        src174 <= 12'h893;
        src175 <= 12'hd01;
        src176 <= 12'h124;
        src177 <= 12'hf99;
        src178 <= 12'h4ad;
        src179 <= 12'he1d;
        src180 <= 12'hcf1;
        src181 <= 12'h764;
        src182 <= 12'hcc8;
        src183 <= 12'hc0e;
        src184 <= 12'h1a9;
        src185 <= 12'h781;
        src186 <= 12'h329;
        src187 <= 12'hc8a;
        src188 <= 12'h46;
        exp <= 20'h60113;
        #1
        src0 <= 12'he85;
        src1 <= 12'h65e;
        src2 <= 12'hd1d;
        src3 <= 12'ha6a;
        src4 <= 12'h535;
        src5 <= 12'hcb2;
        src6 <= 12'h732;
        src7 <= 12'ha2a;
        src8 <= 12'hd55;
        src9 <= 12'hfc3;
        src10 <= 12'hd2b;
        src11 <= 12'hdde;
        src12 <= 12'h78f;
        src13 <= 12'h69d;
        src14 <= 12'h724;
        src15 <= 12'h22;
        src16 <= 12'h83b;
        src17 <= 12'h83a;
        src18 <= 12'h453;
        src19 <= 12'h65d;
        src20 <= 12'h16a;
        src21 <= 12'h4e6;
        src22 <= 12'hb47;
        src23 <= 12'h299;
        src24 <= 12'hb99;
        src25 <= 12'hae4;
        src26 <= 12'h157;
        src27 <= 12'hebc;
        src28 <= 12'h171;
        src29 <= 12'h89d;
        src30 <= 12'h7ad;
        src31 <= 12'h685;
        src32 <= 12'h67b;
        src33 <= 12'hf61;
        src34 <= 12'h3cf;
        src35 <= 12'he32;
        src36 <= 12'hb3;
        src37 <= 12'h53;
        src38 <= 12'h99c;
        src39 <= 12'ha27;
        src40 <= 12'hd9e;
        src41 <= 12'h8bd;
        src42 <= 12'h3d7;
        src43 <= 12'hc6d;
        src44 <= 12'h3cf;
        src45 <= 12'h165;
        src46 <= 12'hef6;
        src47 <= 12'hefa;
        src48 <= 12'hfbf;
        src49 <= 12'h9c2;
        src50 <= 12'h3d6;
        src51 <= 12'h615;
        src52 <= 12'h819;
        src53 <= 12'h157;
        src54 <= 12'h600;
        src55 <= 12'h493;
        src56 <= 12'hd13;
        src57 <= 12'h555;
        src58 <= 12'h8c0;
        src59 <= 12'h313;
        src60 <= 12'h88d;
        src61 <= 12'h31f;
        src62 <= 12'h242;
        src63 <= 12'hac9;
        src64 <= 12'had;
        src65 <= 12'h50b;
        src66 <= 12'ha88;
        src67 <= 12'hb78;
        src68 <= 12'hcd4;
        src69 <= 12'h8ba;
        src70 <= 12'hce5;
        src71 <= 12'h85f;
        src72 <= 12'he42;
        src73 <= 12'hb5c;
        src74 <= 12'hd4b;
        src75 <= 12'h496;
        src76 <= 12'he03;
        src77 <= 12'hdb4;
        src78 <= 12'h12e;
        src79 <= 12'hd0d;
        src80 <= 12'hc3e;
        src81 <= 12'h5b4;
        src82 <= 12'h9ed;
        src83 <= 12'hf21;
        src84 <= 12'hfbf;
        src85 <= 12'hc19;
        src86 <= 12'h5e;
        src87 <= 12'hfc9;
        src88 <= 12'hc9;
        src89 <= 12'hd6b;
        src90 <= 12'h5c2;
        src91 <= 12'h64f;
        src92 <= 12'h768;
        src93 <= 12'h743;
        src94 <= 12'hea9;
        src95 <= 12'h23f;
        src96 <= 12'hebd;
        src97 <= 12'hdc8;
        src98 <= 12'hafe;
        src99 <= 12'hb42;
        src100 <= 12'hbc3;
        src101 <= 12'hd36;
        src102 <= 12'hbc;
        src103 <= 12'hb0;
        src104 <= 12'he24;
        src105 <= 12'heec;
        src106 <= 12'hb90;
        src107 <= 12'h211;
        src108 <= 12'hab;
        src109 <= 12'hea1;
        src110 <= 12'ha10;
        src111 <= 12'hc89;
        src112 <= 12'hd2b;
        src113 <= 12'ha1d;
        src114 <= 12'h5b7;
        src115 <= 12'h94d;
        src116 <= 12'h3c5;
        src117 <= 12'h46e;
        src118 <= 12'h2c0;
        src119 <= 12'hb9;
        src120 <= 12'hd42;
        src121 <= 12'hd9c;
        src122 <= 12'h3;
        src123 <= 12'h505;
        src124 <= 12'h1b1;
        src125 <= 12'hb40;
        src126 <= 12'h26;
        src127 <= 12'h6d0;
        src128 <= 12'h82a;
        src129 <= 12'heb0;
        src130 <= 12'h204;
        src131 <= 12'hc0a;
        src132 <= 12'hb51;
        src133 <= 12'h421;
        src134 <= 12'h560;
        src135 <= 12'h9eb;
        src136 <= 12'he3f;
        src137 <= 12'h49d;
        src138 <= 12'hf7e;
        src139 <= 12'hd90;
        src140 <= 12'h379;
        src141 <= 12'h3f;
        src142 <= 12'hec9;
        src143 <= 12'h6f8;
        src144 <= 12'hb47;
        src145 <= 12'h960;
        src146 <= 12'hbef;
        src147 <= 12'he9b;
        src148 <= 12'h271;
        src149 <= 12'he57;
        src150 <= 12'hf02;
        src151 <= 12'ha7a;
        src152 <= 12'haf2;
        src153 <= 12'h242;
        src154 <= 12'hb23;
        src155 <= 12'h5c0;
        src156 <= 12'h3f4;
        src157 <= 12'ha7d;
        src158 <= 12'h6dc;
        src159 <= 12'h4a;
        src160 <= 12'ha12;
        src161 <= 12'h12d;
        src162 <= 12'ha35;
        src163 <= 12'h6b0;
        src164 <= 12'h13f;
        src165 <= 12'hc88;
        src166 <= 12'h474;
        src167 <= 12'hb45;
        src168 <= 12'h6a6;
        src169 <= 12'hbfd;
        src170 <= 12'h5b6;
        src171 <= 12'h86b;
        src172 <= 12'h1e5;
        src173 <= 12'h88a;
        src174 <= 12'h9f9;
        src175 <= 12'hca1;
        src176 <= 12'h1c3;
        src177 <= 12'heae;
        src178 <= 12'h4ee;
        src179 <= 12'h2ce;
        src180 <= 12'h938;
        src181 <= 12'h5d1;
        src182 <= 12'h71;
        src183 <= 12'hb3;
        src184 <= 12'hf00;
        src185 <= 12'h1a7;
        src186 <= 12'hf9a;
        src187 <= 12'hc0d;
        src188 <= 12'h73b;
        exp <= 20'h62205;
        #1
        src0 <= 12'h133;
        src1 <= 12'hd30;
        src2 <= 12'ha9c;
        src3 <= 12'hd17;
        src4 <= 12'hee7;
        src5 <= 12'h402;
        src6 <= 12'he18;
        src7 <= 12'hdba;
        src8 <= 12'h765;
        src9 <= 12'h71e;
        src10 <= 12'hd8f;
        src11 <= 12'h241;
        src12 <= 12'hef6;
        src13 <= 12'h44f;
        src14 <= 12'h62e;
        src15 <= 12'hfef;
        src16 <= 12'hc6f;
        src17 <= 12'h9d7;
        src18 <= 12'h4fe;
        src19 <= 12'hed0;
        src20 <= 12'h420;
        src21 <= 12'h7c;
        src22 <= 12'hbb3;
        src23 <= 12'h93a;
        src24 <= 12'he78;
        src25 <= 12'h12;
        src26 <= 12'hbc0;
        src27 <= 12'haa7;
        src28 <= 12'hfab;
        src29 <= 12'hdfb;
        src30 <= 12'h5c9;
        src31 <= 12'hd78;
        src32 <= 12'h760;
        src33 <= 12'hdcb;
        src34 <= 12'h2ed;
        src35 <= 12'hf62;
        src36 <= 12'h31e;
        src37 <= 12'hb39;
        src38 <= 12'h3e2;
        src39 <= 12'h787;
        src40 <= 12'haf2;
        src41 <= 12'h705;
        src42 <= 12'hccb;
        src43 <= 12'hc33;
        src44 <= 12'h447;
        src45 <= 12'h38d;
        src46 <= 12'h183;
        src47 <= 12'h7a5;
        src48 <= 12'h90a;
        src49 <= 12'h107;
        src50 <= 12'h5d5;
        src51 <= 12'h5b0;
        src52 <= 12'hfda;
        src53 <= 12'hd81;
        src54 <= 12'h10e;
        src55 <= 12'h97f;
        src56 <= 12'h2de;
        src57 <= 12'h60d;
        src58 <= 12'h4af;
        src59 <= 12'h243;
        src60 <= 12'hb0e;
        src61 <= 12'h316;
        src62 <= 12'hbcf;
        src63 <= 12'hbc8;
        src64 <= 12'h668;
        src65 <= 12'hf6;
        src66 <= 12'he92;
        src67 <= 12'h134;
        src68 <= 12'hd70;
        src69 <= 12'h4a7;
        src70 <= 12'h129;
        src71 <= 12'h568;
        src72 <= 12'he6f;
        src73 <= 12'hf02;
        src74 <= 12'hb4;
        src75 <= 12'hfd9;
        src76 <= 12'h914;
        src77 <= 12'ha0a;
        src78 <= 12'h4a4;
        src79 <= 12'h892;
        src80 <= 12'h747;
        src81 <= 12'hfc2;
        src82 <= 12'hba5;
        src83 <= 12'h9b6;
        src84 <= 12'h4b0;
        src85 <= 12'h457;
        src86 <= 12'h617;
        src87 <= 12'h609;
        src88 <= 12'hc95;
        src89 <= 12'hcd3;
        src90 <= 12'h174;
        src91 <= 12'h596;
        src92 <= 12'h545;
        src93 <= 12'h3f8;
        src94 <= 12'h91;
        src95 <= 12'hf52;
        src96 <= 12'ha19;
        src97 <= 12'h7b4;
        src98 <= 12'hca;
        src99 <= 12'hfcb;
        src100 <= 12'h891;
        src101 <= 12'h534;
        src102 <= 12'hf6b;
        src103 <= 12'h375;
        src104 <= 12'h961;
        src105 <= 12'h8cc;
        src106 <= 12'he04;
        src107 <= 12'hc57;
        src108 <= 12'h911;
        src109 <= 12'h50f;
        src110 <= 12'hd6e;
        src111 <= 12'h71a;
        src112 <= 12'h420;
        src113 <= 12'hb6d;
        src114 <= 12'hd71;
        src115 <= 12'h6df;
        src116 <= 12'h190;
        src117 <= 12'h22d;
        src118 <= 12'h669;
        src119 <= 12'h710;
        src120 <= 12'h207;
        src121 <= 12'h265;
        src122 <= 12'h462;
        src123 <= 12'hd83;
        src124 <= 12'he7c;
        src125 <= 12'h94f;
        src126 <= 12'h7bc;
        src127 <= 12'h9a0;
        src128 <= 12'hec4;
        src129 <= 12'hf91;
        src130 <= 12'h366;
        src131 <= 12'hb08;
        src132 <= 12'hfc;
        src133 <= 12'h73d;
        src134 <= 12'h142;
        src135 <= 12'h24b;
        src136 <= 12'h3e9;
        src137 <= 12'h55f;
        src138 <= 12'he08;
        src139 <= 12'hc97;
        src140 <= 12'h6e0;
        src141 <= 12'h837;
        src142 <= 12'h92a;
        src143 <= 12'h762;
        src144 <= 12'h590;
        src145 <= 12'h67d;
        src146 <= 12'h934;
        src147 <= 12'h801;
        src148 <= 12'h924;
        src149 <= 12'h9ee;
        src150 <= 12'h522;
        src151 <= 12'h227;
        src152 <= 12'h7d3;
        src153 <= 12'h9d3;
        src154 <= 12'h25b;
        src155 <= 12'hab1;
        src156 <= 12'hf8f;
        src157 <= 12'hcd4;
        src158 <= 12'h3c3;
        src159 <= 12'h159;
        src160 <= 12'h33;
        src161 <= 12'h7ca;
        src162 <= 12'ha8f;
        src163 <= 12'h778;
        src164 <= 12'h802;
        src165 <= 12'hb2d;
        src166 <= 12'hc19;
        src167 <= 12'hb49;
        src168 <= 12'h251;
        src169 <= 12'h413;
        src170 <= 12'hc2e;
        src171 <= 12'h461;
        src172 <= 12'h28;
        src173 <= 12'hb1b;
        src174 <= 12'hd58;
        src175 <= 12'hafa;
        src176 <= 12'h7cc;
        src177 <= 12'he46;
        src178 <= 12'h923;
        src179 <= 12'h9bf;
        src180 <= 12'h53f;
        src181 <= 12'hd34;
        src182 <= 12'h6f9;
        src183 <= 12'h9f2;
        src184 <= 12'h86e;
        src185 <= 12'h236;
        src186 <= 12'hfa3;
        src187 <= 12'hda3;
        src188 <= 12'hcb1;
        exp <= 20'h61a24;
        #1
        src0 <= 12'h7c3;
        src1 <= 12'h56;
        src2 <= 12'h1f2;
        src3 <= 12'hbcc;
        src4 <= 12'hfc7;
        src5 <= 12'hd3e;
        src6 <= 12'hed2;
        src7 <= 12'h879;
        src8 <= 12'h91e;
        src9 <= 12'h39b;
        src10 <= 12'hd96;
        src11 <= 12'h92d;
        src12 <= 12'hb09;
        src13 <= 12'he6a;
        src14 <= 12'h6ff;
        src15 <= 12'hab7;
        src16 <= 12'h1dc;
        src17 <= 12'h461;
        src18 <= 12'h309;
        src19 <= 12'h60f;
        src20 <= 12'h6a2;
        src21 <= 12'hd49;
        src22 <= 12'h424;
        src23 <= 12'hce7;
        src24 <= 12'h270;
        src25 <= 12'had3;
        src26 <= 12'h842;
        src27 <= 12'h4e;
        src28 <= 12'h3e0;
        src29 <= 12'h224;
        src30 <= 12'he1a;
        src31 <= 12'hf62;
        src32 <= 12'ha4b;
        src33 <= 12'hf10;
        src34 <= 12'h4a;
        src35 <= 12'h3b7;
        src36 <= 12'h6b7;
        src37 <= 12'h5d;
        src38 <= 12'h3f8;
        src39 <= 12'he92;
        src40 <= 12'h6b5;
        src41 <= 12'hdc3;
        src42 <= 12'h453;
        src43 <= 12'h767;
        src44 <= 12'h943;
        src45 <= 12'h9c;
        src46 <= 12'h93f;
        src47 <= 12'h65a;
        src48 <= 12'hbf4;
        src49 <= 12'h4b6;
        src50 <= 12'h58e;
        src51 <= 12'h620;
        src52 <= 12'h764;
        src53 <= 12'he05;
        src54 <= 12'hcff;
        src55 <= 12'hd1d;
        src56 <= 12'h9a4;
        src57 <= 12'hc3e;
        src58 <= 12'hd96;
        src59 <= 12'h4d6;
        src60 <= 12'h2fe;
        src61 <= 12'hba8;
        src62 <= 12'h8e5;
        src63 <= 12'h528;
        src64 <= 12'h5bd;
        src65 <= 12'hd23;
        src66 <= 12'h9e2;
        src67 <= 12'h904;
        src68 <= 12'hc3f;
        src69 <= 12'h59b;
        src70 <= 12'he7a;
        src71 <= 12'h2ec;
        src72 <= 12'h6b2;
        src73 <= 12'h210;
        src74 <= 12'h59f;
        src75 <= 12'h44d;
        src76 <= 12'hdf3;
        src77 <= 12'hb6b;
        src78 <= 12'h458;
        src79 <= 12'h22b;
        src80 <= 12'h509;
        src81 <= 12'hedc;
        src82 <= 12'h7a;
        src83 <= 12'hbaa;
        src84 <= 12'hce6;
        src85 <= 12'ha4a;
        src86 <= 12'h763;
        src87 <= 12'he4d;
        src88 <= 12'h160;
        src89 <= 12'ha57;
        src90 <= 12'h95;
        src91 <= 12'he7a;
        src92 <= 12'he1b;
        src93 <= 12'h30d;
        src94 <= 12'hcb0;
        src95 <= 12'h88f;
        src96 <= 12'h69d;
        src97 <= 12'hf42;
        src98 <= 12'h537;
        src99 <= 12'h5ff;
        src100 <= 12'h604;
        src101 <= 12'h815;
        src102 <= 12'h6d5;
        src103 <= 12'h841;
        src104 <= 12'h114;
        src105 <= 12'haa0;
        src106 <= 12'h588;
        src107 <= 12'h7e1;
        src108 <= 12'h1db;
        src109 <= 12'hada;
        src110 <= 12'h7;
        src111 <= 12'hac8;
        src112 <= 12'h20;
        src113 <= 12'h793;
        src114 <= 12'h2c4;
        src115 <= 12'h13a;
        src116 <= 12'h2ea;
        src117 <= 12'h482;
        src118 <= 12'h4e0;
        src119 <= 12'heaa;
        src120 <= 12'hee5;
        src121 <= 12'h937;
        src122 <= 12'h2ba;
        src123 <= 12'ha5e;
        src124 <= 12'h24c;
        src125 <= 12'he4e;
        src126 <= 12'h580;
        src127 <= 12'h4c1;
        src128 <= 12'h751;
        src129 <= 12'hd81;
        src130 <= 12'h9c6;
        src131 <= 12'hb2e;
        src132 <= 12'h2d4;
        src133 <= 12'hcde;
        src134 <= 12'h3e4;
        src135 <= 12'h9e9;
        src136 <= 12'hb6b;
        src137 <= 12'he1c;
        src138 <= 12'h92a;
        src139 <= 12'h801;
        src140 <= 12'h6b8;
        src141 <= 12'h11a;
        src142 <= 12'h8ef;
        src143 <= 12'he6;
        src144 <= 12'h573;
        src145 <= 12'h30e;
        src146 <= 12'h719;
        src147 <= 12'hddc;
        src148 <= 12'h4ef;
        src149 <= 12'hefb;
        src150 <= 12'h668;
        src151 <= 12'hb0;
        src152 <= 12'h594;
        src153 <= 12'hed;
        src154 <= 12'h563;
        src155 <= 12'h730;
        src156 <= 12'h742;
        src157 <= 12'h276;
        src158 <= 12'h29;
        src159 <= 12'hfd9;
        src160 <= 12'hcd1;
        src161 <= 12'h7b;
        src162 <= 12'hc2c;
        src163 <= 12'hc62;
        src164 <= 12'h48d;
        src165 <= 12'hbf1;
        src166 <= 12'h7a8;
        src167 <= 12'h73e;
        src168 <= 12'heac;
        src169 <= 12'hc10;
        src170 <= 12'ha67;
        src171 <= 12'h378;
        src172 <= 12'h64a;
        src173 <= 12'h52f;
        src174 <= 12'hc17;
        src175 <= 12'hff5;
        src176 <= 12'hfc6;
        src177 <= 12'hb58;
        src178 <= 12'h539;
        src179 <= 12'h798;
        src180 <= 12'ha4;
        src181 <= 12'h5ad;
        src182 <= 12'hdf4;
        src183 <= 12'h181;
        src184 <= 12'hbd9;
        src185 <= 12'h243;
        src186 <= 12'h62f;
        src187 <= 12'h673;
        src188 <= 12'h962;
        exp <= 20'h5c749;
        #1
        src0 <= 12'hc05;
        src1 <= 12'h752;
        src2 <= 12'he11;
        src3 <= 12'hb97;
        src4 <= 12'h3c2;
        src5 <= 12'h2c7;
        src6 <= 12'he8f;
        src7 <= 12'h4af;
        src8 <= 12'h743;
        src9 <= 12'hcf0;
        src10 <= 12'h780;
        src11 <= 12'hd5f;
        src12 <= 12'h497;
        src13 <= 12'hf90;
        src14 <= 12'h1ab;
        src15 <= 12'h98c;
        src16 <= 12'h1e4;
        src17 <= 12'h1d9;
        src18 <= 12'hb20;
        src19 <= 12'hef;
        src20 <= 12'h2b8;
        src21 <= 12'hfb0;
        src22 <= 12'h877;
        src23 <= 12'h295;
        src24 <= 12'ha18;
        src25 <= 12'h9de;
        src26 <= 12'h7ec;
        src27 <= 12'h407;
        src28 <= 12'h1ab;
        src29 <= 12'h88f;
        src30 <= 12'hdc9;
        src31 <= 12'h772;
        src32 <= 12'h8e3;
        src33 <= 12'he4a;
        src34 <= 12'h217;
        src35 <= 12'h2f0;
        src36 <= 12'h373;
        src37 <= 12'h3e4;
        src38 <= 12'h10b;
        src39 <= 12'hca9;
        src40 <= 12'h402;
        src41 <= 12'h232;
        src42 <= 12'h885;
        src43 <= 12'hcc9;
        src44 <= 12'h711;
        src45 <= 12'h5a4;
        src46 <= 12'he11;
        src47 <= 12'hb17;
        src48 <= 12'h65c;
        src49 <= 12'h8e4;
        src50 <= 12'h6f6;
        src51 <= 12'h40f;
        src52 <= 12'h3da;
        src53 <= 12'h32b;
        src54 <= 12'hd09;
        src55 <= 12'h36c;
        src56 <= 12'h660;
        src57 <= 12'h504;
        src58 <= 12'ha23;
        src59 <= 12'h8de;
        src60 <= 12'h4fa;
        src61 <= 12'h8ef;
        src62 <= 12'h669;
        src63 <= 12'h584;
        src64 <= 12'h245;
        src65 <= 12'hd1e;
        src66 <= 12'h99c;
        src67 <= 12'h7b;
        src68 <= 12'hb93;
        src69 <= 12'h10c;
        src70 <= 12'h366;
        src71 <= 12'hc91;
        src72 <= 12'h8fc;
        src73 <= 12'ha00;
        src74 <= 12'hada;
        src75 <= 12'h478;
        src76 <= 12'h7d7;
        src77 <= 12'h8c6;
        src78 <= 12'h370;
        src79 <= 12'h107;
        src80 <= 12'h1c1;
        src81 <= 12'h61e;
        src82 <= 12'hb84;
        src83 <= 12'hb96;
        src84 <= 12'h7ef;
        src85 <= 12'h866;
        src86 <= 12'ha46;
        src87 <= 12'hdf9;
        src88 <= 12'h12;
        src89 <= 12'hae1;
        src90 <= 12'h27e;
        src91 <= 12'h77d;
        src92 <= 12'h334;
        src93 <= 12'hc96;
        src94 <= 12'hcbe;
        src95 <= 12'h153;
        src96 <= 12'hffe;
        src97 <= 12'h5a;
        src98 <= 12'h4f4;
        src99 <= 12'h960;
        src100 <= 12'h16d;
        src101 <= 12'h15d;
        src102 <= 12'h489;
        src103 <= 12'he62;
        src104 <= 12'h742;
        src105 <= 12'he7e;
        src106 <= 12'he0f;
        src107 <= 12'hb86;
        src108 <= 12'h2a2;
        src109 <= 12'h280;
        src110 <= 12'h91d;
        src111 <= 12'h7f5;
        src112 <= 12'h66a;
        src113 <= 12'h944;
        src114 <= 12'h14b;
        src115 <= 12'h397;
        src116 <= 12'h8b2;
        src117 <= 12'h9e3;
        src118 <= 12'hc2d;
        src119 <= 12'h7c1;
        src120 <= 12'h4ea;
        src121 <= 12'hb2e;
        src122 <= 12'h570;
        src123 <= 12'h3b4;
        src124 <= 12'he3f;
        src125 <= 12'h53d;
        src126 <= 12'h7c;
        src127 <= 12'hae0;
        src128 <= 12'hae4;
        src129 <= 12'hbf7;
        src130 <= 12'ha71;
        src131 <= 12'ha0e;
        src132 <= 12'h312;
        src133 <= 12'h26e;
        src134 <= 12'h19a;
        src135 <= 12'ha2d;
        src136 <= 12'he6e;
        src137 <= 12'h678;
        src138 <= 12'h800;
        src139 <= 12'hf60;
        src140 <= 12'h331;
        src141 <= 12'h65c;
        src142 <= 12'h3a5;
        src143 <= 12'hae6;
        src144 <= 12'hc5e;
        src145 <= 12'h4a6;
        src146 <= 12'hf3c;
        src147 <= 12'h8b;
        src148 <= 12'h995;
        src149 <= 12'h886;
        src150 <= 12'h74;
        src151 <= 12'hfb8;
        src152 <= 12'hfb;
        src153 <= 12'h6a5;
        src154 <= 12'h937;
        src155 <= 12'h425;
        src156 <= 12'h45f;
        src157 <= 12'hfe2;
        src158 <= 12'hcd;
        src159 <= 12'h396;
        src160 <= 12'h12b;
        src161 <= 12'h505;
        src162 <= 12'h9f7;
        src163 <= 12'haa5;
        src164 <= 12'hb72;
        src165 <= 12'h4a9;
        src166 <= 12'ha35;
        src167 <= 12'h9ee;
        src168 <= 12'h316;
        src169 <= 12'h83e;
        src170 <= 12'h490;
        src171 <= 12'hdf0;
        src172 <= 12'h87a;
        src173 <= 12'h2e4;
        src174 <= 12'h4c1;
        src175 <= 12'h856;
        src176 <= 12'hb68;
        src177 <= 12'hf18;
        src178 <= 12'hdde;
        src179 <= 12'h868;
        src180 <= 12'h8fb;
        src181 <= 12'h289;
        src182 <= 12'hc3f;
        src183 <= 12'h8a7;
        src184 <= 12'had4;
        src185 <= 12'hf93;
        src186 <= 12'h166;
        src187 <= 12'h65b;
        src188 <= 12'h2b5;
        exp <= 20'h58a56;
        #1
        src0 <= 12'h7f8;
        src1 <= 12'hb59;
        src2 <= 12'h30c;
        src3 <= 12'h739;
        src4 <= 12'hc82;
        src5 <= 12'hcb9;
        src6 <= 12'heb9;
        src7 <= 12'h608;
        src8 <= 12'ha4f;
        src9 <= 12'hf99;
        src10 <= 12'h83d;
        src11 <= 12'h67f;
        src12 <= 12'h7c7;
        src13 <= 12'h8f1;
        src14 <= 12'hf8c;
        src15 <= 12'h507;
        src16 <= 12'hf15;
        src17 <= 12'h8f2;
        src18 <= 12'h1b9;
        src19 <= 12'h996;
        src20 <= 12'h262;
        src21 <= 12'hb77;
        src22 <= 12'hef7;
        src23 <= 12'h299;
        src24 <= 12'hae3;
        src25 <= 12'hb4d;
        src26 <= 12'h102;
        src27 <= 12'hf5f;
        src28 <= 12'h1b0;
        src29 <= 12'h924;
        src30 <= 12'hc08;
        src31 <= 12'h7dd;
        src32 <= 12'h5a3;
        src33 <= 12'h91b;
        src34 <= 12'h7fb;
        src35 <= 12'h94d;
        src36 <= 12'h742;
        src37 <= 12'hd0d;
        src38 <= 12'h9b8;
        src39 <= 12'hc52;
        src40 <= 12'h45d;
        src41 <= 12'hb3;
        src42 <= 12'ha8d;
        src43 <= 12'h277;
        src44 <= 12'h1f3;
        src45 <= 12'hc58;
        src46 <= 12'hc6d;
        src47 <= 12'h8e9;
        src48 <= 12'he5b;
        src49 <= 12'hbe7;
        src50 <= 12'h88b;
        src51 <= 12'h894;
        src52 <= 12'hd9f;
        src53 <= 12'h78e;
        src54 <= 12'h667;
        src55 <= 12'heab;
        src56 <= 12'h76d;
        src57 <= 12'h6f1;
        src58 <= 12'hbea;
        src59 <= 12'h8e;
        src60 <= 12'h185;
        src61 <= 12'h3cf;
        src62 <= 12'hd60;
        src63 <= 12'he4c;
        src64 <= 12'h34e;
        src65 <= 12'h38;
        src66 <= 12'hfa7;
        src67 <= 12'ha46;
        src68 <= 12'h1d2;
        src69 <= 12'h318;
        src70 <= 12'hd5b;
        src71 <= 12'h9cf;
        src72 <= 12'hd0f;
        src73 <= 12'ha23;
        src74 <= 12'hb7b;
        src75 <= 12'h58f;
        src76 <= 12'hdd4;
        src77 <= 12'h287;
        src78 <= 12'h229;
        src79 <= 12'hca3;
        src80 <= 12'hb13;
        src81 <= 12'h326;
        src82 <= 12'hd40;
        src83 <= 12'ha09;
        src84 <= 12'h496;
        src85 <= 12'h9b6;
        src86 <= 12'h125;
        src87 <= 12'h1dd;
        src88 <= 12'h65c;
        src89 <= 12'h6f6;
        src90 <= 12'h632;
        src91 <= 12'h901;
        src92 <= 12'hcfa;
        src93 <= 12'hd71;
        src94 <= 12'hff;
        src95 <= 12'hddb;
        src96 <= 12'h323;
        src97 <= 12'h42b;
        src98 <= 12'h220;
        src99 <= 12'h8c9;
        src100 <= 12'h295;
        src101 <= 12'h59c;
        src102 <= 12'h81e;
        src103 <= 12'h766;
        src104 <= 12'hd12;
        src105 <= 12'ha2e;
        src106 <= 12'hdeb;
        src107 <= 12'h884;
        src108 <= 12'hf18;
        src109 <= 12'h204;
        src110 <= 12'h6eb;
        src111 <= 12'hadd;
        src112 <= 12'h5ba;
        src113 <= 12'h753;
        src114 <= 12'h133;
        src115 <= 12'h2ec;
        src116 <= 12'h86c;
        src117 <= 12'hb6;
        src118 <= 12'h19c;
        src119 <= 12'h69a;
        src120 <= 12'h590;
        src121 <= 12'h6a6;
        src122 <= 12'hf43;
        src123 <= 12'h47b;
        src124 <= 12'h6b6;
        src125 <= 12'h115;
        src126 <= 12'h897;
        src127 <= 12'hd71;
        src128 <= 12'h71e;
        src129 <= 12'h672;
        src130 <= 12'h8da;
        src131 <= 12'h2e6;
        src132 <= 12'hbb1;
        src133 <= 12'hcf7;
        src134 <= 12'h743;
        src135 <= 12'h924;
        src136 <= 12'hc99;
        src137 <= 12'h42;
        src138 <= 12'h46f;
        src139 <= 12'h62c;
        src140 <= 12'hdf3;
        src141 <= 12'h442;
        src142 <= 12'h7fb;
        src143 <= 12'h19b;
        src144 <= 12'hf9d;
        src145 <= 12'h2b3;
        src146 <= 12'hc78;
        src147 <= 12'h42f;
        src148 <= 12'haed;
        src149 <= 12'hc85;
        src150 <= 12'h2e6;
        src151 <= 12'h5e1;
        src152 <= 12'hb47;
        src153 <= 12'hb4f;
        src154 <= 12'he45;
        src155 <= 12'h88a;
        src156 <= 12'h41b;
        src157 <= 12'h3d9;
        src158 <= 12'h1b5;
        src159 <= 12'h702;
        src160 <= 12'hf02;
        src161 <= 12'h7b5;
        src162 <= 12'h463;
        src163 <= 12'h5a1;
        src164 <= 12'hdc0;
        src165 <= 12'h564;
        src166 <= 12'hece;
        src167 <= 12'hc43;
        src168 <= 12'h221;
        src169 <= 12'hc30;
        src170 <= 12'h57c;
        src171 <= 12'h47;
        src172 <= 12'he67;
        src173 <= 12'h9bc;
        src174 <= 12'h116;
        src175 <= 12'hbb0;
        src176 <= 12'hef;
        src177 <= 12'hfcc;
        src178 <= 12'hc66;
        src179 <= 12'hc64;
        src180 <= 12'h797;
        src181 <= 12'h1d4;
        src182 <= 12'hb45;
        src183 <= 12'ha08;
        src184 <= 12'h51;
        src185 <= 12'h3c8;
        src186 <= 12'ha85;
        src187 <= 12'hfa7;
        src188 <= 12'h35a;
        exp <= 20'h5f40b;
        #1
        src0 <= 12'h71e;
        src1 <= 12'hcf2;
        src2 <= 12'h207;
        src3 <= 12'h74f;
        src4 <= 12'h775;
        src5 <= 12'h1a3;
        src6 <= 12'h3f5;
        src7 <= 12'he3f;
        src8 <= 12'hb00;
        src9 <= 12'hc8c;
        src10 <= 12'h144;
        src11 <= 12'hd52;
        src12 <= 12'h994;
        src13 <= 12'h4c3;
        src14 <= 12'hc8e;
        src15 <= 12'h900;
        src16 <= 12'h9e5;
        src17 <= 12'h945;
        src18 <= 12'hd03;
        src19 <= 12'hff3;
        src20 <= 12'h51;
        src21 <= 12'hef7;
        src22 <= 12'ha4;
        src23 <= 12'hc1e;
        src24 <= 12'ha44;
        src25 <= 12'h473;
        src26 <= 12'hef7;
        src27 <= 12'hdcd;
        src28 <= 12'hf89;
        src29 <= 12'hf04;
        src30 <= 12'h9bc;
        src31 <= 12'hf4b;
        src32 <= 12'h4b0;
        src33 <= 12'h63c;
        src34 <= 12'hd82;
        src35 <= 12'h8f4;
        src36 <= 12'h8ff;
        src37 <= 12'h2f8;
        src38 <= 12'h810;
        src39 <= 12'h46e;
        src40 <= 12'h435;
        src41 <= 12'h35a;
        src42 <= 12'ha50;
        src43 <= 12'hfa;
        src44 <= 12'hc58;
        src45 <= 12'hc41;
        src46 <= 12'hd9e;
        src47 <= 12'h5b2;
        src48 <= 12'h8e6;
        src49 <= 12'h506;
        src50 <= 12'h9bf;
        src51 <= 12'h6a;
        src52 <= 12'h282;
        src53 <= 12'h782;
        src54 <= 12'h955;
        src55 <= 12'hc03;
        src56 <= 12'h67d;
        src57 <= 12'h6cd;
        src58 <= 12'h4ea;
        src59 <= 12'hbb5;
        src60 <= 12'hf5a;
        src61 <= 12'hcbd;
        src62 <= 12'h133;
        src63 <= 12'h3d8;
        src64 <= 12'hcc9;
        src65 <= 12'habb;
        src66 <= 12'h5db;
        src67 <= 12'h7e;
        src68 <= 12'he20;
        src69 <= 12'hf68;
        src70 <= 12'hbb;
        src71 <= 12'h60e;
        src72 <= 12'hf6f;
        src73 <= 12'h55d;
        src74 <= 12'h36;
        src75 <= 12'ha9c;
        src76 <= 12'h3b3;
        src77 <= 12'h7a5;
        src78 <= 12'h26b;
        src79 <= 12'hbc0;
        src80 <= 12'h1a2;
        src81 <= 12'h97b;
        src82 <= 12'h9d;
        src83 <= 12'h8e0;
        src84 <= 12'h8c7;
        src85 <= 12'h31f;
        src86 <= 12'hf6;
        src87 <= 12'hb5e;
        src88 <= 12'h1b1;
        src89 <= 12'hada;
        src90 <= 12'hb09;
        src91 <= 12'h495;
        src92 <= 12'hdf7;
        src93 <= 12'h25e;
        src94 <= 12'h378;
        src95 <= 12'h1b0;
        src96 <= 12'ha7d;
        src97 <= 12'heb0;
        src98 <= 12'h7d1;
        src99 <= 12'h76;
        src100 <= 12'h9c5;
        src101 <= 12'hc7;
        src102 <= 12'h512;
        src103 <= 12'hec5;
        src104 <= 12'h383;
        src105 <= 12'hcfd;
        src106 <= 12'h1b1;
        src107 <= 12'hbbe;
        src108 <= 12'ha75;
        src109 <= 12'h32b;
        src110 <= 12'h105;
        src111 <= 12'h5e6;
        src112 <= 12'h2e6;
        src113 <= 12'h752;
        src114 <= 12'hef9;
        src115 <= 12'ha25;
        src116 <= 12'h3a6;
        src117 <= 12'h5c;
        src118 <= 12'h983;
        src119 <= 12'h396;
        src120 <= 12'hcc0;
        src121 <= 12'hc79;
        src122 <= 12'hb2b;
        src123 <= 12'hecc;
        src124 <= 12'h27b;
        src125 <= 12'h4d2;
        src126 <= 12'h8bb;
        src127 <= 12'hb17;
        src128 <= 12'hb29;
        src129 <= 12'habe;
        src130 <= 12'hc42;
        src131 <= 12'h67e;
        src132 <= 12'h748;
        src133 <= 12'hbe;
        src134 <= 12'habc;
        src135 <= 12'h873;
        src136 <= 12'h6d4;
        src137 <= 12'hbe1;
        src138 <= 12'hc22;
        src139 <= 12'he;
        src140 <= 12'h4fb;
        src141 <= 12'h52;
        src142 <= 12'hc2d;
        src143 <= 12'h879;
        src144 <= 12'h545;
        src145 <= 12'h4d1;
        src146 <= 12'h616;
        src147 <= 12'h852;
        src148 <= 12'h634;
        src149 <= 12'h2ed;
        src150 <= 12'hcad;
        src151 <= 12'he30;
        src152 <= 12'h2b2;
        src153 <= 12'h4be;
        src154 <= 12'hc17;
        src155 <= 12'hb1;
        src156 <= 12'h760;
        src157 <= 12'ha9;
        src158 <= 12'ha3;
        src159 <= 12'h825;
        src160 <= 12'h185;
        src161 <= 12'had6;
        src162 <= 12'h2eb;
        src163 <= 12'hd50;
        src164 <= 12'ha74;
        src165 <= 12'hc00;
        src166 <= 12'h13e;
        src167 <= 12'hf04;
        src168 <= 12'h8f5;
        src169 <= 12'h5a3;
        src170 <= 12'hb5;
        src171 <= 12'h591;
        src172 <= 12'h350;
        src173 <= 12'h406;
        src174 <= 12'hce3;
        src175 <= 12'h8a7;
        src176 <= 12'hf8b;
        src177 <= 12'h759;
        src178 <= 12'hf6f;
        src179 <= 12'hd64;
        src180 <= 12'he90;
        src181 <= 12'h32b;
        src182 <= 12'h96b;
        src183 <= 12'h8d0;
        src184 <= 12'h3da;
        src185 <= 12'hb53;
        src186 <= 12'hca2;
        src187 <= 12'hd17;
        src188 <= 12'h2f1;
        exp <= 20'h5c6a8;
        #1
        src0 <= 12'h612;
        src1 <= 12'h3e7;
        src2 <= 12'h758;
        src3 <= 12'hdb1;
        src4 <= 12'h9bc;
        src5 <= 12'hdd4;
        src6 <= 12'h200;
        src7 <= 12'h59f;
        src8 <= 12'heea;
        src9 <= 12'h30d;
        src10 <= 12'hcf6;
        src11 <= 12'h69;
        src12 <= 12'ha02;
        src13 <= 12'h433;
        src14 <= 12'h3d0;
        src15 <= 12'h1e1;
        src16 <= 12'haf9;
        src17 <= 12'h2c;
        src18 <= 12'hbca;
        src19 <= 12'h682;
        src20 <= 12'h9b9;
        src21 <= 12'h477;
        src22 <= 12'hcdb;
        src23 <= 12'h4fc;
        src24 <= 12'hd0b;
        src25 <= 12'h573;
        src26 <= 12'hda3;
        src27 <= 12'h36f;
        src28 <= 12'h79;
        src29 <= 12'h309;
        src30 <= 12'hea9;
        src31 <= 12'ha6e;
        src32 <= 12'hb83;
        src33 <= 12'h201;
        src34 <= 12'h526;
        src35 <= 12'h846;
        src36 <= 12'h4da;
        src37 <= 12'ha02;
        src38 <= 12'haec;
        src39 <= 12'h720;
        src40 <= 12'h3e7;
        src41 <= 12'h8d7;
        src42 <= 12'h4d2;
        src43 <= 12'h7e2;
        src44 <= 12'hc09;
        src45 <= 12'hcdd;
        src46 <= 12'hf42;
        src47 <= 12'h320;
        src48 <= 12'h663;
        src49 <= 12'ha26;
        src50 <= 12'hcfe;
        src51 <= 12'h71d;
        src52 <= 12'h77;
        src53 <= 12'h502;
        src54 <= 12'h763;
        src55 <= 12'hc0d;
        src56 <= 12'h7ce;
        src57 <= 12'h53a;
        src58 <= 12'hdc3;
        src59 <= 12'h919;
        src60 <= 12'hb58;
        src61 <= 12'hb9c;
        src62 <= 12'hf51;
        src63 <= 12'h392;
        src64 <= 12'hda2;
        src65 <= 12'h1c5;
        src66 <= 12'hd39;
        src67 <= 12'h785;
        src68 <= 12'h7fc;
        src69 <= 12'hd21;
        src70 <= 12'hc75;
        src71 <= 12'h9ca;
        src72 <= 12'h407;
        src73 <= 12'h7b4;
        src74 <= 12'h96e;
        src75 <= 12'h273;
        src76 <= 12'h14c;
        src77 <= 12'h145;
        src78 <= 12'hbff;
        src79 <= 12'hc62;
        src80 <= 12'hb27;
        src81 <= 12'h74b;
        src82 <= 12'h102;
        src83 <= 12'hc62;
        src84 <= 12'h798;
        src85 <= 12'h354;
        src86 <= 12'h1cf;
        src87 <= 12'h1ac;
        src88 <= 12'h4c1;
        src89 <= 12'h2aa;
        src90 <= 12'h751;
        src91 <= 12'had8;
        src92 <= 12'h57f;
        src93 <= 12'hc5;
        src94 <= 12'h608;
        src95 <= 12'hc1c;
        src96 <= 12'hb87;
        src97 <= 12'h68;
        src98 <= 12'h3a4;
        src99 <= 12'h2bc;
        src100 <= 12'h8cc;
        src101 <= 12'hfb5;
        src102 <= 12'hdf;
        src103 <= 12'h82d;
        src104 <= 12'hcd4;
        src105 <= 12'h175;
        src106 <= 12'h8a6;
        src107 <= 12'h917;
        src108 <= 12'h5f4;
        src109 <= 12'hc0d;
        src110 <= 12'hae4;
        src111 <= 12'h99d;
        src112 <= 12'h69f;
        src113 <= 12'hec4;
        src114 <= 12'h183;
        src115 <= 12'h53c;
        src116 <= 12'h12;
        src117 <= 12'h129;
        src118 <= 12'h647;
        src119 <= 12'hbeb;
        src120 <= 12'h1f3;
        src121 <= 12'hee7;
        src122 <= 12'hfb2;
        src123 <= 12'h4f8;
        src124 <= 12'h215;
        src125 <= 12'h515;
        src126 <= 12'hcab;
        src127 <= 12'hf18;
        src128 <= 12'h1b2;
        src129 <= 12'h524;
        src130 <= 12'ha9e;
        src131 <= 12'hdf6;
        src132 <= 12'he7f;
        src133 <= 12'h2be;
        src134 <= 12'h350;
        src135 <= 12'h259;
        src136 <= 12'h92a;
        src137 <= 12'hc87;
        src138 <= 12'h9d3;
        src139 <= 12'h8f;
        src140 <= 12'h670;
        src141 <= 12'h5cb;
        src142 <= 12'ha2e;
        src143 <= 12'h4d2;
        src144 <= 12'h3c1;
        src145 <= 12'hc6f;
        src146 <= 12'hff5;
        src147 <= 12'hc85;
        src148 <= 12'ha9b;
        src149 <= 12'hae5;
        src150 <= 12'hd26;
        src151 <= 12'he47;
        src152 <= 12'h40c;
        src153 <= 12'h86;
        src154 <= 12'h329;
        src155 <= 12'hfa8;
        src156 <= 12'hb62;
        src157 <= 12'h51a;
        src158 <= 12'h7db;
        src159 <= 12'h168;
        src160 <= 12'hbf7;
        src161 <= 12'h355;
        src162 <= 12'h96b;
        src163 <= 12'h4c3;
        src164 <= 12'hd;
        src165 <= 12'h72c;
        src166 <= 12'h9aa;
        src167 <= 12'h216;
        src168 <= 12'habc;
        src169 <= 12'hbe0;
        src170 <= 12'h3dd;
        src171 <= 12'h54e;
        src172 <= 12'h65e;
        src173 <= 12'hc62;
        src174 <= 12'h1ec;
        src175 <= 12'h6bf;
        src176 <= 12'h8e7;
        src177 <= 12'hb4e;
        src178 <= 12'h9a;
        src179 <= 12'h55e;
        src180 <= 12'hab8;
        src181 <= 12'h6ea;
        src182 <= 12'h1a2;
        src183 <= 12'ha3;
        src184 <= 12'hcc7;
        src185 <= 12'h14e;
        src186 <= 12'ha34;
        src187 <= 12'h4a1;
        src188 <= 12'hbed;
        exp <= 20'h5927b;
        #1
        src0 <= 12'h8c4;
        src1 <= 12'h74f;
        src2 <= 12'h610;
        src3 <= 12'h752;
        src4 <= 12'h667;
        src5 <= 12'h9a5;
        src6 <= 12'hf22;
        src7 <= 12'he5a;
        src8 <= 12'hfc;
        src9 <= 12'h9d1;
        src10 <= 12'hf8;
        src11 <= 12'he0c;
        src12 <= 12'h2f4;
        src13 <= 12'h163;
        src14 <= 12'h527;
        src15 <= 12'hc43;
        src16 <= 12'h985;
        src17 <= 12'h562;
        src18 <= 12'h303;
        src19 <= 12'h12d;
        src20 <= 12'h8cb;
        src21 <= 12'h4ec;
        src22 <= 12'h8b0;
        src23 <= 12'hf76;
        src24 <= 12'hf6;
        src25 <= 12'h582;
        src26 <= 12'h87a;
        src27 <= 12'hf83;
        src28 <= 12'h346;
        src29 <= 12'h730;
        src30 <= 12'hcf;
        src31 <= 12'hb80;
        src32 <= 12'hef3;
        src33 <= 12'hc7e;
        src34 <= 12'hfca;
        src35 <= 12'hb28;
        src36 <= 12'h47d;
        src37 <= 12'h2cb;
        src38 <= 12'heb5;
        src39 <= 12'hf4d;
        src40 <= 12'h5a1;
        src41 <= 12'h9;
        src42 <= 12'h405;
        src43 <= 12'hfb4;
        src44 <= 12'h6b3;
        src45 <= 12'h24a;
        src46 <= 12'h5bc;
        src47 <= 12'ha3d;
        src48 <= 12'h3f6;
        src49 <= 12'h85b;
        src50 <= 12'h668;
        src51 <= 12'h22d;
        src52 <= 12'hf18;
        src53 <= 12'had5;
        src54 <= 12'h566;
        src55 <= 12'ha29;
        src56 <= 12'h29d;
        src57 <= 12'h9f0;
        src58 <= 12'hdf2;
        src59 <= 12'h6a7;
        src60 <= 12'h65f;
        src61 <= 12'h7f1;
        src62 <= 12'hfaf;
        src63 <= 12'h79f;
        src64 <= 12'h448;
        src65 <= 12'h388;
        src66 <= 12'hec4;
        src67 <= 12'hfba;
        src68 <= 12'h653;
        src69 <= 12'hd33;
        src70 <= 12'h895;
        src71 <= 12'h983;
        src72 <= 12'h7c7;
        src73 <= 12'h15e;
        src74 <= 12'hfb;
        src75 <= 12'hbd1;
        src76 <= 12'hd84;
        src77 <= 12'h627;
        src78 <= 12'h3f;
        src79 <= 12'h42d;
        src80 <= 12'hf87;
        src81 <= 12'h207;
        src82 <= 12'he9d;
        src83 <= 12'hbc6;
        src84 <= 12'ha71;
        src85 <= 12'h4ee;
        src86 <= 12'hbc9;
        src87 <= 12'h2c8;
        src88 <= 12'hdc3;
        src89 <= 12'hd16;
        src90 <= 12'h8b;
        src91 <= 12'hd56;
        src92 <= 12'ha67;
        src93 <= 12'h642;
        src94 <= 12'hd79;
        src95 <= 12'h2bc;
        src96 <= 12'hcaf;
        src97 <= 12'h70d;
        src98 <= 12'h1c;
        src99 <= 12'h607;
        src100 <= 12'h205;
        src101 <= 12'h886;
        src102 <= 12'hdc7;
        src103 <= 12'h76a;
        src104 <= 12'ha82;
        src105 <= 12'hdaa;
        src106 <= 12'h8a;
        src107 <= 12'h54c;
        src108 <= 12'h231;
        src109 <= 12'hf34;
        src110 <= 12'h472;
        src111 <= 12'h788;
        src112 <= 12'hd18;
        src113 <= 12'h9bb;
        src114 <= 12'hab4;
        src115 <= 12'hcd9;
        src116 <= 12'h8ae;
        src117 <= 12'h7b3;
        src118 <= 12'hb39;
        src119 <= 12'h494;
        src120 <= 12'h977;
        src121 <= 12'h216;
        src122 <= 12'he52;
        src123 <= 12'h33;
        src124 <= 12'he76;
        src125 <= 12'h59;
        src126 <= 12'ha50;
        src127 <= 12'h138;
        src128 <= 12'hafd;
        src129 <= 12'h48;
        src130 <= 12'h507;
        src131 <= 12'h76a;
        src132 <= 12'hf23;
        src133 <= 12'h6c6;
        src134 <= 12'h132;
        src135 <= 12'hfad;
        src136 <= 12'hb84;
        src137 <= 12'hcc6;
        src138 <= 12'ha79;
        src139 <= 12'hb74;
        src140 <= 12'h5a7;
        src141 <= 12'hd9b;
        src142 <= 12'h17f;
        src143 <= 12'hc66;
        src144 <= 12'h844;
        src145 <= 12'h100;
        src146 <= 12'hfa8;
        src147 <= 12'h8bf;
        src148 <= 12'hd1b;
        src149 <= 12'h824;
        src150 <= 12'h3a6;
        src151 <= 12'h2dd;
        src152 <= 12'h93b;
        src153 <= 12'h8c2;
        src154 <= 12'h7e2;
        src155 <= 12'h19f;
        src156 <= 12'hf6a;
        src157 <= 12'h1c2;
        src158 <= 12'h7d8;
        src159 <= 12'hd83;
        src160 <= 12'h78e;
        src161 <= 12'ha35;
        src162 <= 12'hba;
        src163 <= 12'hbe7;
        src164 <= 12'h847;
        src165 <= 12'hd68;
        src166 <= 12'h68b;
        src167 <= 12'haf6;
        src168 <= 12'he05;
        src169 <= 12'h821;
        src170 <= 12'he69;
        src171 <= 12'h96c;
        src172 <= 12'haf3;
        src173 <= 12'hf95;
        src174 <= 12'habb;
        src175 <= 12'hfb2;
        src176 <= 12'he45;
        src177 <= 12'hfa8;
        src178 <= 12'h6fa;
        src179 <= 12'hd1;
        src180 <= 12'h27a;
        src181 <= 12'he91;
        src182 <= 12'he31;
        src183 <= 12'hb9d;
        src184 <= 12'h270;
        src185 <= 12'h969;
        src186 <= 12'h20c;
        src187 <= 12'hfbd;
        src188 <= 12'h53;
        exp <= 20'h625a1;
        #1
        src0 <= 12'h2d5;
        src1 <= 12'h962;
        src2 <= 12'h305;
        src3 <= 12'h942;
        src4 <= 12'ha90;
        src5 <= 12'hb47;
        src6 <= 12'h1fe;
        src7 <= 12'h94c;
        src8 <= 12'hd0d;
        src9 <= 12'habb;
        src10 <= 12'h777;
        src11 <= 12'h9d5;
        src12 <= 12'h8ca;
        src13 <= 12'hc31;
        src14 <= 12'h111;
        src15 <= 12'h37a;
        src16 <= 12'h48c;
        src17 <= 12'hdc0;
        src18 <= 12'h9e8;
        src19 <= 12'h3c6;
        src20 <= 12'hf33;
        src21 <= 12'h44c;
        src22 <= 12'h9f5;
        src23 <= 12'h182;
        src24 <= 12'h210;
        src25 <= 12'ha29;
        src26 <= 12'h5c6;
        src27 <= 12'he8b;
        src28 <= 12'h9c;
        src29 <= 12'h9b;
        src30 <= 12'h2f5;
        src31 <= 12'hb9c;
        src32 <= 12'h18c;
        src33 <= 12'h185;
        src34 <= 12'hc7;
        src35 <= 12'hbde;
        src36 <= 12'h342;
        src37 <= 12'h6f1;
        src38 <= 12'h70f;
        src39 <= 12'h420;
        src40 <= 12'h9c;
        src41 <= 12'h4ab;
        src42 <= 12'hc61;
        src43 <= 12'hbea;
        src44 <= 12'h2c8;
        src45 <= 12'hba9;
        src46 <= 12'h1f9;
        src47 <= 12'h838;
        src48 <= 12'h521;
        src49 <= 12'hd81;
        src50 <= 12'h4cc;
        src51 <= 12'h1dd;
        src52 <= 12'hd6c;
        src53 <= 12'h6cc;
        src54 <= 12'h8c;
        src55 <= 12'hcfa;
        src56 <= 12'h700;
        src57 <= 12'h4ab;
        src58 <= 12'h6d1;
        src59 <= 12'h81e;
        src60 <= 12'h389;
        src61 <= 12'h7e0;
        src62 <= 12'hf26;
        src63 <= 12'h9e;
        src64 <= 12'hbc4;
        src65 <= 12'h195;
        src66 <= 12'h966;
        src67 <= 12'had0;
        src68 <= 12'h9e0;
        src69 <= 12'h185;
        src70 <= 12'ha25;
        src71 <= 12'hbe;
        src72 <= 12'h845;
        src73 <= 12'h4c9;
        src74 <= 12'he33;
        src75 <= 12'h603;
        src76 <= 12'h1da;
        src77 <= 12'h4f2;
        src78 <= 12'hea5;
        src79 <= 12'h554;
        src80 <= 12'h6b3;
        src81 <= 12'he88;
        src82 <= 12'h755;
        src83 <= 12'h62;
        src84 <= 12'h868;
        src85 <= 12'h473;
        src86 <= 12'h894;
        src87 <= 12'hecb;
        src88 <= 12'hd1a;
        src89 <= 12'hc11;
        src90 <= 12'he2c;
        src91 <= 12'h582;
        src92 <= 12'h687;
        src93 <= 12'hde3;
        src94 <= 12'h39e;
        src95 <= 12'h6ee;
        src96 <= 12'h22d;
        src97 <= 12'hc21;
        src98 <= 12'hdca;
        src99 <= 12'hb0f;
        src100 <= 12'hebe;
        src101 <= 12'h319;
        src102 <= 12'hef1;
        src103 <= 12'h9e;
        src104 <= 12'h1ec;
        src105 <= 12'h66c;
        src106 <= 12'hc5f;
        src107 <= 12'hd5;
        src108 <= 12'h6e7;
        src109 <= 12'h20d;
        src110 <= 12'h2d0;
        src111 <= 12'h904;
        src112 <= 12'hd00;
        src113 <= 12'hb76;
        src114 <= 12'h821;
        src115 <= 12'h869;
        src116 <= 12'h7d8;
        src117 <= 12'h3f8;
        src118 <= 12'h96e;
        src119 <= 12'h63;
        src120 <= 12'h69b;
        src121 <= 12'hc48;
        src122 <= 12'h456;
        src123 <= 12'h1d5;
        src124 <= 12'hed;
        src125 <= 12'h8ce;
        src126 <= 12'he68;
        src127 <= 12'he77;
        src128 <= 12'hd28;
        src129 <= 12'he7;
        src130 <= 12'h71e;
        src131 <= 12'h5eb;
        src132 <= 12'he22;
        src133 <= 12'h798;
        src134 <= 12'hf3a;
        src135 <= 12'ha13;
        src136 <= 12'h249;
        src137 <= 12'h4d8;
        src138 <= 12'h31e;
        src139 <= 12'h904;
        src140 <= 12'h2f7;
        src141 <= 12'h3f0;
        src142 <= 12'hd26;
        src143 <= 12'h716;
        src144 <= 12'hed2;
        src145 <= 12'ha1f;
        src146 <= 12'hbac;
        src147 <= 12'ha2d;
        src148 <= 12'h743;
        src149 <= 12'h703;
        src150 <= 12'hac5;
        src151 <= 12'h2f4;
        src152 <= 12'h5b1;
        src153 <= 12'ha79;
        src154 <= 12'h575;
        src155 <= 12'hbbf;
        src156 <= 12'hdd3;
        src157 <= 12'h9ff;
        src158 <= 12'h32c;
        src159 <= 12'h87c;
        src160 <= 12'hcb9;
        src161 <= 12'hc36;
        src162 <= 12'h3de;
        src163 <= 12'h652;
        src164 <= 12'h68;
        src165 <= 12'h51a;
        src166 <= 12'h619;
        src167 <= 12'h6b1;
        src168 <= 12'h211;
        src169 <= 12'h3b3;
        src170 <= 12'h156;
        src171 <= 12'h87e;
        src172 <= 12'h156;
        src173 <= 12'h40;
        src174 <= 12'hd48;
        src175 <= 12'hbc0;
        src176 <= 12'h726;
        src177 <= 12'hb86;
        src178 <= 12'hadc;
        src179 <= 12'hb6e;
        src180 <= 12'h9ca;
        src181 <= 12'h1be;
        src182 <= 12'ha5d;
        src183 <= 12'h10c;
        src184 <= 12'h8fb;
        src185 <= 12'h33c;
        src186 <= 12'hc3a;
        src187 <= 12'h830;
        src188 <= 12'hbc2;
        exp <= 20'h57dad;
        #1
        src0 <= 12'h41d;
        src1 <= 12'h79c;
        src2 <= 12'h201;
        src3 <= 12'h9f8;
        src4 <= 12'h5a1;
        src5 <= 12'h9be;
        src6 <= 12'h849;
        src7 <= 12'h526;
        src8 <= 12'h969;
        src9 <= 12'h62;
        src10 <= 12'h7ca;
        src11 <= 12'hebe;
        src12 <= 12'hd08;
        src13 <= 12'h5c2;
        src14 <= 12'hbcd;
        src15 <= 12'h7ca;
        src16 <= 12'hfe7;
        src17 <= 12'hbd1;
        src18 <= 12'h702;
        src19 <= 12'hd2e;
        src20 <= 12'h718;
        src21 <= 12'h287;
        src22 <= 12'h85f;
        src23 <= 12'h52a;
        src24 <= 12'h234;
        src25 <= 12'h214;
        src26 <= 12'h9e7;
        src27 <= 12'hfc5;
        src28 <= 12'h2bc;
        src29 <= 12'h3ac;
        src30 <= 12'h49b;
        src31 <= 12'hadf;
        src32 <= 12'h119;
        src33 <= 12'h8c8;
        src34 <= 12'h29f;
        src35 <= 12'h576;
        src36 <= 12'hf32;
        src37 <= 12'h402;
        src38 <= 12'hcf0;
        src39 <= 12'he09;
        src40 <= 12'h3c;
        src41 <= 12'h46b;
        src42 <= 12'h965;
        src43 <= 12'h97b;
        src44 <= 12'hc6f;
        src45 <= 12'hb87;
        src46 <= 12'h11e;
        src47 <= 12'h54c;
        src48 <= 12'hbe5;
        src49 <= 12'hf1;
        src50 <= 12'hc4e;
        src51 <= 12'h80d;
        src52 <= 12'h4ab;
        src53 <= 12'hbe4;
        src54 <= 12'hb4f;
        src55 <= 12'hb3e;
        src56 <= 12'h7c4;
        src57 <= 12'hc9b;
        src58 <= 12'h93d;
        src59 <= 12'h7c6;
        src60 <= 12'h96d;
        src61 <= 12'h4e9;
        src62 <= 12'h9d3;
        src63 <= 12'he53;
        src64 <= 12'haa5;
        src65 <= 12'h8b9;
        src66 <= 12'hbeb;
        src67 <= 12'h4d9;
        src68 <= 12'h698;
        src69 <= 12'hd1b;
        src70 <= 12'h308;
        src71 <= 12'h32c;
        src72 <= 12'h74e;
        src73 <= 12'h50;
        src74 <= 12'h739;
        src75 <= 12'h11e;
        src76 <= 12'h116;
        src77 <= 12'hfcf;
        src78 <= 12'h86;
        src79 <= 12'hef0;
        src80 <= 12'ha3c;
        src81 <= 12'hfb;
        src82 <= 12'head;
        src83 <= 12'h21a;
        src84 <= 12'he3c;
        src85 <= 12'h1ed;
        src86 <= 12'h5e4;
        src87 <= 12'h3f8;
        src88 <= 12'h5a1;
        src89 <= 12'hc04;
        src90 <= 12'h331;
        src91 <= 12'h50;
        src92 <= 12'h69a;
        src93 <= 12'h8ac;
        src94 <= 12'ha56;
        src95 <= 12'h591;
        src96 <= 12'h5c9;
        src97 <= 12'h62b;
        src98 <= 12'hc19;
        src99 <= 12'h1e9;
        src100 <= 12'ha8b;
        src101 <= 12'h637;
        src102 <= 12'hc39;
        src103 <= 12'h18c;
        src104 <= 12'hbbf;
        src105 <= 12'ha55;
        src106 <= 12'h83a;
        src107 <= 12'h6c7;
        src108 <= 12'h423;
        src109 <= 12'hd8d;
        src110 <= 12'h73f;
        src111 <= 12'h1fb;
        src112 <= 12'h6d1;
        src113 <= 12'hb96;
        src114 <= 12'h5c4;
        src115 <= 12'hdf;
        src116 <= 12'h472;
        src117 <= 12'h187;
        src118 <= 12'h3c1;
        src119 <= 12'h102;
        src120 <= 12'h9ba;
        src121 <= 12'h5af;
        src122 <= 12'h4d5;
        src123 <= 12'h306;
        src124 <= 12'hb15;
        src125 <= 12'h5a6;
        src126 <= 12'h729;
        src127 <= 12'hd6d;
        src128 <= 12'h219;
        src129 <= 12'h283;
        src130 <= 12'hd0c;
        src131 <= 12'h229;
        src132 <= 12'h773;
        src133 <= 12'hf38;
        src134 <= 12'h622;
        src135 <= 12'h6e3;
        src136 <= 12'h96f;
        src137 <= 12'hfe7;
        src138 <= 12'hd31;
        src139 <= 12'h438;
        src140 <= 12'h29;
        src141 <= 12'hfee;
        src142 <= 12'h58;
        src143 <= 12'hf4b;
        src144 <= 12'h900;
        src145 <= 12'hbcd;
        src146 <= 12'h47c;
        src147 <= 12'h495;
        src148 <= 12'hb90;
        src149 <= 12'haf8;
        src150 <= 12'h55a;
        src151 <= 12'h530;
        src152 <= 12'h952;
        src153 <= 12'hbc1;
        src154 <= 12'h90c;
        src155 <= 12'hd49;
        src156 <= 12'h74f;
        src157 <= 12'h81e;
        src158 <= 12'hf29;
        src159 <= 12'h770;
        src160 <= 12'hf14;
        src161 <= 12'h815;
        src162 <= 12'h731;
        src163 <= 12'he1c;
        src164 <= 12'h83b;
        src165 <= 12'hbab;
        src166 <= 12'h803;
        src167 <= 12'h721;
        src168 <= 12'h50d;
        src169 <= 12'h879;
        src170 <= 12'hbc3;
        src171 <= 12'h647;
        src172 <= 12'h712;
        src173 <= 12'ha3f;
        src174 <= 12'hb8c;
        src175 <= 12'h6c6;
        src176 <= 12'h7f6;
        src177 <= 12'h378;
        src178 <= 12'hed4;
        src179 <= 12'h184;
        src180 <= 12'h11a;
        src181 <= 12'h92c;
        src182 <= 12'ha98;
        src183 <= 12'h976;
        src184 <= 12'heab;
        src185 <= 12'h1db;
        src186 <= 12'hc6a;
        src187 <= 12'h70e;
        src188 <= 12'he4;
        exp <= 20'h5b5dc;
        #1
        src0 <= 12'h5f0;
        src1 <= 12'h6d6;
        src2 <= 12'hf85;
        src3 <= 12'he05;
        src4 <= 12'h69b;
        src5 <= 12'hc35;
        src6 <= 12'hd63;
        src7 <= 12'hb90;
        src8 <= 12'h931;
        src9 <= 12'hda4;
        src10 <= 12'h4f3;
        src11 <= 12'h427;
        src12 <= 12'heee;
        src13 <= 12'hf87;
        src14 <= 12'h143;
        src15 <= 12'h351;
        src16 <= 12'h839;
        src17 <= 12'hb5f;
        src18 <= 12'h6c;
        src19 <= 12'hb80;
        src20 <= 12'h265;
        src21 <= 12'hda;
        src22 <= 12'h9b1;
        src23 <= 12'hbfd;
        src24 <= 12'h5e8;
        src25 <= 12'h540;
        src26 <= 12'h8fb;
        src27 <= 12'h65f;
        src28 <= 12'he3e;
        src29 <= 12'hefc;
        src30 <= 12'hfa0;
        src31 <= 12'h955;
        src32 <= 12'hdeb;
        src33 <= 12'h46c;
        src34 <= 12'hcd0;
        src35 <= 12'hda2;
        src36 <= 12'h2ee;
        src37 <= 12'h3ea;
        src38 <= 12'h84d;
        src39 <= 12'hf5c;
        src40 <= 12'h55b;
        src41 <= 12'h47a;
        src42 <= 12'hf12;
        src43 <= 12'he5e;
        src44 <= 12'hc94;
        src45 <= 12'hf10;
        src46 <= 12'h738;
        src47 <= 12'h98b;
        src48 <= 12'h65;
        src49 <= 12'h641;
        src50 <= 12'h77e;
        src51 <= 12'ha1d;
        src52 <= 12'h1bb;
        src53 <= 12'h54f;
        src54 <= 12'h108;
        src55 <= 12'h78e;
        src56 <= 12'h49d;
        src57 <= 12'hadc;
        src58 <= 12'hfd5;
        src59 <= 12'h68c;
        src60 <= 12'h812;
        src61 <= 12'h2b2;
        src62 <= 12'ha00;
        src63 <= 12'h9cf;
        src64 <= 12'hdd2;
        src65 <= 12'h4a8;
        src66 <= 12'hb55;
        src67 <= 12'he24;
        src68 <= 12'h484;
        src69 <= 12'hd1c;
        src70 <= 12'h853;
        src71 <= 12'h64b;
        src72 <= 12'h7e;
        src73 <= 12'h70c;
        src74 <= 12'h8ce;
        src75 <= 12'h483;
        src76 <= 12'hd7a;
        src77 <= 12'h90d;
        src78 <= 12'h942;
        src79 <= 12'h28d;
        src80 <= 12'he18;
        src81 <= 12'ha7a;
        src82 <= 12'h532;
        src83 <= 12'h6fd;
        src84 <= 12'h5b9;
        src85 <= 12'h586;
        src86 <= 12'he0c;
        src87 <= 12'h355;
        src88 <= 12'h6ca;
        src89 <= 12'h110;
        src90 <= 12'had2;
        src91 <= 12'habb;
        src92 <= 12'h486;
        src93 <= 12'h515;
        src94 <= 12'h988;
        src95 <= 12'h788;
        src96 <= 12'h550;
        src97 <= 12'h747;
        src98 <= 12'hcd2;
        src99 <= 12'h12f;
        src100 <= 12'h4ae;
        src101 <= 12'h7a4;
        src102 <= 12'h871;
        src103 <= 12'hb66;
        src104 <= 12'h67b;
        src105 <= 12'h9c5;
        src106 <= 12'hc8b;
        src107 <= 12'h3d8;
        src108 <= 12'h5ec;
        src109 <= 12'h725;
        src110 <= 12'h9e2;
        src111 <= 12'h41c;
        src112 <= 12'hed0;
        src113 <= 12'h2bc;
        src114 <= 12'hfaf;
        src115 <= 12'hb2f;
        src116 <= 12'h97;
        src117 <= 12'h956;
        src118 <= 12'hd05;
        src119 <= 12'h79a;
        src120 <= 12'h54b;
        src121 <= 12'h7cd;
        src122 <= 12'h594;
        src123 <= 12'h5a8;
        src124 <= 12'h85d;
        src125 <= 12'h9cb;
        src126 <= 12'hcc6;
        src127 <= 12'hdee;
        src128 <= 12'h17a;
        src129 <= 12'h23c;
        src130 <= 12'h9dd;
        src131 <= 12'hb1;
        src132 <= 12'h381;
        src133 <= 12'h8d0;
        src134 <= 12'h656;
        src135 <= 12'h469;
        src136 <= 12'hd9e;
        src137 <= 12'hb14;
        src138 <= 12'hb31;
        src139 <= 12'hba5;
        src140 <= 12'hf3e;
        src141 <= 12'h1c9;
        src142 <= 12'h8e7;
        src143 <= 12'hb0;
        src144 <= 12'hf55;
        src145 <= 12'he41;
        src146 <= 12'hca7;
        src147 <= 12'h984;
        src148 <= 12'h1b5;
        src149 <= 12'hc5c;
        src150 <= 12'h9e2;
        src151 <= 12'h161;
        src152 <= 12'h93e;
        src153 <= 12'hce;
        src154 <= 12'hc96;
        src155 <= 12'h1f;
        src156 <= 12'hbb1;
        src157 <= 12'h52a;
        src158 <= 12'h493;
        src159 <= 12'h3a7;
        src160 <= 12'hfe5;
        src161 <= 12'h84f;
        src162 <= 12'h7fc;
        src163 <= 12'h486;
        src164 <= 12'hee7;
        src165 <= 12'h1ab;
        src166 <= 12'he0a;
        src167 <= 12'he56;
        src168 <= 12'hcc0;
        src169 <= 12'hce0;
        src170 <= 12'h4f;
        src171 <= 12'h9b3;
        src172 <= 12'h86a;
        src173 <= 12'h6d7;
        src174 <= 12'h7fa;
        src175 <= 12'hcf7;
        src176 <= 12'hd1;
        src177 <= 12'hf12;
        src178 <= 12'hef2;
        src179 <= 12'hab5;
        src180 <= 12'h57a;
        src181 <= 12'hd4;
        src182 <= 12'h6c4;
        src183 <= 12'hf26;
        src184 <= 12'hd51;
        src185 <= 12'h152;
        src186 <= 12'h168;
        src187 <= 12'hdc8;
        src188 <= 12'hcba;
        exp <= 20'h6270f;
        #1
        $finish;
    end
endmodule

