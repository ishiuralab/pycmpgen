module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    compressor2_1_64_16 compressor2_1_64_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_64_16(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [0:0] comp_out20;
    wire [0:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    rowadder2_1_22 rowadder2_1inst(
        .src0({comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [19:0] stage1_0;
   wire [29:0] stage1_1;
   wire [23:0] stage1_2;
   wire [26:0] stage1_3;
   wire [39:0] stage1_4;
   wire [28:0] stage1_5;
   wire [26:0] stage1_6;
   wire [22:0] stage1_7;
   wire [28:0] stage1_8;
   wire [29:0] stage1_9;
   wire [27:0] stage1_10;
   wire [23:0] stage1_11;
   wire [29:0] stage1_12;
   wire [32:0] stage1_13;
   wire [24:0] stage1_14;
   wire [23:0] stage1_15;
   wire [18:0] stage1_16;
   wire [9:0] stage1_17;
   wire [3:0] stage2_0;
   wire [21:0] stage2_1;
   wire [7:0] stage2_2;
   wire [10:0] stage2_3;
   wire [15:0] stage2_4;
   wire [17:0] stage2_5;
   wire [11:0] stage2_6;
   wire [11:0] stage2_7;
   wire [15:0] stage2_8;
   wire [7:0] stage2_9;
   wire [12:0] stage2_10;
   wire [17:0] stage2_11;
   wire [7:0] stage2_12;
   wire [18:0] stage2_13;
   wire [23:0] stage2_14;
   wire [7:0] stage2_15;
   wire [12:0] stage2_16;
   wire [5:0] stage2_17;
   wire [3:0] stage2_18;
   wire [1:0] stage2_19;
   wire [1:0] stage3_0;
   wire [6:0] stage3_1;
   wire [3:0] stage3_2;
   wire [6:0] stage3_3;
   wire [5:0] stage3_4;
   wire [9:0] stage3_5;
   wire [4:0] stage3_6;
   wire [3:0] stage3_7;
   wire [7:0] stage3_8;
   wire [6:0] stage3_9;
   wire [2:0] stage3_10;
   wire [6:0] stage3_11;
   wire [6:0] stage3_12;
   wire [4:0] stage3_13;
   wire [13:0] stage3_14;
   wire [6:0] stage3_15;
   wire [4:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [2:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [5:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [3:0] stage4_8;
   wire [3:0] stage4_9;
   wire [3:0] stage4_10;
   wire [1:0] stage4_11;
   wire [2:0] stage4_12;
   wire [2:0] stage4_13;
   wire [8:0] stage4_14;
   wire [2:0] stage4_15;
   wire [2:0] stage4_16;
   wire [3:0] stage4_17;
   wire [1:0] stage4_18;
   wire [3:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [0:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[50]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc615_5 gpc18 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[51]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[9],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[13],stage1_4[22]}
   );
   gpc615_5 gpc23 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_5[6]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[14],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[7]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[15],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_5[8]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[16],stage1_4[25]}
   );
   gpc615_5 gpc26 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50]},
      {stage0_5[9]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[12],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[13],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[14],stage1_5[22]}
   );
   gpc606_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[15],stage1_5[23]}
   );
   gpc606_5 gpc33 (
      {stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc34 (
      {stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[17],stage1_5[25]}
   );
   gpc615_5 gpc35 (
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_6[43]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[18],stage1_5[26]}
   );
   gpc615_5 gpc36 (
      {stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[19]}
   );
   gpc615_5 gpc37 (
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[17],stage1_7[18],stage1_6[20]}
   );
   gpc615_5 gpc38 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[18],stage1_7[19],stage1_6[21]}
   );
   gpc615_5 gpc39 (
      {stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[12],stage1_8[19],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[4],stage1_9[13],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[5],stage1_9[14],stage1_8[21]}
   );
   gpc606_5 gpc42 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[6],stage1_9[15],stage1_8[22]}
   );
   gpc606_5 gpc43 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[7],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc44 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_9[6]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[8],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc45 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_9[7]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[9],stage1_9[18],stage1_8[25]}
   );
   gpc615_5 gpc46 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_9[8]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[10],stage1_9[19],stage1_8[26]}
   );
   gpc615_5 gpc47 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62]},
      {stage0_9[9]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[11],stage1_9[20],stage1_8[27]}
   );
   gpc606_5 gpc48 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc52 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc53 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[17],stage1_9[26]}
   );
   gpc606_5 gpc54 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[18],stage1_9[27]}
   );
   gpc606_5 gpc55 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[19],stage1_9[28]}
   );
   gpc606_5 gpc56 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[16],stage1_11[17],stage1_10[20],stage1_9[29]}
   );
   gpc606_5 gpc57 (
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[17],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc58 (
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58]},
      {stage0_11[54]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[18],stage1_11[19],stage1_10[22]}
   );
   gpc606_5 gpc59 (
      {stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[11],stage1_12[19],stage1_11[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[3],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc61 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[4],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc62 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[5],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc63 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[6],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc64 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[7],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc65 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[8],stage1_13[17],stage1_12[25]}
   );
   gpc615_5 gpc66 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_13[6]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[9],stage1_13[18],stage1_12[26]}
   );
   gpc615_5 gpc67 (
      {stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage0_13[7]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[10],stage1_13[19],stage1_12[27]}
   );
   gpc615_5 gpc68 (
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_13[8]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[11],stage1_13[20],stage1_12[28]}
   );
   gpc606_5 gpc69 (
      {stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[12],stage1_13[21]}
   );
   gpc606_5 gpc70 (
      {stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[13],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[14],stage1_13[23]}
   );
   gpc615_5 gpc72 (
      {stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage0_14[54]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[15],stage1_13[24]}
   );
   gpc615_5 gpc73 (
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36]},
      {stage0_14[55]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[16],stage1_13[25]}
   );
   gpc615_5 gpc74 (
      {stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_14[56]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[17],stage1_13[26]}
   );
   gpc615_5 gpc75 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_14[57]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[18],stage1_13[27]}
   );
   gpc615_5 gpc76 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage0_14[58]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[19],stage1_13[28]}
   );
   gpc615_5 gpc77 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56]},
      {stage0_14[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[17],stage1_15[18],stage1_14[20],stage1_13[29]}
   );
   gpc615_5 gpc78 (
      {stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_14[60]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[18],stage1_15[19],stage1_14[21],stage1_13[30]}
   );
   gpc1_1 gpc79 (
      {stage0_0[53]},
      {stage1_0[9]}
   );
   gpc1_1 gpc80 (
      {stage0_0[54]},
      {stage1_0[10]}
   );
   gpc1_1 gpc81 (
      {stage0_0[55]},
      {stage1_0[11]}
   );
   gpc1_1 gpc82 (
      {stage0_0[56]},
      {stage1_0[12]}
   );
   gpc1_1 gpc83 (
      {stage0_0[57]},
      {stage1_0[13]}
   );
   gpc1_1 gpc84 (
      {stage0_0[58]},
      {stage1_0[14]}
   );
   gpc1_1 gpc85 (
      {stage0_0[59]},
      {stage1_0[15]}
   );
   gpc1_1 gpc86 (
      {stage0_0[60]},
      {stage1_0[16]}
   );
   gpc1_1 gpc87 (
      {stage0_0[61]},
      {stage1_0[17]}
   );
   gpc1_1 gpc88 (
      {stage0_0[62]},
      {stage1_0[18]}
   );
   gpc1_1 gpc89 (
      {stage0_0[63]},
      {stage1_0[19]}
   );
   gpc1_1 gpc90 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc91 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc92 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc93 (
      {stage0_1[54]},
      {stage1_1[20]}
   );
   gpc1_1 gpc94 (
      {stage0_1[55]},
      {stage1_1[21]}
   );
   gpc1_1 gpc95 (
      {stage0_1[56]},
      {stage1_1[22]}
   );
   gpc1_1 gpc96 (
      {stage0_1[57]},
      {stage1_1[23]}
   );
   gpc1_1 gpc97 (
      {stage0_1[58]},
      {stage1_1[24]}
   );
   gpc1_1 gpc98 (
      {stage0_1[59]},
      {stage1_1[25]}
   );
   gpc1_1 gpc99 (
      {stage0_1[60]},
      {stage1_1[26]}
   );
   gpc1_1 gpc100 (
      {stage0_1[61]},
      {stage1_1[27]}
   );
   gpc1_1 gpc101 (
      {stage0_1[62]},
      {stage1_1[28]}
   );
   gpc1_1 gpc102 (
      {stage0_1[63]},
      {stage1_1[29]}
   );
   gpc1_1 gpc103 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc104 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc105 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc106 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc107 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc108 (
      {stage0_3[57]},
      {stage1_3[20]}
   );
   gpc1_1 gpc109 (
      {stage0_3[58]},
      {stage1_3[21]}
   );
   gpc1_1 gpc110 (
      {stage0_3[59]},
      {stage1_3[22]}
   );
   gpc1_1 gpc111 (
      {stage0_3[60]},
      {stage1_3[23]}
   );
   gpc1_1 gpc112 (
      {stage0_3[61]},
      {stage1_3[24]}
   );
   gpc1_1 gpc113 (
      {stage0_3[62]},
      {stage1_3[25]}
   );
   gpc1_1 gpc114 (
      {stage0_3[63]},
      {stage1_3[26]}
   );
   gpc1_1 gpc115 (
      {stage0_4[51]},
      {stage1_4[27]}
   );
   gpc1_1 gpc116 (
      {stage0_4[52]},
      {stage1_4[28]}
   );
   gpc1_1 gpc117 (
      {stage0_4[53]},
      {stage1_4[29]}
   );
   gpc1_1 gpc118 (
      {stage0_4[54]},
      {stage1_4[30]}
   );
   gpc1_1 gpc119 (
      {stage0_4[55]},
      {stage1_4[31]}
   );
   gpc1_1 gpc120 (
      {stage0_4[56]},
      {stage1_4[32]}
   );
   gpc1_1 gpc121 (
      {stage0_4[57]},
      {stage1_4[33]}
   );
   gpc1_1 gpc122 (
      {stage0_4[58]},
      {stage1_4[34]}
   );
   gpc1_1 gpc123 (
      {stage0_4[59]},
      {stage1_4[35]}
   );
   gpc1_1 gpc124 (
      {stage0_4[60]},
      {stage1_4[36]}
   );
   gpc1_1 gpc125 (
      {stage0_4[61]},
      {stage1_4[37]}
   );
   gpc1_1 gpc126 (
      {stage0_4[62]},
      {stage1_4[38]}
   );
   gpc1_1 gpc127 (
      {stage0_4[63]},
      {stage1_4[39]}
   );
   gpc1_1 gpc128 (
      {stage0_5[62]},
      {stage1_5[27]}
   );
   gpc1_1 gpc129 (
      {stage0_5[63]},
      {stage1_5[28]}
   );
   gpc1_1 gpc130 (
      {stage0_6[59]},
      {stage1_6[22]}
   );
   gpc1_1 gpc131 (
      {stage0_6[60]},
      {stage1_6[23]}
   );
   gpc1_1 gpc132 (
      {stage0_6[61]},
      {stage1_6[24]}
   );
   gpc1_1 gpc133 (
      {stage0_6[62]},
      {stage1_6[25]}
   );
   gpc1_1 gpc134 (
      {stage0_6[63]},
      {stage1_6[26]}
   );
   gpc1_1 gpc135 (
      {stage0_7[62]},
      {stage1_7[21]}
   );
   gpc1_1 gpc136 (
      {stage0_7[63]},
      {stage1_7[22]}
   );
   gpc1_1 gpc137 (
      {stage0_8[63]},
      {stage1_8[28]}
   );
   gpc1_1 gpc138 (
      {stage0_10[59]},
      {stage1_10[23]}
   );
   gpc1_1 gpc139 (
      {stage0_10[60]},
      {stage1_10[24]}
   );
   gpc1_1 gpc140 (
      {stage0_10[61]},
      {stage1_10[25]}
   );
   gpc1_1 gpc141 (
      {stage0_10[62]},
      {stage1_10[26]}
   );
   gpc1_1 gpc142 (
      {stage0_10[63]},
      {stage1_10[27]}
   );
   gpc1_1 gpc143 (
      {stage0_11[61]},
      {stage1_11[21]}
   );
   gpc1_1 gpc144 (
      {stage0_11[62]},
      {stage1_11[22]}
   );
   gpc1_1 gpc145 (
      {stage0_11[63]},
      {stage1_11[23]}
   );
   gpc1_1 gpc146 (
      {stage0_12[63]},
      {stage1_12[29]}
   );
   gpc1_1 gpc147 (
      {stage0_13[62]},
      {stage1_13[31]}
   );
   gpc1_1 gpc148 (
      {stage0_13[63]},
      {stage1_13[32]}
   );
   gpc1_1 gpc149 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc150 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc151 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc152 (
      {stage0_15[60]},
      {stage1_15[20]}
   );
   gpc1_1 gpc153 (
      {stage0_15[61]},
      {stage1_15[21]}
   );
   gpc1_1 gpc154 (
      {stage0_15[62]},
      {stage1_15[22]}
   );
   gpc1_1 gpc155 (
      {stage0_15[63]},
      {stage1_15[23]}
   );
   gpc2135_5 gpc156 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc157 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc158 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc159 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc160 (
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_3[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc161 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage1_3[9]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc162 (
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_3[10]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc163 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[11]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc164 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[4],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc165 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[25]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[5],stage2_5[5],stage2_4[9],stage2_3[9]}
   );
   gpc615_5 gpc166 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[26]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[6],stage2_5[6],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc167 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31]},
      {stage1_5[18]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[7],stage2_5[7],stage2_4[11]}
   );
   gpc615_5 gpc168 (
      {stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36]},
      {stage1_5[19]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[8],stage2_5[8],stage2_4[12]}
   );
   gpc615_5 gpc169 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[0]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[5],stage2_6[9]}
   );
   gpc615_5 gpc170 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[1]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[6],stage2_6[10]}
   );
   gpc615_5 gpc171 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[2]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[4],stage2_7[7],stage2_6[11]}
   );
   gpc615_5 gpc172 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[3],stage2_8[5],stage2_7[8]}
   );
   gpc615_5 gpc173 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[4],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc174 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[5],stage2_8[7],stage2_7[10]}
   );
   gpc615_5 gpc175 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[6],stage2_8[8],stage2_7[11]}
   );
   gpc606_5 gpc176 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[4],stage2_10[7],stage2_9[7]}
   );
   gpc606_5 gpc177 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc178 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc179 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[7],stage2_10[10]}
   );
   gpc606_5 gpc180 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[8],stage2_10[11]}
   );
   gpc606_5 gpc181 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], 1'b0, 1'b0},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[9],stage2_10[12]}
   );
   gpc606_5 gpc182 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[10]}
   );
   gpc606_5 gpc183 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[11]}
   );
   gpc606_5 gpc184 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[2],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc185 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[3],stage2_14[8],stage2_13[9]}
   );
   gpc606_5 gpc186 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[4],stage2_14[9]}
   );
   gpc606_5 gpc187 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[5],stage2_14[10]}
   );
   gpc606_5 gpc188 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[6]}
   );
   gpc606_5 gpc189 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], 1'b0, 1'b0},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[7]}
   );
   gpc1_1 gpc190 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc191 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc192 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc193 (
      {stage1_1[15]},
      {stage2_1[7]}
   );
   gpc1_1 gpc194 (
      {stage1_1[16]},
      {stage2_1[8]}
   );
   gpc1_1 gpc195 (
      {stage1_1[17]},
      {stage2_1[9]}
   );
   gpc1_1 gpc196 (
      {stage1_1[18]},
      {stage2_1[10]}
   );
   gpc1_1 gpc197 (
      {stage1_1[19]},
      {stage2_1[11]}
   );
   gpc1_1 gpc198 (
      {stage1_1[20]},
      {stage2_1[12]}
   );
   gpc1_1 gpc199 (
      {stage1_1[21]},
      {stage2_1[13]}
   );
   gpc1_1 gpc200 (
      {stage1_1[22]},
      {stage2_1[14]}
   );
   gpc1_1 gpc201 (
      {stage1_1[23]},
      {stage2_1[15]}
   );
   gpc1_1 gpc202 (
      {stage1_1[24]},
      {stage2_1[16]}
   );
   gpc1_1 gpc203 (
      {stage1_1[25]},
      {stage2_1[17]}
   );
   gpc1_1 gpc204 (
      {stage1_1[26]},
      {stage2_1[18]}
   );
   gpc1_1 gpc205 (
      {stage1_1[27]},
      {stage2_1[19]}
   );
   gpc1_1 gpc206 (
      {stage1_1[28]},
      {stage2_1[20]}
   );
   gpc1_1 gpc207 (
      {stage1_1[29]},
      {stage2_1[21]}
   );
   gpc1_1 gpc208 (
      {stage1_4[37]},
      {stage2_4[13]}
   );
   gpc1_1 gpc209 (
      {stage1_4[38]},
      {stage2_4[14]}
   );
   gpc1_1 gpc210 (
      {stage1_4[39]},
      {stage2_4[15]}
   );
   gpc1_1 gpc211 (
      {stage1_5[20]},
      {stage2_5[9]}
   );
   gpc1_1 gpc212 (
      {stage1_5[21]},
      {stage2_5[10]}
   );
   gpc1_1 gpc213 (
      {stage1_5[22]},
      {stage2_5[11]}
   );
   gpc1_1 gpc214 (
      {stage1_5[23]},
      {stage2_5[12]}
   );
   gpc1_1 gpc215 (
      {stage1_5[24]},
      {stage2_5[13]}
   );
   gpc1_1 gpc216 (
      {stage1_5[25]},
      {stage2_5[14]}
   );
   gpc1_1 gpc217 (
      {stage1_5[26]},
      {stage2_5[15]}
   );
   gpc1_1 gpc218 (
      {stage1_5[27]},
      {stage2_5[16]}
   );
   gpc1_1 gpc219 (
      {stage1_5[28]},
      {stage2_5[17]}
   );
   gpc1_1 gpc220 (
      {stage1_8[22]},
      {stage2_8[9]}
   );
   gpc1_1 gpc221 (
      {stage1_8[23]},
      {stage2_8[10]}
   );
   gpc1_1 gpc222 (
      {stage1_8[24]},
      {stage2_8[11]}
   );
   gpc1_1 gpc223 (
      {stage1_8[25]},
      {stage2_8[12]}
   );
   gpc1_1 gpc224 (
      {stage1_8[26]},
      {stage2_8[13]}
   );
   gpc1_1 gpc225 (
      {stage1_8[27]},
      {stage2_8[14]}
   );
   gpc1_1 gpc226 (
      {stage1_8[28]},
      {stage2_8[15]}
   );
   gpc1_1 gpc227 (
      {stage1_11[18]},
      {stage2_11[12]}
   );
   gpc1_1 gpc228 (
      {stage1_11[19]},
      {stage2_11[13]}
   );
   gpc1_1 gpc229 (
      {stage1_11[20]},
      {stage2_11[14]}
   );
   gpc1_1 gpc230 (
      {stage1_11[21]},
      {stage2_11[15]}
   );
   gpc1_1 gpc231 (
      {stage1_11[22]},
      {stage2_11[16]}
   );
   gpc1_1 gpc232 (
      {stage1_11[23]},
      {stage2_11[17]}
   );
   gpc1_1 gpc233 (
      {stage1_13[24]},
      {stage2_13[10]}
   );
   gpc1_1 gpc234 (
      {stage1_13[25]},
      {stage2_13[11]}
   );
   gpc1_1 gpc235 (
      {stage1_13[26]},
      {stage2_13[12]}
   );
   gpc1_1 gpc236 (
      {stage1_13[27]},
      {stage2_13[13]}
   );
   gpc1_1 gpc237 (
      {stage1_13[28]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[29]},
      {stage2_13[15]}
   );
   gpc1_1 gpc239 (
      {stage1_13[30]},
      {stage2_13[16]}
   );
   gpc1_1 gpc240 (
      {stage1_13[31]},
      {stage2_13[17]}
   );
   gpc1_1 gpc241 (
      {stage1_13[32]},
      {stage2_13[18]}
   );
   gpc1_1 gpc242 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc243 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc244 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc245 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc246 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc247 (
      {stage1_14[17]},
      {stage2_14[16]}
   );
   gpc1_1 gpc248 (
      {stage1_14[18]},
      {stage2_14[17]}
   );
   gpc1_1 gpc249 (
      {stage1_14[19]},
      {stage2_14[18]}
   );
   gpc1_1 gpc250 (
      {stage1_14[20]},
      {stage2_14[19]}
   );
   gpc1_1 gpc251 (
      {stage1_14[21]},
      {stage2_14[20]}
   );
   gpc1_1 gpc252 (
      {stage1_14[22]},
      {stage2_14[21]}
   );
   gpc1_1 gpc253 (
      {stage1_14[23]},
      {stage2_14[22]}
   );
   gpc1_1 gpc254 (
      {stage1_14[24]},
      {stage2_14[23]}
   );
   gpc1_1 gpc255 (
      {stage1_16[12]},
      {stage2_16[6]}
   );
   gpc1_1 gpc256 (
      {stage1_16[13]},
      {stage2_16[7]}
   );
   gpc1_1 gpc257 (
      {stage1_16[14]},
      {stage2_16[8]}
   );
   gpc1_1 gpc258 (
      {stage1_16[15]},
      {stage2_16[9]}
   );
   gpc1_1 gpc259 (
      {stage1_16[16]},
      {stage2_16[10]}
   );
   gpc1_1 gpc260 (
      {stage1_16[17]},
      {stage2_16[11]}
   );
   gpc1_1 gpc261 (
      {stage1_16[18]},
      {stage2_16[12]}
   );
   gpc1163_5 gpc262 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc263 (
      {stage2_0[3], 1'b0, 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc264 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc265 (
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc266 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[0]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4]}
   );
   gpc615_5 gpc267 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[1]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5]}
   );
   gpc606_5 gpc268 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[4]}
   );
   gpc606_5 gpc269 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12], stage2_5[13]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[5]}
   );
   gpc1163_5 gpc270 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[0]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[2],stage3_8[4]}
   );
   gpc606_5 gpc271 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7], stage2_8[8]},
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc272 (
      {stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14]},
      {stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc273 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[3]}
   );
   gpc615_5 gpc274 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[4]}
   );
   gpc615_5 gpc275 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[5]}
   );
   gpc606_5 gpc276 (
      {stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6]}
   );
   gpc615_5 gpc277 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[4],stage3_14[4]}
   );
   gpc615_5 gpc278 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[5],stage3_14[5]}
   );
   gpc606_5 gpc279 (
      {stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[6]}
   );
   gpc1_1 gpc280 (
      {stage2_1[18]},
      {stage3_1[3]}
   );
   gpc1_1 gpc281 (
      {stage2_1[19]},
      {stage3_1[4]}
   );
   gpc1_1 gpc282 (
      {stage2_1[20]},
      {stage3_1[5]}
   );
   gpc1_1 gpc283 (
      {stage2_1[21]},
      {stage3_1[6]}
   );
   gpc1_1 gpc284 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc285 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc286 (
      {stage2_3[10]},
      {stage3_3[6]}
   );
   gpc1_1 gpc287 (
      {stage2_5[14]},
      {stage3_5[6]}
   );
   gpc1_1 gpc288 (
      {stage2_5[15]},
      {stage3_5[7]}
   );
   gpc1_1 gpc289 (
      {stage2_5[16]},
      {stage3_5[8]}
   );
   gpc1_1 gpc290 (
      {stage2_5[17]},
      {stage3_5[9]}
   );
   gpc1_1 gpc291 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc292 (
      {stage2_9[6]},
      {stage3_9[5]}
   );
   gpc1_1 gpc293 (
      {stage2_9[7]},
      {stage3_9[6]}
   );
   gpc1_1 gpc294 (
      {stage2_11[17]},
      {stage3_11[6]}
   );
   gpc1_1 gpc295 (
      {stage2_13[18]},
      {stage3_13[4]}
   );
   gpc1_1 gpc296 (
      {stage2_14[16]},
      {stage3_14[6]}
   );
   gpc1_1 gpc297 (
      {stage2_14[17]},
      {stage3_14[7]}
   );
   gpc1_1 gpc298 (
      {stage2_14[18]},
      {stage3_14[8]}
   );
   gpc1_1 gpc299 (
      {stage2_14[19]},
      {stage3_14[9]}
   );
   gpc1_1 gpc300 (
      {stage2_14[20]},
      {stage3_14[10]}
   );
   gpc1_1 gpc301 (
      {stage2_14[21]},
      {stage3_14[11]}
   );
   gpc1_1 gpc302 (
      {stage2_14[22]},
      {stage3_14[12]}
   );
   gpc1_1 gpc303 (
      {stage2_14[23]},
      {stage3_14[13]}
   );
   gpc1_1 gpc304 (
      {stage2_16[12]},
      {stage3_16[4]}
   );
   gpc1_1 gpc305 (
      {stage2_18[0]},
      {stage3_18[3]}
   );
   gpc1_1 gpc306 (
      {stage2_18[1]},
      {stage3_18[4]}
   );
   gpc1_1 gpc307 (
      {stage2_18[2]},
      {stage3_18[5]}
   );
   gpc1_1 gpc308 (
      {stage2_18[3]},
      {stage3_18[6]}
   );
   gpc1_1 gpc309 (
      {stage2_19[0]},
      {stage3_19[1]}
   );
   gpc1_1 gpc310 (
      {stage2_19[1]},
      {stage3_19[2]}
   );
   gpc606_5 gpc311 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc312 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], 1'b0},
      {stage3_3[6]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc207_4 gpc313 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[2]}
   );
   gpc615_5 gpc314 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2]}
   );
   gpc615_5 gpc315 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc606_5 gpc316 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc615_5 gpc317 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4]},
      {stage3_14[6]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc318 (
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[2]}
   );
   gpc1_1 gpc319 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc320 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc321 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc322 (
      {stage3_5[7]},
      {stage4_5[3]}
   );
   gpc1_1 gpc323 (
      {stage3_5[8]},
      {stage4_5[4]}
   );
   gpc1_1 gpc324 (
      {stage3_5[9]},
      {stage4_5[5]}
   );
   gpc1_1 gpc325 (
      {stage3_7[3]},
      {stage4_7[2]}
   );
   gpc1_1 gpc326 (
      {stage3_8[6]},
      {stage4_8[2]}
   );
   gpc1_1 gpc327 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc328 (
      {stage3_9[5]},
      {stage4_9[2]}
   );
   gpc1_1 gpc329 (
      {stage3_9[6]},
      {stage4_9[3]}
   );
   gpc1_1 gpc330 (
      {stage3_10[1]},
      {stage4_10[2]}
   );
   gpc1_1 gpc331 (
      {stage3_10[2]},
      {stage4_10[3]}
   );
   gpc1_1 gpc332 (
      {stage3_11[6]},
      {stage4_11[1]}
   );
   gpc1_1 gpc333 (
      {stage3_12[6]},
      {stage4_12[2]}
   );
   gpc1_1 gpc334 (
      {stage3_14[7]},
      {stage4_14[2]}
   );
   gpc1_1 gpc335 (
      {stage3_14[8]},
      {stage4_14[3]}
   );
   gpc1_1 gpc336 (
      {stage3_14[9]},
      {stage4_14[4]}
   );
   gpc1_1 gpc337 (
      {stage3_14[10]},
      {stage4_14[5]}
   );
   gpc1_1 gpc338 (
      {stage3_14[11]},
      {stage4_14[6]}
   );
   gpc1_1 gpc339 (
      {stage3_14[12]},
      {stage4_14[7]}
   );
   gpc1_1 gpc340 (
      {stage3_14[13]},
      {stage4_14[8]}
   );
   gpc1_1 gpc341 (
      {stage3_15[6]},
      {stage4_15[2]}
   );
   gpc1_1 gpc342 (
      {stage3_17[1]},
      {stage4_17[2]}
   );
   gpc1_1 gpc343 (
      {stage3_17[2]},
      {stage4_17[3]}
   );
   gpc1_1 gpc344 (
      {stage3_18[6]},
      {stage4_18[1]}
   );
   gpc1_1 gpc345 (
      {stage3_19[0]},
      {stage4_19[1]}
   );
   gpc1_1 gpc346 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc347 (
      {stage3_19[2]},
      {stage4_19[3]}
   );
   gpc1325_5 gpc348 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0], stage4_6[1]},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0]}
   );
   gpc1343_5 gpc349 (
      {stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc623_5 gpc350 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc1343_5 gpc351 (
      {stage4_14[6], stage4_14[7], stage4_14[8]},
      {stage4_15[0], stage4_15[1], stage4_15[2], 1'b0},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc352 (
      {stage4_17[1], stage4_17[2], stage4_17[3]},
      {stage4_18[0], stage4_18[1]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3]},
      {stage4_20[0]},
      {stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1]}
   );
   gpc1_1 gpc353 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc354 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc355 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc356 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc357 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc358 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc359 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc360 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc361 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc362 (
      {stage4_4[1]},
      {stage5_4[1]}
   );
   gpc1_1 gpc363 (
      {stage4_5[5]},
      {stage5_5[1]}
   );
   gpc1_1 gpc364 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc365 (
      {stage4_10[3]},
      {stage5_10[1]}
   );
   gpc1_1 gpc366 (
      {stage4_11[1]},
      {stage5_11[1]}
   );
   gpc1_1 gpc367 (
      {stage4_13[2]},
      {stage5_13[1]}
   );
endmodule
module rowadder2_1_22(input [21:0] src0, input [21:0] src1, output [22:0] dst0);
    wire [21:0] gene;
    wire [21:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[21:20]}),
        .S({2'h0, prop[21:20]})
    );
    assign dst0 = {carryout[21], out[21:0]};
endmodule


module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor2_1_64_16 compressor2_1_64_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h521534f7019ba947408991153a61ef2002dca621a3cd46109316c95fc81fdc8175d780eb3e2dca76c0ebd726e52f5e15a29412ed12e8bc0c233beb38a5c9cd587ac12e6ce6deb9a9dbe89f71eda2633a11ad9e69ee1b9c9949aef761bd641f6c8b6fe65b2b0f0f3277424fc2f5daf03546f26a7bf998e768f6a10baa94c2a855;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43c3c050fc49c83ca6db39af0e6a3d94e56a2327d9da2b8da0e31300ab71d283f468c4083094edd9e26308ad21f3db914ccee7241c2e8045577b60ca4edcccbd3bbde28e265ed69a0351c9d3d6e62cfae4696d9b20d36a91d9121b628571d6360e74584bac43719fcb37839a2b3b61ac8b98ba09c257ee9c59d9b43f9469e8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbe82e879dcf6919889a31c39b4954d07db66b8ca11afeefa82754c970052d59e28a8b32d01477eaaeb7b4a75e6311b694c4a2710717ae76ed96d21bcb677752aeaf0cd760bd131f00891fb120efc28ab053703985a9d81bc0bed7ddf5ae07e61c065ce1b4e946a4dd82c85a6da1d986bf250b1c8116b4e027d560c710310021;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80e598ea8d14326724ee253af83b595a94c16b1dce525f232dc95f0a8773dff54c61ca0f5460e33ed6d3c6d7349b2b6d735dfc66866b6ec20f7a91a6d4bcf90d3d84f3be923e876b565de224cbd50807dc67f2f4eeaf780857943ca8ecfc8e41867025d16813df0e6ee3b7e2224363bb7eac92c58082227585dea04376448964;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcef49129db3def436667b416917d72f50ea9884a96ce6d9b52b531f865c378f0e3d6d4c617ed07a23338d13e8432272a6054b70050abb4b20275f6b73be512068385b503111ccbbaaca35d584c18d2f16a59899cd0e8c4483311cf9c98fe25b48df1e12cfab4635edc2fde1f4059d163f45895a81a0fb3bd9c961d16f84ed294;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeb5ee490b45dba30f4ec91ba53f7998b5a07d07823a3b25a52eea2f94a7ea5691e5c4e7755c42d5ba546d119ff691ab42ef0d907b3d79dd1b12b619251842aadb5d27c2935de752e8102bbfea94b7d2cde40c7d1117c362f5176c5d89eb440d2e59b5ad907117866f68c462990691f750e40cbfd5c1c97b12674f332a759f67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fb30501a30b4c3aef5b897fd8f294dc22793c4a84a1594cb224a67238185675fe7dfc441ccf67f0600a9abf816bb484c0e40208ce9cca5beec508679aae70a3e5eb378d25573df0dfe97ab31513a98304ff51c7e2f5626fc9554794dd3d0a5fbe6785218586329de5705a6898b7a7e36b7ea8b6b9f5c8ab6454a9e5c0868b07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ec8bdc5ece3fceebfb7d8b690c747970d743e3b8b521253dff8c23fdc82d84f0e4706ef36ce08fdf75a23225db2733be014ce2b88bac89f2b77e2a3c6be63244c7f92b84fd36c2d4e88607f91b5c8da33c54a259b18fcfcbfd48726eca6642b5190c0dc1fcdbefab71cb4c94d33d3550b4cad0183a13e85dfffb3a6bf3ea1db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h413a331b1bb3820fb24fd893404ee9c1b5a9de3ebaa5f69e26f93834bf832249da2f24045bf4831e539636c9a422f94e33752d7dbdd8095b1fcad8da21c8af0d23d164f13fcdceb8e465c8153d0f6ea5eca6b23aba04d4da6a18216d65d6cc9f4161061e1a2729a56a4f4e2b929916a4514938879eb6c8984216deef53b0c1e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fabc2d85fbc4edbfcc510bfbddbb7fe4376d1cad72d749de198c1be2df253f4813bba5ba5bc2b27dd63e7ccd142325fabd0bc2290ef61cf1ae2b525a1ded45463278fef0c579909b18b6238c845a413d4d011e9bee107a74c4750beafa30e04bb885879857fb5801006302eb272e4af0d122506116bdce85cd8a3d860a11d76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5698dc6752aad4ff5ac2cfe9fb43e4b819c49d4abcd60ecb500c2f3e61b71f99820957375138fa60fcf71a4ef023c38ca2ce6310c3074172d1bbe1eff86e4843f78fb838de8225ae094eb364c1edfd5cafee6dee1217dd811e3daf9af92ab63f45783c60d3d9b6f377e2f0b9969ec6da2908ab4cbe41bdf6665eef804017ebdd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac02c22946fd13aa05c63f52030743f2a4656a9f503802b9b0ac4565f8405ad9d7d1494f0390e93ed455d764f4fcd58bb5b92d6a118224b9e1a6484b9c6f484d50cd332c175314f1311c88013b9a917c7dd06a933c60d7592b6e0101e4e062f3a9779e8224c34427864395c1cde8b18d839da0ce80f39dce79535a0816ace4b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h369d5ecae1d5bd00fc454006d7f9314cda8b4031390478d69b8933fb5d3fd2e213fafc9d3ebe4e82ac0cd5937bb98f67623441a69887b521e4faca4b2c5c41c79bc1db5711d4f1761d759402abd82be3a723a529795abef53aff7688b07c082e17437bc3696bda5eedd78f69c3301801d24b10f1f379ed1df48a127495ea361f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a0261c5e98b14a64aa76b02a276ceb61dfd89f87dede031cdefe9fa071ac931f2f87f99de0b0c1fa33909b85e97d633a88107a622720040a8c7e4ecf6f5c73da24d7556665e2449f44b79870aff9616b3f2e378d5f4ad1ebe8d6836b19cbe16b011aad02feb55ad5a8fc54567744c6f5ab7138186818df0aa7ff74214776fd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91837ddaa666ea0ba5305afeb5145f04345910c04e0926ce5ef7e887ce938abde38d8aceb06ccad0f4af1080ae837472c1451dfd0eedd89ec0078e539f302da70e0e69b49c45431838feb06496fb339881723031d5fcb5b71a11d1c632e536d7ffd2ed977cafe092f0e0a8837244b65be68e61240c273e4054fa77b7cef9f861;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc360fc2dc408ede4167923d83ef51188614864291f960affaeef0f2113f4c868a11c2effc71418eb6118b033854d2b704a3caf254d807be98b502e72c5bd6d86c8e3a4bc61eb09dd7a78447270a7d58c3a6e1c7afd04358b575c93d63ecff29eddbd9b4d3627b387ab91301263c3d95a77a0b2e856cd3727921a8d6225a608da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5759bd7ea114da58f9e62ab838ea6d36c529b4b8b7f42a81331d355ca8777d337e6f319ecd449b9a2a9c14d844df0639429b6caaa27e90221ae129ed73b7895909f82057bfa8c7368e562f0fba09660eba5b38375c3caa328639a26a41736862b104c8d48c5613921a46bf2fcfbf2e3231050c827bd63c1099697efe0aab27e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf7d3bcbf55a76594a4b79b6f37f4ad92292737d9456e0781243eec59fd9e036d602574a8b35babcb51d10a2f0a91260f60de977002084a821f5b7b7df771668ac3103970392663ff29d9a478f2f2ac036f8a3b958a61873d1e71a4a9b2ec8d169c069d4e03524f835d35af3ba9879cb691150743d26d7c978af331ede6b3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35876c790d35c34e1acf4db8a1d1b4a2833f06254338678f0cbe5393d1f47f31b20f341e1ccac7554c35e4dbb45f4d03e4af634ce8b2cdc3ca9bd24713fb79eb5cf84479bd372b92da6c410e3fa2861b5e74ffb98fc18ff7c67ae9219b262e2712a8c6a06a4cfeddf05cd60bec1a3fd7a96ac7b44e4ae6cd8aad508ed404025b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2edc290fb2a71b74d153cd6806f58877cbbc658ce17ecf5d34ce81daf6954ea1ed594f1db5e12070d22093cffd76519c9ed72fcf66a4c0fba90e2ddd17d74a47b5b4d3bce4580e842debbb0f130fb3fd539c24e89372bed655b758ff05aaf3f8bdd7a05574e4b2216f427aa49735433473eb01ac37109e8e4568a168bf8e3b89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f4e4563e86d30146aba06d1c833fec44b92df9d48cb0c2c760f37da1103a47813ce065646ebe354353debc39d87eb078082b090955e1bab58edf9870e005cb997d36f56fb4bc61bad7822affc97653b0a3021959ab7f5f51677bf773a7ff12d7437b4b9785d3a851001887ec30cc5754db6e64652a1d32410e13db9ad992290;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd61dfc9952b86bbfd158712a809d62ae9f0f5f70862af6fbb5b87f47df73cbf37a930516286b7d14ec5d5d780f9140f5c656afcf1fc2bc7720bd615a6e2c12a1e4ae68aa98e392fcfaf9e5fb43488e12dc1fab3c3089a1c58d350d44667e429cf2b2ff7bb3a2297e1cf6b841c9b1305aed9181d7187b3249a8e4cd297c9e6bdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8849e10dad41f78c36f336b178b15ec340e694cc2b12fb3f86102d195e13b0b18226332f6ad8e605fb26a0bb9e192ea973b8aa9d0c5af88b35c44a2d583a01ffd21ced60123e501be6622159c6473494241e2494b47855bb42324ec77b06f6442147ed5191016ce3a02b685a79390698a0d1843d568db021020cbaca50fae07d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b20ebc54cf86fe251bfbe9a351f2952ec9c7cba70e6ed91c6a22ad40975936bb0dd4480e2e6b2af1c452e6059420924767b57f9deb1a00cf83ac333de6a92b0428fdb9c7aebcebeb1b5b97c17e151ef3d3f65877f83441fdd9da8f09d929ea8a51a6223fb84ff47e34046e13352970beddc85468fc2e9e22e6c1336d4f905f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb000af4a33f687700d42cf83b725d833b374dea2962a48a993190622a235d7547acac031e50ea276da6314070b754fc5dee203926d05e2d1360263e3de78b45d25297bf2b37d4163430b51d8410e15460c5190c306ff5a1edce90d6eb8c5ed37dc523e067f2a94456c3b0b8bfde54650a3ae638cad655defe37f0a8f80429d13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde55d4f949b506ea0ed1a4241c17fcc10e47ffeaf62b2ce76ed7fc0b6e3b2e86eee146c9f7c54b6bb037e48901d2cab8ef43ee4fbf60787040b1a61eec38fc5e854ea74e46f6cfaf3c6bca724f61f52fe2d4ca3e8e4bc2d82cb927445fcf5c877c1dd218a3bd757811c28ef051aeadfc35fc64b263e4e949f6a7c9701286b72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ff7f4791dd871d91d26cb8e95e5bec7c32164f324f76cb533bd1a27380824010c352a1042f1ddc353dec7bd08470c2fff30151189ac7c4517f796cf136a4353350b8118408cb1efacf4926afe61f26796e57015ec931324fe77618e46bf000c1379d001067d99abe45bab92e4fd42785b3b34a5efc74fc1d552bfdcf5e814d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74d60cfdba92b91ff7cd85a991feefc840d5f6986c2a5e5057bc4c9d4f8e6665a1e10c97391b4fe203b7fe3aad581d8db69c3e5ca240aa5c88d68c777a3b4da09c038458dc17eda3ee2d67895d7ca5ffd7662a6a601d89c4dd2e0dd9f9cd286efc346cd2468c0b57c3d6b729004362e04abf4bf1431c85523f55f3e5f2af1839;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd0ac38e6e0de19139cb1484ba2b49130e6b41cc40eba2c511178a30f4b342e0e9350e53d8069df5d93ad3481f6e442ba0bc7319c8653cc4c95e42d367a7c292df48b5b9c373ddd0988bfa40b41765c30f43f98babd6e617fe2c606621865588c16caef978068a03ea432a2b55d874d396ce0837b665db4aa94da0e3b109e47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b16a4327f7aa62c15fc59417b1fc91ec689137ef11e2aa93193e1dee6661877b8ecd1fe0751fec4343169500d6b81c654c626ad954ca56e072383353f69b69ed9ef0f81071e4a2ca7b9833d956f828b76d5d026e3dd39c713e94104af728c2f763a703e455150e8e648836b13175203ba6a812e683c4d8ecd06c539639fa0cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdb19c376d57018edd957bc221b84aff3bf61590f8b2ead1fde23f7c752830c4760951b37e9b017910594f17fcb9c3bf5fb4b92052d9cd0c2853a52d99aa18041abb62c64fbb340f8ce7eed5af7b59b577aed8e77b3775952af33fb8d727e74cc5dba72d8fd388aa8ff13e719bee1799d308ea75f8c483accbe9a88da249fb2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf89dbac59a19c8460b722e9c77366ae99d1921b08ff25376f2096f237632dee1d53337131c399577a528535cc40d9d0706d186f766ae187144defa65341bc06e3c2cf7e74f669ddedd88dad8f0595f0e1c26665c63a185d93af4daf4d606c70c8ae3dcbad78d34bdba3b5d125f989654d0c0ac2a96b3e90695891215afa40c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1efa07b0aa54006d8a2463d9da9253445fe516d769f875940e9d90aad21ab8ba2fcb8b025cbf8322ff0cbaa4b727be4632acb43c5866acce9dd864acfbeb76d5d79657d63f1e70f7cc38d103c95d52c29ebbbf01332245240c9dde136c53fa4cd828ca2a235b0818dac8cdcec0ad98f83559a1724675338e0d7534ef4c4a1faa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53399ebbceb05aaee476563adfa7084d9d1d8ee86688d1de687e75de138c055e5fe62fd943b48c8c0b0a4e142743f422ca3d1011f3ed031cde3954dd27c4a197788c9caea4cb5e38eacdf7d94e6fe9037f7b7ebc6a21bd47da2bc4e14464cb0f224e6585d23a8812e39f4da5f014dde670bec845b40bda7718b0b22365438d84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72631accb60ba9a2c7b8863fab497d40018be51e2653363c025d99181dd30b6ea083e472f50cddf93ac8eac84a4cc506259185110baf6a41a3947018c55eb8f36a0a1981c2dabcc50151027c027e48ec4ca9ea267b5a729bca035102a17e3719e83d2ba4714672627c25fe77787529e4d806933f7e4d7497f5e696f097a3f45;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f31a7db50dcaa2a8c57837815e259ef8ee9c6d1e1d9b61c39c8461f4032144a8606d111fa2847d38c02d301bdf871adf5ec66df67f3ac016611c3e3aaec22f73c43ccb828e66eec9886c3656ca2779646e5a62228f87049fd896db4b2842c1bb1383b39b7ffe1bc6ed4fadb4ee419db55415ab99ab10ff7fd1f357cc896b3a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73a63c39b324a6921503425f7746c73cba16c569e969f2ff3af19630840f858923f55e14c19a8aeb8bfe5487cdcc2e6470e71630a7bf5ed53e0dc7dd89f966e0dba42e55a4d7d8adec471ddf64a96d70691b943017ac4a1f019d30356852545447b551d6635e904bdf031ee5ae92e72790baecdd9d0554682a26cb053d8e4fb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h656ffc616ac29e1057464b4a496f93b9b62ca237d06435ba82934abd7097d3cb13fdc960054adb089947ac45601edd3cbbb590cc0b524f4a06fdc95dbaa2edc0b2fb8ba29665ee32e88f8bca229122cafe135fadd73b286fcfc7e057237e6a9e11bc7e717256e72608c71856eb7431bca14e35d484d9e7b6d45cd0221c59848f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd086185954b8862c534a15e73ce59c698222dc7a68036bb8fa83576d0517adae6d51fbd917fc5ca86b0fa5b865acbf347197100b5958ba167ba08c0e774b7687d5f39ac97b8cabbd7ace36bcc4699619dcc7138de8bcfeed330a3a50f391d4ba6169d7a5d097495d339051f1ec02055680da47a54934f9055d80aa967f2197a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20ec22d9c4848da8a5cbb8cab89396c3ebdda9db51943ade89477fbca38856a3cedcf8b3ca11437edbe2ae6f001033596714fd68039cf2e1ae652eee3630f41cdf793b7b4fd60d3ec621e1a4cd6c41bfb33e06644abd28846176e0e5bef624436cf0a821edb2661832bc85961b38a7641420ee8cfd2f40fd4356a8fe7721bd26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf98d3415821c2be8953272526572f3177f30d5433b0ba9c9824f81debaa9bff287a4b7c322382d7e80ffd0c0e439245b1b20e86f57793e0ed0cdf6632caeb7c4b40eed66fe1ab3817b30b8aba5cc26cdb971207a54c8681ef2ee62d14ddb4897410f3765683676bea0dc19191802dd30e0104121e368d9c49aa9ee52b845645d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d084655eea07ee3872b67135cde5f333e43c9cfe199e89564ade57e53c1f95055e7f29fc6f786a663dabbc62ab953c5f17242b5066f60b03430f1651251352c99277dca589ab02adae826d384d98d472cab6c99d271db9d28b14ccda52b01d02275622eedf654c5cb151ac8831a7790d798109583e78c863a808b78f7ecd5ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h507945b368cc4af7e11e53d81ba916aed834b04452db4dd888065d5cbd46e2fc3d0ada7c9629ddeb54148a9ec07bc63ba8f6316d36993f977c8343413ab1bf264340d9848e5eac13ba3fd5bf9b7ac2bd59bee9a19bfe6fa349df5ee656ecbcc3926b2e8086777d6c5ca9660b4d8b5eb770860f45dff59137ed12d733c444e3d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34455f3f604816ce482da8a93522642f69bc8c7aa3a3b9da4cad12d0847843203c92c69b8e5f6b1f9eff72cf011bc20aab265548f04d9fcb94bbd6e06d45324b787c3fce39b18807a5374ae2616cbe1772dafd4b4af73710787225e6f2474cfb8eddf6f9e7b30c6274225a9b10ac9bd62bd0b10452f2e8942f3fb98f6d1b82a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc155d643c1aff818fa47b1c5a231c5cdcc8d06273ece507db8b2c5ccf91efcf0384bae761dd08c4b8d5b12d709f8de4f28818f2834f06b09cf5aa7ca574d027a9efa8df3287bad42bea00cff875588be5ce7580d18d898db907208ea0206e4bc4815faa2b509be0c50279e36fc5fed0cb3bab5c54ec45cb3f7f002195a0e17cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21f9bbe7b226681488cbcd103b444cc44d7b1d3458a3c6994f0cca012020ec7f7c2752a34af5a27c1bd2639ca3cf8a702fab9dee2371374535dc36e7bd7ef0cfcd23f10c1507adb219c76869e66c1acb059aceafef0cebe7566b5cc4199d424f2a72f52a3ff36d607fc7e4b841e16cfe5d604fd52b5258de9d5ddd50c403b37b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb1226b1840292074d89213b6806be94f77090a72a7696f35e11f1c89f9f0fb6518d8335345e690bd9a099cc0145bfdddff07ccc683879b6399ae86e1a4c2a15f6486af723d11d907b074cf31471f2632c0c3882dac5a06683fc90c52ac40e171a5b1bc33bd1c234955bb61b42fb042c7c4912016611489d66d3910c8c62ace9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8255e258fad5555268bc9ff92d57dd1a53aab05147eccae5718d29d222d1979419c7d56d027aed427a46ff8a107322b18188b3d044ca8c09f1473855ca92fe0ef0b93d68271239d8c9b54d6789405472960c4170b41039a1f2b135af2db5e5666c255aeebde2e2d85cf1b6566b9bb9907142bc517050473ac95dbd060be9fb52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0ac2ee463a1d85e1cf9a30ddd1026294189f4afc7d509bfbaf8b83b9b1b92a94e20eb2c254d5be9e701283adf5110e550d8a7e208ad77037596fb4a5ec7119a266b39bc308f1718d7f52c8ea85a1e5858dfce40cfd83937092eb16fa5eede76d6eecee630c12f32d25e01b866dfb027951e04dc4c0879316f3ba05f08a0fba6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd19b195cdb6270a9c6fe7ce79714e9ab21587094eac7e0df51e9115d7434ec21a28ad8d938fcdc74d30dcd568c9d852b5a430cb6b0754c809f40d24e84d5927ec3c22b04df6a6d89f3e184e56b52ea79e8e180cd90a27c167944d6269b2bffb598739c240d15ac622e220a96c25ec38fe520fd707e79a83ec28170c41c2e5d75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a7ac16ca1620e418d41b2c7e782d577a6b99ebd3c5183d456f865b9400d8b3f9ede380f74d1423369bff3e3552f63bd99c6093be86086c9263acb644f47c55a843e18745cf02feb604c4139877e3d785734856a0e251d29f1dfbb6a5140f51da263b49c055d1b2dd2e9898deed9a0413dad20e20f5de0794414d766a05d4c96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h353e94221b076d7f411fff7aa2d4aabe8950bc4885d3919d6f15972dc6301c87dcc9b15fa240eca9ce165daa44b41cd1210137851fb569eeddf1e027b3a1de99e90c2ca8068a43122a9cebb334341d5f3334cb8ac14415580a246c40a65bc956a14e9edd6f86607d5ffe0bbd85e8256805e58c0c5d5d2fa0d5e35b78d1c5c4dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d9668c59f37400ca6f6567ef3c8892bec7bc0a851cc942beca4c79988e855cc703ef502e40db9cd70c0316ce0f24b06cd606ce2ebb8c911502bf76d2361c933c4b65d9d497eb9e7946cff69282493a645e80a498a072bd2a6d0aed06270e3f915dd9387454ac81ecf6c97eef6aeb5640c473bb2125e7308cd5309d63bcd6f0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6977ec9fedb76580d4c7199385cb81a22eaa51a5fb73f39b134f76c43c09de87987d564fc7be019be5573b5ee326bbf0513068e9391e1a402549ab77e3e8a552e49946351f889f5f404311cb6a064f4ee4f35fd536deef7bc930a34dd96cb12257176745a21521d018bb8f5b633954a128a41bfa95d7d3a0d349cd2d3912d05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37cef7d88974d92bcbea4dc3a6a5317514fc60c0c4cc504ceb69c8938dbbeb4a5b27f1be440a2f749e2d3ecd8ad6492bbf7311f22411c626c3e376906825b8cd4d37c369cdeb886b51074d5e567b7854f9ead5acfbb8794db49c263653f774b17e294792f0150529beae16f307fd72940c127e2ecd49083bc8f46b8e435aa944;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b243dfb1ff2bd30730dc2be172035b5064fc913305c7d21206ed33480ca99e57e85ddd7081c757acc1b9110f5c3883dd7db6cc18f4bb7d7a74c9c384093c7b532852184dc72735614fa9bd768d29a2511b7fcf4b862ccd4e13ef37aa2bb0527c12d62314951067d6d2337d8353ea4a2e46b936bf20369ba1f52dac49582768;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2ffc05333230f77955ba90f3ed8f68b19da2bd514454ad29ca4adea0ce59b79431b69e47c98c291187aa64df656a79e9f1a281a948dd82991ab5813194ca9c010acee41734f9847dfcbfbe8f5ed035f2bbb36425fdb3d3b99450af89239d7d2ac86f4906c1612e1836b77918050ac04765b6986be0922e5c9a80461fdd4c40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2241e11c577057b9c78acf3fae75e3996c1505eb1799ae6357e7f5a62285024ac5d54b10994747cf48f8628bf18a183ee1fe7c5d021da261932dfea11dacc1ff479a8c4c5ddbb05a3c7f7e6045541eee428f5996e2b7524fb7fd230cba170c3d0a2617c5eb17c77d550fe16a73f779cc245792ac61a04f05f4582f92a77d0662;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e1a33e5dc285bf3c72b7acd8fa8ba34713b724df1c299adbed0bf5ce01e54edd0fbc7035b3e161474de108e63821268ef4e891177561475ad926309933d3ba38f14d41f3b953cb111e9c81399bdfd60bc5461c7cff4b378911b021780cf8fb7e63d19585d44ee6f2091c975162e2e39b81aa81dcdc5ac7de60cdc68611b2cbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb81b5f6de16934e9740d8a122d2b6ce6d876ca4ed7056e74df5924930d293c56b68c29a0986fa0efdde5be529ba81fd7c4b57485f88a25f36f82839f766744a3966fd07cc66072104dd8d7a798d907966cdd8c90908a1fdd069da9db9ce1fba4828f2fe29cd400e0594196cf0946ac33e0a7d7fc42ac78280e05a4c2080db98a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95d37570bd9bffbdfcf7845ac7f8e49caee325e7c31f287ec28375c9bcd4e5e692b67b3d06a631ecfa979b105a3966291b8f3f35c7672b23539fda7493d7cf4294360c33afad39e36439e34063766bc93815ef4d2680901c8899eae9d24f83a0b38eb15205a3dd1d5daac37f2be66f6f32fdf1614addd1551de5477989721379;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h560442664e3e12f12f23af8906286d69cbe287d1d27e12c60596d7ddcd6f99353d169aa7ce1c5c4fe9c34bb6cb7e9f622a4d4301f48115ddfb55f96ee094a1571d0089c46da04c7045a720f98758ddb49082505cd9d2e845fae724d10184aaf507da3754655e93510dd8b9bd3621128cf6d31c93ddef283011746b760b7a3c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87fd90dff6a51ffb897a2b7818e8ad36e243c7c7a8595e29fa0f510173310541b125ca60a12d5fbe7488f8ce22db0afd3dbedac4d15062f15ada2b6a5049e704521a1e0efcab6d3284944f7b744b213f87697d26e8c522a0b2d1235490b231eaa1a1be2df558b550a28e563ce98e052c8a872b215e96fc20383d551ee3f4d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7d716c48a8cf80e5d5e5d1d0d258ea985a6eea6a5f8114779ee29cea1c715356dcbcf5961af546921892518e9767ed3157606482556c6f6df678261a6a03e4ef148ea2e45595119a0dfc7eeb3c65c1850dfaa010187a14911fb35c473dee7c0181294dc3fe7ee110acd2389bb56e3d3a6372ac7f91ac9e827301707b9f6bea7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he40061233eb12b03fd9c48e7b19232ea8d065de1043105ad8c1a24df9ecda65e5109785ed116103f468c38d7a96912695a76879462c9d95cc8c9cb5bfcadb6e87955e47f0a144696c2c2b148937c160e5964284d1a2c411095831f50a3ae243272367f87911a3769d6c92ffb67343bd36eb9f7994ffebfd9de656665b3a619df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6da82b8c1ea1a3c9e47a4510c48c0f332f654c2c35059e6685f84d961079c3f70e9defa00a8a544a8fbac8694d23c563111bb16f6696e2dd5f714155efa3e3f84e3df413914e5a207c75270f7c286eeb6464edf1e4fe62d782bad5db0d50641855bef8cfcaa75c39bd61c7fbdf819964756c7bfd8828b7cab8a53b9eb0e1abc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha66a9a338e23bf0751466d4be0a42bd3ec9c8ceaab702b3b4fdb50f89a32dca8326f5ac68c5c87a18c07a96f25ea2b6c9786373df0a6838d87a6b7be85547c58b4f40b2d239329d299e50387572049d11d081388409bd190282a39525e14313596ec5556343a67e34f45a36f089be9644e3bf83fd553f9148af060752b1a963e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h823463fb5d26175e227c99d4c1bfcb38dd89ae7741a1dee5cd25e890432a3f0cf1233159b10676db04d897eb5feba783257fe7569ca434e6d7424ea6d8eb4672a924c077f32e856019b5b3d83bafe837da08950b3dafdbb878fb51cba0bfa948065636374a7415ef3065ffc1fd5d956c85112f95cf2fe710b4bf3399f14a2eb6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97d010a36f103f71cf8e7707110d6d037f58aa9ff2dd4a94b5143203a9387a18411eb29f6a8232a4d8b8771ee743d0a0ffb3c9e5a55a15c0dc9655773d74da1d14ff63dce5a37536d986cf7e1b3a88d90f23ed50675f239e8306d9d73f95e6245c74698e24eb0a73caec4c8a51e4ff32a2cbad169c0e2791de5883becac0d3a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3607cd4c9c160b9a6b5ab5d816fb947d4b538dcdcd6e38231f62fd47da92a730e3b160a23e35a9402b14c44d35311e84a0492f102f49a285f929224a52681e875092fbd533b5da7c8e61c62bc846695fad715afc8ca0f4eb2ca1f2ff22131d931771ebd474ded2b4c8314d0e9ef9560325bcd1f886211862a62fcc432a648f18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h665f387f828ff8c4b7f60f41c056d34353fd677c15dc7fb1f32664add745eb26e994b15303ba669e3d36d6443974068a58184c3b592af50c6508c60c7bf25e1cfbe90bc8d045ef6af3ae0d242d96cce88e95bb728bba4461cc04598e7fadaf11942dc77e4a8164ef9f8108170bf4e7cb3a7112bb355bfdb6fbf74fa3dc694fda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heffac50a154a2a76ba43d7fc2fe3bc52cf7323ae98749ab9a61eb5536b6943a393478b31f0f47c6a70fbf0c23487f5fe682476ef8c6435f076260310f3e5ea786144898ce301a5a213cdf05951286b4da60d0c3d9a3424cba8e82c6b7730773ecf3ee7c6ddddb61969a76f12aef8475e2a134517fa040da5eb57a7af31a2e7a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he55a23d3e3f49c69dc5db53591e98af8ede5df2520d495f5ca2fa820aa7305af1acc7ac43d1be12b34a7746578fa4008d2b4ae36a6affcae2309d93e916b3455dd6f54930f3885887c0eb5df07d6acd2df9c7b61de5070e2ab986cf93f82a1d31df9a44522cb47e5cda83ee04984c264387348315da5501ec9844437a3a17e56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c22f5dad53110590aca8974325613e6b7349c22e1d62fc4f575182cab3e94c913f00c505a8226f5d5e4fe293fd5d4a245ee12a2fea60a1bd7e3b3b2fe97487b78f8b80c3df953c268ecf6b9f800876d5046b37e65fd1a0741987f9bd27f8114b991d7b528d05e5913ecd4b34a9d7e02fd5d0a2ef6799b5f9c26f090092ef7ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee2196c7658ffdf9bbdea264febfc159fe8aecbef6344a857c76ecf381fa0b7826aec371b07288f273ab83a3ab7d6e749a11c14eb6cf33374de11e3c70c9717faf85af948036b712e4fdae7370039e1ca01fc2075bdcf4f14e8091426181b54114c770785b53283c0ad81b0d3bda44658f0c5eb5623357cffba555b1262edeb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4ee84e1472cc546d5b553a1948466e7091b18e5906d5b6383d202e7f821df4b3dbd71ae6c0044742b30ca24723a1dacc23ab108c0886049196a26ccfabe3417e9456623fd40203e2363f7f9d1dabb44ad5c1e43bcb6095b478a89e3d61f1db67b16d1ae06f28be7ee24aab91a037a086fde0a19946f2710f0c574acff328866;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54e06f7f7989ff264ede3b058cd14a28fe2ead4c6971ff7be9644732517ff8d2b458c3849be3888178d741d08b391db314b315ca6ef32b5a1bcdd091ee07dcbd5ea5729a183a3e9d931fc07a2f8350ee8c81a1a3241cd396b4d56e2351639490d6d4b4e47260c9e21df5e442fef3033e3b3b410e51ecc2741f926f4305ae0547;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ed0d8f6c2ff51c71df1d5c21da96bda7db343050af420e1b498b7b26395ab7bd50298d96f053575af10a0a5e6b9ea2bf7ba9fda7b697812232bd0c774427516c6e2c03a6e8371064ae844b7b77db59518cd7cb7dcf04f2b6106e45d3bfbf0c5ce870971f7dce4d00310fe44aecabc91534d969e17e61c106b0d2930b3044685;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6df9e1d4068ab6edaf7dcbad2128df51c49c933b37a3b931811a3c86ebb9d9f3f7047737543798b16a8c409f3224d8db0a24924d2dc98ac5d605cf0b2ec0534bf9c0a091fe1af8057739048b61eaba40ce11a842ef47f2c76649e172744b52f60f87c11df9d64be81a3fda07b50ea2f76a3c5ebec7c5d7806862b9cfeaab12f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8422fd04d09d8184b4c4edfc7c8975f58ba2d43d9a7043f5dd75cd3c0f6958f5672fe0a2edca86636cbe336fb76ec349a9621b87d1ba6ae4f46304b163a110ed45f2aee7bdfd59f4c743e024a91161bf5e28afbd621be1730f7cffa3a81ff31573538c840508ab0a6dd663c14b42a628b1f026f125d5098372ac22a5a6233dbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2d54ec7577282764b1a09f5bc8f9141b0940dc298cdd55d77067d0b6396f8e0fff8854eafd8ff9b4093198c81dfc202bd2214086eeb25e56bf3be8d60c570cb13d3763bd49ed12e8a07065d956c9fa7dd57a34f0fde94e3333cceb5feae1b1ab0c72fc907dad49aca34fe50200278090f1f731b5ccc9457351ba0fae899008f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32a049947877e224ab53b24a0089480feddec837381818349c20e96e2090461cf7eb53f44e1bda7338da847e31ed91f5e2bc4384e523d98a784fad9d5b1be7d8b13112bca3001083e13da0f56d26da885afd26d9a37e10da25703f3f34fa7f6ef560401fa512fa215f10385ee9c4bf93bb0fa94e71e9c27f97b6bd28e7be32c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2762e021c2b1688092525ecd7086841bd25163474b7ec15d12d3a24568040927b876e1cf303f633ee93987001981c545ae432813c7651e56cc7a405d03c12c667428e4f8057b25eb9090104b7466b799d5d0e0332b0fb14bab8c1cddf220b756cdf69e96ef092d68c5148fbaf1376f1505978d71744d83892727abebac4afe9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h901f70024148890b8f7b3f68d8948e84fad11bab6e5cb84654beb53d28c3888d07924968f4a2b085fcff2580b802cb28933ee60a36c4c353d9399451662aa7af635d709abac9836c2bea4d97dda20c0dc7bd6c4ad881ea1183b6dd5a520fc84dc03aaefce3834ab4f592757127df247f133c11b1c0ea630de4037901f3d2cb3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1cd10ef54d32ddba5f4c148138c674825becc7a93eeb0d596337c36c3174c5c3c640270ddc7bf9b3df46fc05ca8a32ca161c3053430b296d5fc83337e8682086ff576918ba867be30087fd1c43d4b5a37b355108ae73db63ecf6480eec84540ad7d9f0c97de172970b372ee21549234d82cff17105ea3462f36870d6c194a86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h318c011fb52f5d33bdbeee1c3224a5673787d5a9d2a83086ac0c865272ac607957a6ad3f3553b4ede15a1ad3bac33ef5010f2d06778757da9135c4a2ef6a83b5469ea813ce9cc8b5f2875efaa63bc07cbf7178e714b3e637cfd0f724e5e7c3c042131724a1cca232f7dfc4b7d5c64d68fc69f91544784b54e6b241249ea6b646;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34f6fec4282a37099af6f3085cfca940de8ac561adfd612adb333223161fd523076d3404c8819b2bfff4c11bf0892b8df5edb3157138b53fbfdb2e03e6bf0ca763ecf6169b757b848115bd7c22b924a0a85749de9cfaa401d26e1485f0c31e360f669e44c9a0aa51d4fc511d0ab0547ad4271669bd9df327c6462fd05acb6cab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h963957c93f7588d7186924f6c02143173f17a91f758acbc97dfe0d44afd56a7716b619a2745e11648f82913b92cf1f52998457031470cc91d603d7ab4901205b7e4c7a5f4909f68394731a0c71c2015e3527b763c2ee00e1bff7efa6d9151c284f75e717e73ea512d448562cd403ab6914a4a38178a50c5d1187dbb5d963cb8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66be8c9d4ed9ba5cef250acb1e119dc46ec7398c7db6d7529570eaa0bd542649b42457aa48e3d68bc100df96804c7c75a0e414749c71b3888c316cdb93012134ef517b5c43b580fd870bc1a52560c696d401d888d9e2fa03a727863e5ff5b5412ddaab854f2f5f0a4e94447923370eb063a1b5d0aea131bcdc379b96bbefe75d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d12c1612bc83200b27bf8cbe12f17f2e7ad340b2904851797e3dd7b2b4b7938dde4bb3f58f5dc3df533ae7dc4c20c65244ba93feed729d23f9cd835fead5147a19ba90839b11c05757520772274804fb77cc35b1341dcc3e008a7bbf3bd5dc9a722c29081e76269d161e1b198fed73d73ca1265db0d16457f4a28d67dde4db4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94319e7d75e598e7e8197e1335514760161c4ba7676a900b64dcd3fa89abe799e937aad6d039be8a8fa9f4a54f297faeb9bb0c0207a6eeb0de7fbe1d96a5bd8b33285d6a446d20fe19195653ad5bc21c19f41a39b596cb6d9c7f51c84b739f4cbc3f02dd591b5616840c1db372e8e669e113bc354d897eaff1b7009e00466369;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1575dad2b19d486d499aafedcc123730fc5ec53378e5f079ae982aa519093a21b461bba898b81cdf386ea1903861ac5394f156d4eac75cc5f1a601f54eba62605389b5e4a4b80b3473ec1383f8726ffd91031d9a1dc810f9c1b40a095d7e0818998784f7b67042e2f29dfeb7f794939fc36530735373746590aefc2f620de827;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dc9917e886e9d9b41e9a19f42668760f5a027c5bb57c49c07fbd1a57450949ee41fd25331e70afad3bdb3ffe8bf3d8976cbf8540c032abad9a752bdb325435858e089c17ebc38b7d5b8d0649d9d86ec9bb732d288763202750a8695d27fac15f2ec1d6c04b130a056954fc1649f47b6be0da45e43f806c8789aa81f5afe54a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dd6dba7546c974471dfcdd7477db82c925b29752bba0f14c9c03cb7154e91a21e20eb96a9eb11b0f62e7bff365f1864629231dc9235c27d8e70c10ebbd7c470eba2519011ddd025f750789c449b7cee4d684972a762c254f0251249af77a85b0dd52c5bdf8a2d64c83ea2c73c14a874c3a0575f08fd5c1a653a2090b8f01ce4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13cb201088b0af21ac24d0c89bcdf95c4b619f58a6de77eda7375acd9b2535fb7d015a36d7893fa34b5cc460208532610b4b11381a724e8dddfbbb7473f101aab0d0062a08be036ff86316274487b4dbf3137979df6e1c7389e749c7f6d460e7831ed6e690e8a23564098ea2ad61b08edc7996a54007bd9838f8538bfd25ce7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55650d8efc977dbe3567c1171ff02930549f2ddc026d1b275e456f442c2fb1854f4e2013530af59db5cbdfc10b6081bb1f13857b85c0b76f132646922f4fb51794d727316206b8e6176488baecfce410c7309fef1d1bcc1e04a8b484ed4612a3a743fab2835c70cc0ceece847f1276529bc239bef4faac9b49c8e4b63d6d9ccf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70966969621ccb70618c66bed022da4a38530e98393ab672c175bcaa719038b7a6dceb611f288833b118a52e8c362de792563db24029a1e4b0bf626e742da9d032a1adafb8acb8d47f60b295632621bc8a3ab4448f93c9cd34679b44d9e20fe6be02ebec6771c2b57d81b16851eac59275dc112d24dab31ee1da6ae086ae3023;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e468c85585d0118f4ab39fe1398ec63d4f4c8458307eb4416ed83e38311e38b74ffff34b1205fbb40157ada3741192f32e76eec352571236463aa25ebdf7b6f4d5d4da373b1aa5eb830714614938b14b4f5627248a31f8646231007cdb35390f9ef94048b2ae3e25d9859e9701bccf39eb3393099a9f2eca2da6a44bb014bf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c9f7ad9e1e2e46922e7b5a2cf0f1b1ce444ceb912437f2f503f022fefbccc452ed14032f7ea6548d8f34b3ba42aa4ce640773535b7469fe6e20135dd2803b4eec3e99f8f802b6007fb2374a533f2ceb76b3102c2e0988fdb3db65398c248e4f2e9d74290a41e2d82c1e2411f4d852b1c7840fa21e4e304681538e950aaad79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f51bc255d53937338ccc2e5105ecaac8f51952472ea8347a32673928eae06e019067c774814af8a9f977d3121f87b3290fbb2af36ce164e89772b67b8f9831f682f98bcf37671ac8ba097db1360e3b4cb13fc335a7bfe230041977ab0c9583655b4f568e21652fd845b5011087d4340794adbdb51bf012b54f5ecb6cb89441e;
        #1
        $finish();
    end
endmodule
