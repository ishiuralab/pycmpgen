module compressor2_1_185_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, input in_data128, input in_data129, input in_data130, input in_data131, input in_data132, input in_data133, input in_data134, input in_data135, input in_data136, input in_data137, input in_data138, input in_data139, input in_data140, input in_data141, input in_data142, input in_data143, input in_data144, input in_data145, input in_data146, input in_data147, input in_data148, input in_data149, input in_data150, input in_data151, input in_data152, input in_data153, input in_data154, input in_data155, input in_data156, input in_data157, input in_data158, input in_data159, input in_data160, input in_data161, input in_data162, input in_data163, input in_data164, input in_data165, input in_data166, input in_data167, input in_data168, input in_data169, input in_data170, input in_data171, input in_data172, input in_data173, input in_data174, input in_data175, input in_data176, input in_data177, input in_data178, input in_data179, input in_data180, input in_data181, input in_data182, input in_data183, input in_data184, output [23:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    reg [15:0] src128;
    reg [15:0] src129;
    reg [15:0] src130;
    reg [15:0] src131;
    reg [15:0] src132;
    reg [15:0] src133;
    reg [15:0] src134;
    reg [15:0] src135;
    reg [15:0] src136;
    reg [15:0] src137;
    reg [15:0] src138;
    reg [15:0] src139;
    reg [15:0] src140;
    reg [15:0] src141;
    reg [15:0] src142;
    reg [15:0] src143;
    reg [15:0] src144;
    reg [15:0] src145;
    reg [15:0] src146;
    reg [15:0] src147;
    reg [15:0] src148;
    reg [15:0] src149;
    reg [15:0] src150;
    reg [15:0] src151;
    reg [15:0] src152;
    reg [15:0] src153;
    reg [15:0] src154;
    reg [15:0] src155;
    reg [15:0] src156;
    reg [15:0] src157;
    reg [15:0] src158;
    reg [15:0] src159;
    reg [15:0] src160;
    reg [15:0] src161;
    reg [15:0] src162;
    reg [15:0] src163;
    reg [15:0] src164;
    reg [15:0] src165;
    reg [15:0] src166;
    reg [15:0] src167;
    reg [15:0] src168;
    reg [15:0] src169;
    reg [15:0] src170;
    reg [15:0] src171;
    reg [15:0] src172;
    reg [15:0] src173;
    reg [15:0] src174;
    reg [15:0] src175;
    reg [15:0] src176;
    reg [15:0] src177;
    reg [15:0] src178;
    reg [15:0] src179;
    reg [15:0] src180;
    reg [15:0] src181;
    reg [15:0] src182;
    reg [15:0] src183;
    reg [15:0] src184;
    compressor2_1_185_16 compressor2_1_185_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .src128(src128), .src129(src129), .src130(src130), .src131(src131), .src132(src132), .src133(src133), .src134(src134), .src135(src135), .src136(src136), .src137(src137), .src138(src138), .src139(src139), .src140(src140), .src141(src141), .src142(src142), .src143(src143), .src144(src144), .src145(src145), .src146(src146), .src147(src147), .src148(src148), .src149(src149), .src150(src150), .src151(src151), .src152(src152), .src153(src153), .src154(src154), .src155(src155), .src156(src156), .src157(src157), .src158(src158), .src159(src159), .src160(src160), .src161(src161), .src162(src162), .src163(src163), .src164(src164), .src165(src165), .src166(src166), .src167(src167), .src168(src168), .src169(src169), .src170(src170), .src171(src171), .src172(src172), .src173(src173), .src174(src174), .src175(src175), .src176(src176), .src177(src177), .src178(src178), .src179(src179), .src180(src180), .src181(src181), .src182(src182), .src183(src183), .src184(src184), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
        src128 <= 0;
        src129 <= 0;
        src130 <= 0;
        src131 <= 0;
        src132 <= 0;
        src133 <= 0;
        src134 <= 0;
        src135 <= 0;
        src136 <= 0;
        src137 <= 0;
        src138 <= 0;
        src139 <= 0;
        src140 <= 0;
        src141 <= 0;
        src142 <= 0;
        src143 <= 0;
        src144 <= 0;
        src145 <= 0;
        src146 <= 0;
        src147 <= 0;
        src148 <= 0;
        src149 <= 0;
        src150 <= 0;
        src151 <= 0;
        src152 <= 0;
        src153 <= 0;
        src154 <= 0;
        src155 <= 0;
        src156 <= 0;
        src157 <= 0;
        src158 <= 0;
        src159 <= 0;
        src160 <= 0;
        src161 <= 0;
        src162 <= 0;
        src163 <= 0;
        src164 <= 0;
        src165 <= 0;
        src166 <= 0;
        src167 <= 0;
        src168 <= 0;
        src169 <= 0;
        src170 <= 0;
        src171 <= 0;
        src172 <= 0;
        src173 <= 0;
        src174 <= 0;
        src175 <= 0;
        src176 <= 0;
        src177 <= 0;
        src178 <= 0;
        src179 <= 0;
        src180 <= 0;
        src181 <= 0;
        src182 <= 0;
        src183 <= 0;
        src184 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
        src32 <= {src32[14:0], in_data32};
        src33 <= {src33[14:0], in_data33};
        src34 <= {src34[14:0], in_data34};
        src35 <= {src35[14:0], in_data35};
        src36 <= {src36[14:0], in_data36};
        src37 <= {src37[14:0], in_data37};
        src38 <= {src38[14:0], in_data38};
        src39 <= {src39[14:0], in_data39};
        src40 <= {src40[14:0], in_data40};
        src41 <= {src41[14:0], in_data41};
        src42 <= {src42[14:0], in_data42};
        src43 <= {src43[14:0], in_data43};
        src44 <= {src44[14:0], in_data44};
        src45 <= {src45[14:0], in_data45};
        src46 <= {src46[14:0], in_data46};
        src47 <= {src47[14:0], in_data47};
        src48 <= {src48[14:0], in_data48};
        src49 <= {src49[14:0], in_data49};
        src50 <= {src50[14:0], in_data50};
        src51 <= {src51[14:0], in_data51};
        src52 <= {src52[14:0], in_data52};
        src53 <= {src53[14:0], in_data53};
        src54 <= {src54[14:0], in_data54};
        src55 <= {src55[14:0], in_data55};
        src56 <= {src56[14:0], in_data56};
        src57 <= {src57[14:0], in_data57};
        src58 <= {src58[14:0], in_data58};
        src59 <= {src59[14:0], in_data59};
        src60 <= {src60[14:0], in_data60};
        src61 <= {src61[14:0], in_data61};
        src62 <= {src62[14:0], in_data62};
        src63 <= {src63[14:0], in_data63};
        src64 <= {src64[14:0], in_data64};
        src65 <= {src65[14:0], in_data65};
        src66 <= {src66[14:0], in_data66};
        src67 <= {src67[14:0], in_data67};
        src68 <= {src68[14:0], in_data68};
        src69 <= {src69[14:0], in_data69};
        src70 <= {src70[14:0], in_data70};
        src71 <= {src71[14:0], in_data71};
        src72 <= {src72[14:0], in_data72};
        src73 <= {src73[14:0], in_data73};
        src74 <= {src74[14:0], in_data74};
        src75 <= {src75[14:0], in_data75};
        src76 <= {src76[14:0], in_data76};
        src77 <= {src77[14:0], in_data77};
        src78 <= {src78[14:0], in_data78};
        src79 <= {src79[14:0], in_data79};
        src80 <= {src80[14:0], in_data80};
        src81 <= {src81[14:0], in_data81};
        src82 <= {src82[14:0], in_data82};
        src83 <= {src83[14:0], in_data83};
        src84 <= {src84[14:0], in_data84};
        src85 <= {src85[14:0], in_data85};
        src86 <= {src86[14:0], in_data86};
        src87 <= {src87[14:0], in_data87};
        src88 <= {src88[14:0], in_data88};
        src89 <= {src89[14:0], in_data89};
        src90 <= {src90[14:0], in_data90};
        src91 <= {src91[14:0], in_data91};
        src92 <= {src92[14:0], in_data92};
        src93 <= {src93[14:0], in_data93};
        src94 <= {src94[14:0], in_data94};
        src95 <= {src95[14:0], in_data95};
        src96 <= {src96[14:0], in_data96};
        src97 <= {src97[14:0], in_data97};
        src98 <= {src98[14:0], in_data98};
        src99 <= {src99[14:0], in_data99};
        src100 <= {src100[14:0], in_data100};
        src101 <= {src101[14:0], in_data101};
        src102 <= {src102[14:0], in_data102};
        src103 <= {src103[14:0], in_data103};
        src104 <= {src104[14:0], in_data104};
        src105 <= {src105[14:0], in_data105};
        src106 <= {src106[14:0], in_data106};
        src107 <= {src107[14:0], in_data107};
        src108 <= {src108[14:0], in_data108};
        src109 <= {src109[14:0], in_data109};
        src110 <= {src110[14:0], in_data110};
        src111 <= {src111[14:0], in_data111};
        src112 <= {src112[14:0], in_data112};
        src113 <= {src113[14:0], in_data113};
        src114 <= {src114[14:0], in_data114};
        src115 <= {src115[14:0], in_data115};
        src116 <= {src116[14:0], in_data116};
        src117 <= {src117[14:0], in_data117};
        src118 <= {src118[14:0], in_data118};
        src119 <= {src119[14:0], in_data119};
        src120 <= {src120[14:0], in_data120};
        src121 <= {src121[14:0], in_data121};
        src122 <= {src122[14:0], in_data122};
        src123 <= {src123[14:0], in_data123};
        src124 <= {src124[14:0], in_data124};
        src125 <= {src125[14:0], in_data125};
        src126 <= {src126[14:0], in_data126};
        src127 <= {src127[14:0], in_data127};
        src128 <= {src128[14:0], in_data128};
        src129 <= {src129[14:0], in_data129};
        src130 <= {src130[14:0], in_data130};
        src131 <= {src131[14:0], in_data131};
        src132 <= {src132[14:0], in_data132};
        src133 <= {src133[14:0], in_data133};
        src134 <= {src134[14:0], in_data134};
        src135 <= {src135[14:0], in_data135};
        src136 <= {src136[14:0], in_data136};
        src137 <= {src137[14:0], in_data137};
        src138 <= {src138[14:0], in_data138};
        src139 <= {src139[14:0], in_data139};
        src140 <= {src140[14:0], in_data140};
        src141 <= {src141[14:0], in_data141};
        src142 <= {src142[14:0], in_data142};
        src143 <= {src143[14:0], in_data143};
        src144 <= {src144[14:0], in_data144};
        src145 <= {src145[14:0], in_data145};
        src146 <= {src146[14:0], in_data146};
        src147 <= {src147[14:0], in_data147};
        src148 <= {src148[14:0], in_data148};
        src149 <= {src149[14:0], in_data149};
        src150 <= {src150[14:0], in_data150};
        src151 <= {src151[14:0], in_data151};
        src152 <= {src152[14:0], in_data152};
        src153 <= {src153[14:0], in_data153};
        src154 <= {src154[14:0], in_data154};
        src155 <= {src155[14:0], in_data155};
        src156 <= {src156[14:0], in_data156};
        src157 <= {src157[14:0], in_data157};
        src158 <= {src158[14:0], in_data158};
        src159 <= {src159[14:0], in_data159};
        src160 <= {src160[14:0], in_data160};
        src161 <= {src161[14:0], in_data161};
        src162 <= {src162[14:0], in_data162};
        src163 <= {src163[14:0], in_data163};
        src164 <= {src164[14:0], in_data164};
        src165 <= {src165[14:0], in_data165};
        src166 <= {src166[14:0], in_data166};
        src167 <= {src167[14:0], in_data167};
        src168 <= {src168[14:0], in_data168};
        src169 <= {src169[14:0], in_data169};
        src170 <= {src170[14:0], in_data170};
        src171 <= {src171[14:0], in_data171};
        src172 <= {src172[14:0], in_data172};
        src173 <= {src173[14:0], in_data173};
        src174 <= {src174[14:0], in_data174};
        src175 <= {src175[14:0], in_data175};
        src176 <= {src176[14:0], in_data176};
        src177 <= {src177[14:0], in_data177};
        src178 <= {src178[14:0], in_data178};
        src179 <= {src179[14:0], in_data179};
        src180 <= {src180[14:0], in_data180};
        src181 <= {src181[14:0], in_data181};
        src182 <= {src182[14:0], in_data182};
        src183 <= {src183[14:0], in_data183};
        src184 <= {src184[14:0], in_data184};
    end
endmodule

module compressor2_1_185_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    input [15:0]src64,
    input [15:0]src65,
    input [15:0]src66,
    input [15:0]src67,
    input [15:0]src68,
    input [15:0]src69,
    input [15:0]src70,
    input [15:0]src71,
    input [15:0]src72,
    input [15:0]src73,
    input [15:0]src74,
    input [15:0]src75,
    input [15:0]src76,
    input [15:0]src77,
    input [15:0]src78,
    input [15:0]src79,
    input [15:0]src80,
    input [15:0]src81,
    input [15:0]src82,
    input [15:0]src83,
    input [15:0]src84,
    input [15:0]src85,
    input [15:0]src86,
    input [15:0]src87,
    input [15:0]src88,
    input [15:0]src89,
    input [15:0]src90,
    input [15:0]src91,
    input [15:0]src92,
    input [15:0]src93,
    input [15:0]src94,
    input [15:0]src95,
    input [15:0]src96,
    input [15:0]src97,
    input [15:0]src98,
    input [15:0]src99,
    input [15:0]src100,
    input [15:0]src101,
    input [15:0]src102,
    input [15:0]src103,
    input [15:0]src104,
    input [15:0]src105,
    input [15:0]src106,
    input [15:0]src107,
    input [15:0]src108,
    input [15:0]src109,
    input [15:0]src110,
    input [15:0]src111,
    input [15:0]src112,
    input [15:0]src113,
    input [15:0]src114,
    input [15:0]src115,
    input [15:0]src116,
    input [15:0]src117,
    input [15:0]src118,
    input [15:0]src119,
    input [15:0]src120,
    input [15:0]src121,
    input [15:0]src122,
    input [15:0]src123,
    input [15:0]src124,
    input [15:0]src125,
    input [15:0]src126,
    input [15:0]src127,
    input [15:0]src128,
    input [15:0]src129,
    input [15:0]src130,
    input [15:0]src131,
    input [15:0]src132,
    input [15:0]src133,
    input [15:0]src134,
    input [15:0]src135,
    input [15:0]src136,
    input [15:0]src137,
    input [15:0]src138,
    input [15:0]src139,
    input [15:0]src140,
    input [15:0]src141,
    input [15:0]src142,
    input [15:0]src143,
    input [15:0]src144,
    input [15:0]src145,
    input [15:0]src146,
    input [15:0]src147,
    input [15:0]src148,
    input [15:0]src149,
    input [15:0]src150,
    input [15:0]src151,
    input [15:0]src152,
    input [15:0]src153,
    input [15:0]src154,
    input [15:0]src155,
    input [15:0]src156,
    input [15:0]src157,
    input [15:0]src158,
    input [15:0]src159,
    input [15:0]src160,
    input [15:0]src161,
    input [15:0]src162,
    input [15:0]src163,
    input [15:0]src164,
    input [15:0]src165,
    input [15:0]src166,
    input [15:0]src167,
    input [15:0]src168,
    input [15:0]src169,
    input [15:0]src170,
    input [15:0]src171,
    input [15:0]src172,
    input [15:0]src173,
    input [15:0]src174,
    input [15:0]src175,
    input [15:0]src176,
    input [15:0]src177,
    input [15:0]src178,
    input [15:0]src179,
    input [15:0]src180,
    input [15:0]src181,
    input [15:0]src182,
    input [15:0]src183,
    input [15:0]src184,
    output [23:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [0:0] comp_out22;
    wire [0:0] comp_out23;
    wire [24:0] out;
    compressor compressor_inst(
        .src0({src184[0], src183[0], src182[0], src181[0], src180[0], src179[0], src178[0], src177[0], src176[0], src175[0], src174[0], src173[0], src172[0], src171[0], src170[0], src169[0], src168[0], src167[0], src166[0], src165[0], src164[0], src163[0], src162[0], src161[0], src160[0], src159[0], src158[0], src157[0], src156[0], src155[0], src154[0], src153[0], src152[0], src151[0], src150[0], src149[0], src148[0], src147[0], src146[0], src145[0], src144[0], src143[0], src142[0], src141[0], src140[0], src139[0], src138[0], src137[0], src136[0], src135[0], src134[0], src133[0], src132[0], src131[0], src130[0], src129[0], src128[0], src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src184[1], src183[1], src182[1], src181[1], src180[1], src179[1], src178[1], src177[1], src176[1], src175[1], src174[1], src173[1], src172[1], src171[1], src170[1], src169[1], src168[1], src167[1], src166[1], src165[1], src164[1], src163[1], src162[1], src161[1], src160[1], src159[1], src158[1], src157[1], src156[1], src155[1], src154[1], src153[1], src152[1], src151[1], src150[1], src149[1], src148[1], src147[1], src146[1], src145[1], src144[1], src143[1], src142[1], src141[1], src140[1], src139[1], src138[1], src137[1], src136[1], src135[1], src134[1], src133[1], src132[1], src131[1], src130[1], src129[1], src128[1], src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src184[2], src183[2], src182[2], src181[2], src180[2], src179[2], src178[2], src177[2], src176[2], src175[2], src174[2], src173[2], src172[2], src171[2], src170[2], src169[2], src168[2], src167[2], src166[2], src165[2], src164[2], src163[2], src162[2], src161[2], src160[2], src159[2], src158[2], src157[2], src156[2], src155[2], src154[2], src153[2], src152[2], src151[2], src150[2], src149[2], src148[2], src147[2], src146[2], src145[2], src144[2], src143[2], src142[2], src141[2], src140[2], src139[2], src138[2], src137[2], src136[2], src135[2], src134[2], src133[2], src132[2], src131[2], src130[2], src129[2], src128[2], src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src184[3], src183[3], src182[3], src181[3], src180[3], src179[3], src178[3], src177[3], src176[3], src175[3], src174[3], src173[3], src172[3], src171[3], src170[3], src169[3], src168[3], src167[3], src166[3], src165[3], src164[3], src163[3], src162[3], src161[3], src160[3], src159[3], src158[3], src157[3], src156[3], src155[3], src154[3], src153[3], src152[3], src151[3], src150[3], src149[3], src148[3], src147[3], src146[3], src145[3], src144[3], src143[3], src142[3], src141[3], src140[3], src139[3], src138[3], src137[3], src136[3], src135[3], src134[3], src133[3], src132[3], src131[3], src130[3], src129[3], src128[3], src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src184[4], src183[4], src182[4], src181[4], src180[4], src179[4], src178[4], src177[4], src176[4], src175[4], src174[4], src173[4], src172[4], src171[4], src170[4], src169[4], src168[4], src167[4], src166[4], src165[4], src164[4], src163[4], src162[4], src161[4], src160[4], src159[4], src158[4], src157[4], src156[4], src155[4], src154[4], src153[4], src152[4], src151[4], src150[4], src149[4], src148[4], src147[4], src146[4], src145[4], src144[4], src143[4], src142[4], src141[4], src140[4], src139[4], src138[4], src137[4], src136[4], src135[4], src134[4], src133[4], src132[4], src131[4], src130[4], src129[4], src128[4], src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src184[5], src183[5], src182[5], src181[5], src180[5], src179[5], src178[5], src177[5], src176[5], src175[5], src174[5], src173[5], src172[5], src171[5], src170[5], src169[5], src168[5], src167[5], src166[5], src165[5], src164[5], src163[5], src162[5], src161[5], src160[5], src159[5], src158[5], src157[5], src156[5], src155[5], src154[5], src153[5], src152[5], src151[5], src150[5], src149[5], src148[5], src147[5], src146[5], src145[5], src144[5], src143[5], src142[5], src141[5], src140[5], src139[5], src138[5], src137[5], src136[5], src135[5], src134[5], src133[5], src132[5], src131[5], src130[5], src129[5], src128[5], src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src184[6], src183[6], src182[6], src181[6], src180[6], src179[6], src178[6], src177[6], src176[6], src175[6], src174[6], src173[6], src172[6], src171[6], src170[6], src169[6], src168[6], src167[6], src166[6], src165[6], src164[6], src163[6], src162[6], src161[6], src160[6], src159[6], src158[6], src157[6], src156[6], src155[6], src154[6], src153[6], src152[6], src151[6], src150[6], src149[6], src148[6], src147[6], src146[6], src145[6], src144[6], src143[6], src142[6], src141[6], src140[6], src139[6], src138[6], src137[6], src136[6], src135[6], src134[6], src133[6], src132[6], src131[6], src130[6], src129[6], src128[6], src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src184[7], src183[7], src182[7], src181[7], src180[7], src179[7], src178[7], src177[7], src176[7], src175[7], src174[7], src173[7], src172[7], src171[7], src170[7], src169[7], src168[7], src167[7], src166[7], src165[7], src164[7], src163[7], src162[7], src161[7], src160[7], src159[7], src158[7], src157[7], src156[7], src155[7], src154[7], src153[7], src152[7], src151[7], src150[7], src149[7], src148[7], src147[7], src146[7], src145[7], src144[7], src143[7], src142[7], src141[7], src140[7], src139[7], src138[7], src137[7], src136[7], src135[7], src134[7], src133[7], src132[7], src131[7], src130[7], src129[7], src128[7], src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src184[8], src183[8], src182[8], src181[8], src180[8], src179[8], src178[8], src177[8], src176[8], src175[8], src174[8], src173[8], src172[8], src171[8], src170[8], src169[8], src168[8], src167[8], src166[8], src165[8], src164[8], src163[8], src162[8], src161[8], src160[8], src159[8], src158[8], src157[8], src156[8], src155[8], src154[8], src153[8], src152[8], src151[8], src150[8], src149[8], src148[8], src147[8], src146[8], src145[8], src144[8], src143[8], src142[8], src141[8], src140[8], src139[8], src138[8], src137[8], src136[8], src135[8], src134[8], src133[8], src132[8], src131[8], src130[8], src129[8], src128[8], src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src184[9], src183[9], src182[9], src181[9], src180[9], src179[9], src178[9], src177[9], src176[9], src175[9], src174[9], src173[9], src172[9], src171[9], src170[9], src169[9], src168[9], src167[9], src166[9], src165[9], src164[9], src163[9], src162[9], src161[9], src160[9], src159[9], src158[9], src157[9], src156[9], src155[9], src154[9], src153[9], src152[9], src151[9], src150[9], src149[9], src148[9], src147[9], src146[9], src145[9], src144[9], src143[9], src142[9], src141[9], src140[9], src139[9], src138[9], src137[9], src136[9], src135[9], src134[9], src133[9], src132[9], src131[9], src130[9], src129[9], src128[9], src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src184[10], src183[10], src182[10], src181[10], src180[10], src179[10], src178[10], src177[10], src176[10], src175[10], src174[10], src173[10], src172[10], src171[10], src170[10], src169[10], src168[10], src167[10], src166[10], src165[10], src164[10], src163[10], src162[10], src161[10], src160[10], src159[10], src158[10], src157[10], src156[10], src155[10], src154[10], src153[10], src152[10], src151[10], src150[10], src149[10], src148[10], src147[10], src146[10], src145[10], src144[10], src143[10], src142[10], src141[10], src140[10], src139[10], src138[10], src137[10], src136[10], src135[10], src134[10], src133[10], src132[10], src131[10], src130[10], src129[10], src128[10], src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src184[11], src183[11], src182[11], src181[11], src180[11], src179[11], src178[11], src177[11], src176[11], src175[11], src174[11], src173[11], src172[11], src171[11], src170[11], src169[11], src168[11], src167[11], src166[11], src165[11], src164[11], src163[11], src162[11], src161[11], src160[11], src159[11], src158[11], src157[11], src156[11], src155[11], src154[11], src153[11], src152[11], src151[11], src150[11], src149[11], src148[11], src147[11], src146[11], src145[11], src144[11], src143[11], src142[11], src141[11], src140[11], src139[11], src138[11], src137[11], src136[11], src135[11], src134[11], src133[11], src132[11], src131[11], src130[11], src129[11], src128[11], src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src184[12], src183[12], src182[12], src181[12], src180[12], src179[12], src178[12], src177[12], src176[12], src175[12], src174[12], src173[12], src172[12], src171[12], src170[12], src169[12], src168[12], src167[12], src166[12], src165[12], src164[12], src163[12], src162[12], src161[12], src160[12], src159[12], src158[12], src157[12], src156[12], src155[12], src154[12], src153[12], src152[12], src151[12], src150[12], src149[12], src148[12], src147[12], src146[12], src145[12], src144[12], src143[12], src142[12], src141[12], src140[12], src139[12], src138[12], src137[12], src136[12], src135[12], src134[12], src133[12], src132[12], src131[12], src130[12], src129[12], src128[12], src127[12], src126[12], src125[12], src124[12], src123[12], src122[12], src121[12], src120[12], src119[12], src118[12], src117[12], src116[12], src115[12], src114[12], src113[12], src112[12], src111[12], src110[12], src109[12], src108[12], src107[12], src106[12], src105[12], src104[12], src103[12], src102[12], src101[12], src100[12], src99[12], src98[12], src97[12], src96[12], src95[12], src94[12], src93[12], src92[12], src91[12], src90[12], src89[12], src88[12], src87[12], src86[12], src85[12], src84[12], src83[12], src82[12], src81[12], src80[12], src79[12], src78[12], src77[12], src76[12], src75[12], src74[12], src73[12], src72[12], src71[12], src70[12], src69[12], src68[12], src67[12], src66[12], src65[12], src64[12], src63[12], src62[12], src61[12], src60[12], src59[12], src58[12], src57[12], src56[12], src55[12], src54[12], src53[12], src52[12], src51[12], src50[12], src49[12], src48[12], src47[12], src46[12], src45[12], src44[12], src43[12], src42[12], src41[12], src40[12], src39[12], src38[12], src37[12], src36[12], src35[12], src34[12], src33[12], src32[12], src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src184[13], src183[13], src182[13], src181[13], src180[13], src179[13], src178[13], src177[13], src176[13], src175[13], src174[13], src173[13], src172[13], src171[13], src170[13], src169[13], src168[13], src167[13], src166[13], src165[13], src164[13], src163[13], src162[13], src161[13], src160[13], src159[13], src158[13], src157[13], src156[13], src155[13], src154[13], src153[13], src152[13], src151[13], src150[13], src149[13], src148[13], src147[13], src146[13], src145[13], src144[13], src143[13], src142[13], src141[13], src140[13], src139[13], src138[13], src137[13], src136[13], src135[13], src134[13], src133[13], src132[13], src131[13], src130[13], src129[13], src128[13], src127[13], src126[13], src125[13], src124[13], src123[13], src122[13], src121[13], src120[13], src119[13], src118[13], src117[13], src116[13], src115[13], src114[13], src113[13], src112[13], src111[13], src110[13], src109[13], src108[13], src107[13], src106[13], src105[13], src104[13], src103[13], src102[13], src101[13], src100[13], src99[13], src98[13], src97[13], src96[13], src95[13], src94[13], src93[13], src92[13], src91[13], src90[13], src89[13], src88[13], src87[13], src86[13], src85[13], src84[13], src83[13], src82[13], src81[13], src80[13], src79[13], src78[13], src77[13], src76[13], src75[13], src74[13], src73[13], src72[13], src71[13], src70[13], src69[13], src68[13], src67[13], src66[13], src65[13], src64[13], src63[13], src62[13], src61[13], src60[13], src59[13], src58[13], src57[13], src56[13], src55[13], src54[13], src53[13], src52[13], src51[13], src50[13], src49[13], src48[13], src47[13], src46[13], src45[13], src44[13], src43[13], src42[13], src41[13], src40[13], src39[13], src38[13], src37[13], src36[13], src35[13], src34[13], src33[13], src32[13], src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src184[14], src183[14], src182[14], src181[14], src180[14], src179[14], src178[14], src177[14], src176[14], src175[14], src174[14], src173[14], src172[14], src171[14], src170[14], src169[14], src168[14], src167[14], src166[14], src165[14], src164[14], src163[14], src162[14], src161[14], src160[14], src159[14], src158[14], src157[14], src156[14], src155[14], src154[14], src153[14], src152[14], src151[14], src150[14], src149[14], src148[14], src147[14], src146[14], src145[14], src144[14], src143[14], src142[14], src141[14], src140[14], src139[14], src138[14], src137[14], src136[14], src135[14], src134[14], src133[14], src132[14], src131[14], src130[14], src129[14], src128[14], src127[14], src126[14], src125[14], src124[14], src123[14], src122[14], src121[14], src120[14], src119[14], src118[14], src117[14], src116[14], src115[14], src114[14], src113[14], src112[14], src111[14], src110[14], src109[14], src108[14], src107[14], src106[14], src105[14], src104[14], src103[14], src102[14], src101[14], src100[14], src99[14], src98[14], src97[14], src96[14], src95[14], src94[14], src93[14], src92[14], src91[14], src90[14], src89[14], src88[14], src87[14], src86[14], src85[14], src84[14], src83[14], src82[14], src81[14], src80[14], src79[14], src78[14], src77[14], src76[14], src75[14], src74[14], src73[14], src72[14], src71[14], src70[14], src69[14], src68[14], src67[14], src66[14], src65[14], src64[14], src63[14], src62[14], src61[14], src60[14], src59[14], src58[14], src57[14], src56[14], src55[14], src54[14], src53[14], src52[14], src51[14], src50[14], src49[14], src48[14], src47[14], src46[14], src45[14], src44[14], src43[14], src42[14], src41[14], src40[14], src39[14], src38[14], src37[14], src36[14], src35[14], src34[14], src33[14], src32[14], src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src184[15], src183[15], src182[15], src181[15], src180[15], src179[15], src178[15], src177[15], src176[15], src175[15], src174[15], src173[15], src172[15], src171[15], src170[15], src169[15], src168[15], src167[15], src166[15], src165[15], src164[15], src163[15], src162[15], src161[15], src160[15], src159[15], src158[15], src157[15], src156[15], src155[15], src154[15], src153[15], src152[15], src151[15], src150[15], src149[15], src148[15], src147[15], src146[15], src145[15], src144[15], src143[15], src142[15], src141[15], src140[15], src139[15], src138[15], src137[15], src136[15], src135[15], src134[15], src133[15], src132[15], src131[15], src130[15], src129[15], src128[15], src127[15], src126[15], src125[15], src124[15], src123[15], src122[15], src121[15], src120[15], src119[15], src118[15], src117[15], src116[15], src115[15], src114[15], src113[15], src112[15], src111[15], src110[15], src109[15], src108[15], src107[15], src106[15], src105[15], src104[15], src103[15], src102[15], src101[15], src100[15], src99[15], src98[15], src97[15], src96[15], src95[15], src94[15], src93[15], src92[15], src91[15], src90[15], src89[15], src88[15], src87[15], src86[15], src85[15], src84[15], src83[15], src82[15], src81[15], src80[15], src79[15], src78[15], src77[15], src76[15], src75[15], src74[15], src73[15], src72[15], src71[15], src70[15], src69[15], src68[15], src67[15], src66[15], src65[15], src64[15], src63[15], src62[15], src61[15], src60[15], src59[15], src58[15], src57[15], src56[15], src55[15], src54[15], src53[15], src52[15], src51[15], src50[15], src49[15], src48[15], src47[15], src46[15], src45[15], src44[15], src43[15], src42[15], src41[15], src40[15], src39[15], src38[15], src37[15], src36[15], src35[15], src34[15], src33[15], src32[15], src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23)
    );
    rowadder2_1_24 rowadder2_1inst(
        .src0({comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[23:0];
endmodule
module compressor (
      input wire [184:0] src0,
      input wire [184:0] src1,
      input wire [184:0] src2,
      input wire [184:0] src3,
      input wire [184:0] src4,
      input wire [184:0] src5,
      input wire [184:0] src6,
      input wire [184:0] src7,
      input wire [184:0] src8,
      input wire [184:0] src9,
      input wire [184:0] src10,
      input wire [184:0] src11,
      input wire [184:0] src12,
      input wire [184:0] src13,
      input wire [184:0] src14,
      input wire [184:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [0:0] dst22,
      output wire [0:0] dst23);

   wire [184:0] stage0_0;
   wire [184:0] stage0_1;
   wire [184:0] stage0_2;
   wire [184:0] stage0_3;
   wire [184:0] stage0_4;
   wire [184:0] stage0_5;
   wire [184:0] stage0_6;
   wire [184:0] stage0_7;
   wire [184:0] stage0_8;
   wire [184:0] stage0_9;
   wire [184:0] stage0_10;
   wire [184:0] stage0_11;
   wire [184:0] stage0_12;
   wire [184:0] stage0_13;
   wire [184:0] stage0_14;
   wire [184:0] stage0_15;
   wire [48:0] stage1_0;
   wire [55:0] stage1_1;
   wire [66:0] stage1_2;
   wire [81:0] stage1_3;
   wire [84:0] stage1_4;
   wire [129:0] stage1_5;
   wire [63:0] stage1_6;
   wire [89:0] stage1_7;
   wire [80:0] stage1_8;
   wire [83:0] stage1_9;
   wire [93:0] stage1_10;
   wire [58:0] stage1_11;
   wire [104:0] stage1_12;
   wire [85:0] stage1_13;
   wire [68:0] stage1_14;
   wire [81:0] stage1_15;
   wire [52:0] stage1_16;
   wire [26:0] stage1_17;
   wire [12:0] stage2_0;
   wire [19:0] stage2_1;
   wire [24:0] stage2_2;
   wire [30:0] stage2_3;
   wire [37:0] stage2_4;
   wire [33:0] stage2_5;
   wire [37:0] stage2_6;
   wire [39:0] stage2_7;
   wire [45:0] stage2_8;
   wire [31:0] stage2_9;
   wire [39:0] stage2_10;
   wire [32:0] stage2_11;
   wire [51:0] stage2_12;
   wire [39:0] stage2_13;
   wire [36:0] stage2_14;
   wire [27:0] stage2_15;
   wire [27:0] stage2_16;
   wire [24:0] stage2_17;
   wire [11:0] stage2_18;
   wire [3:0] stage2_19;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [11:0] stage3_4;
   wire [14:0] stage3_5;
   wire [15:0] stage3_6;
   wire [21:0] stage3_7;
   wire [18:0] stage3_8;
   wire [14:0] stage3_9;
   wire [20:0] stage3_10;
   wire [16:0] stage3_11;
   wire [21:0] stage3_12;
   wire [18:0] stage3_13;
   wire [15:0] stage3_14;
   wire [13:0] stage3_15;
   wire [14:0] stage3_16;
   wire [21:0] stage3_17;
   wire [5:0] stage3_18;
   wire [7:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage4_0;
   wire [5:0] stage4_1;
   wire [3:0] stage4_2;
   wire [7:0] stage4_3;
   wire [3:0] stage4_4;
   wire [5:0] stage4_5;
   wire [5:0] stage4_6;
   wire [10:0] stage4_7;
   wire [6:0] stage4_8;
   wire [7:0] stage4_9;
   wire [7:0] stage4_10;
   wire [13:0] stage4_11;
   wire [7:0] stage4_12;
   wire [7:0] stage4_13;
   wire [7:0] stage4_14;
   wire [6:0] stage4_15;
   wire [5:0] stage4_16;
   wire [8:0] stage4_17;
   wire [8:0] stage4_18;
   wire [4:0] stage4_19;
   wire [3:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [3:0] stage5_4;
   wire [7:0] stage5_5;
   wire [1:0] stage5_6;
   wire [4:0] stage5_7;
   wire [2:0] stage5_8;
   wire [3:0] stage5_9;
   wire [3:0] stage5_10;
   wire [3:0] stage5_11;
   wire [3:0] stage5_12;
   wire [5:0] stage5_13;
   wire [4:0] stage5_14;
   wire [2:0] stage5_15;
   wire [1:0] stage5_16;
   wire [3:0] stage5_17;
   wire [3:0] stage5_18;
   wire [2:0] stage5_19;
   wire [2:0] stage5_20;
   wire [2:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [0:0] stage6_22;
   wire [0:0] stage6_23;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc2135_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[12]},
      {stage0_3[24], stage0_3[25]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc615_5 gpc25 (
      {stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[39]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc615_5 gpc26 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_1[40]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc615_5 gpc27 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[41]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc615_5 gpc28 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[42]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc615_5 gpc29 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_1[43]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc615_5 gpc30 (
      {stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166]},
      {stage0_1[44]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[0],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[1],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[2],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[3],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[4],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[5],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[6],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[7],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[8],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[9],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[10],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[11],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[12],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[13],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[14],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[15],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[16],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[17],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[18],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[19],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[20],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157]},
      {stage1_5[21],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163]},
      {stage1_5[22],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[23],stage1_4[54],stage1_3[54],stage1_2[54]}
   );
   gpc606_5 gpc55 (
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[24],stage1_4[55],stage1_3[55],stage1_2[55]}
   );
   gpc606_5 gpc56 (
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[25],stage1_4[56],stage1_3[56],stage1_2[56]}
   );
   gpc606_5 gpc57 (
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[26],stage1_4[57],stage1_3[57],stage1_2[57]}
   );
   gpc606_5 gpc58 (
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[27],stage1_4[58],stage1_3[58],stage1_2[58]}
   );
   gpc606_5 gpc59 (
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[28],stage1_4[59],stage1_3[59],stage1_2[59]}
   );
   gpc606_5 gpc60 (
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[29],stage1_4[60],stage1_3[60],stage1_2[60]}
   );
   gpc615_5 gpc61 (
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage0_3[164]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[30],stage1_4[61],stage1_3[61],stage1_2[61]}
   );
   gpc615_5 gpc62 (
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172]},
      {stage0_3[165]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[31],stage1_4[62],stage1_3[62],stage1_2[62]}
   );
   gpc615_5 gpc63 (
      {stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177]},
      {stage0_3[166]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[32],stage1_4[63],stage1_3[63],stage1_2[63]}
   );
   gpc615_5 gpc64 (
      {stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage0_3[167]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[33],stage1_4[64],stage1_3[64],stage1_2[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[11],stage1_5[34],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[12],stage1_5[35],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[13],stage1_5[36],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[14],stage1_5[37],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[15],stage1_5[38],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[16],stage1_5[39],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[17],stage1_5[40],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[18],stage1_5[41],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[19],stage1_5[42],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[20],stage1_5[43],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[21],stage1_5[44],stage1_4[75]}
   );
   gpc606_5 gpc76 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[22],stage1_5[45],stage1_4[76]}
   );
   gpc606_5 gpc77 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[23],stage1_5[46],stage1_4[77]}
   );
   gpc606_5 gpc78 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[24],stage1_5[47],stage1_4[78]}
   );
   gpc606_5 gpc79 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[25],stage1_5[48],stage1_4[79]}
   );
   gpc606_5 gpc80 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[26],stage1_5[49],stage1_4[80]}
   );
   gpc606_5 gpc81 (
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[27],stage1_5[50],stage1_4[81]}
   );
   gpc606_5 gpc82 (
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[28],stage1_5[51],stage1_4[82]}
   );
   gpc606_5 gpc83 (
      {stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[29],stage1_5[52],stage1_4[83]}
   );
   gpc615_5 gpc84 (
      {stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_5[0]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[30],stage1_5[53],stage1_4[84]}
   );
   gpc606_5 gpc85 (
      {stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[20],stage1_7[20],stage1_6[31],stage1_5[54]}
   );
   gpc606_5 gpc86 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[21],stage1_7[21],stage1_6[32],stage1_5[55]}
   );
   gpc606_5 gpc87 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[22],stage1_7[22],stage1_6[33],stage1_5[56]}
   );
   gpc606_5 gpc88 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[23],stage1_7[23],stage1_6[34],stage1_5[57]}
   );
   gpc606_5 gpc89 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[24],stage1_7[24],stage1_6[35],stage1_5[58]}
   );
   gpc606_5 gpc90 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[25],stage1_7[25],stage1_6[36],stage1_5[59]}
   );
   gpc606_5 gpc91 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[26],stage1_7[26],stage1_6[37],stage1_5[60]}
   );
   gpc606_5 gpc92 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[27],stage1_7[27],stage1_6[38],stage1_5[61]}
   );
   gpc606_5 gpc93 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[28],stage1_7[28],stage1_6[39],stage1_5[62]}
   );
   gpc606_5 gpc94 (
      {stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[29],stage1_7[29],stage1_6[40],stage1_5[63]}
   );
   gpc606_5 gpc95 (
      {stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[30],stage1_7[30],stage1_6[41],stage1_5[64]}
   );
   gpc606_5 gpc96 (
      {stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[31],stage1_7[31],stage1_6[42],stage1_5[65]}
   );
   gpc606_5 gpc97 (
      {stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[32],stage1_7[32],stage1_6[43],stage1_5[66]}
   );
   gpc606_5 gpc98 (
      {stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[33],stage1_7[33],stage1_6[44],stage1_5[67]}
   );
   gpc606_5 gpc99 (
      {stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[34],stage1_7[34],stage1_6[45],stage1_5[68]}
   );
   gpc606_5 gpc100 (
      {stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[35],stage1_7[35],stage1_6[46],stage1_5[69]}
   );
   gpc615_5 gpc101 (
      {stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_6[120]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[36],stage1_7[36],stage1_6[47],stage1_5[70]}
   );
   gpc615_5 gpc102 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106]},
      {stage0_6[121]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[37],stage1_7[37],stage1_6[48],stage1_5[71]}
   );
   gpc615_5 gpc103 (
      {stage0_5[107], stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111]},
      {stage0_6[122]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[38],stage1_7[38],stage1_6[49],stage1_5[72]}
   );
   gpc615_5 gpc104 (
      {stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116]},
      {stage0_6[123]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[39],stage1_7[39],stage1_6[50],stage1_5[73]}
   );
   gpc615_5 gpc105 (
      {stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121]},
      {stage0_6[124]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[40],stage1_7[40],stage1_6[51],stage1_5[74]}
   );
   gpc615_5 gpc106 (
      {stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126]},
      {stage0_6[125]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[41],stage1_7[41],stage1_6[52],stage1_5[75]}
   );
   gpc615_5 gpc107 (
      {stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_6[126]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[42],stage1_7[42],stage1_6[53],stage1_5[76]}
   );
   gpc606_5 gpc108 (
      {stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[23],stage1_8[43],stage1_7[43],stage1_6[54]}
   );
   gpc606_5 gpc109 (
      {stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[24],stage1_8[44],stage1_7[44],stage1_6[55]}
   );
   gpc606_5 gpc110 (
      {stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143], stage0_6[144]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[25],stage1_8[45],stage1_7[45],stage1_6[56]}
   );
   gpc606_5 gpc111 (
      {stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149], stage0_6[150]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[26],stage1_8[46],stage1_7[46],stage1_6[57]}
   );
   gpc606_5 gpc112 (
      {stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155], stage0_6[156]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[27],stage1_8[47],stage1_7[47],stage1_6[58]}
   );
   gpc606_5 gpc113 (
      {stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161], stage0_6[162]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[28],stage1_8[48],stage1_7[48],stage1_6[59]}
   );
   gpc606_5 gpc114 (
      {stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167], stage0_6[168]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[29],stage1_8[49],stage1_7[49],stage1_6[60]}
   );
   gpc606_5 gpc115 (
      {stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173], stage0_6[174]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[30],stage1_8[50],stage1_7[50],stage1_6[61]}
   );
   gpc615_5 gpc116 (
      {stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage0_7[138]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[31],stage1_8[51],stage1_7[51],stage1_6[62]}
   );
   gpc615_5 gpc117 (
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184]},
      {stage0_7[139]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[32],stage1_8[52],stage1_7[52],stage1_6[63]}
   );
   gpc615_5 gpc118 (
      {stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143], stage0_7[144]},
      {stage0_8[60]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[10],stage1_9[33],stage1_8[53],stage1_7[53]}
   );
   gpc615_5 gpc119 (
      {stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage0_8[61]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[11],stage1_9[34],stage1_8[54],stage1_7[54]}
   );
   gpc606_5 gpc120 (
      {stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[12],stage1_9[35],stage1_8[55]}
   );
   gpc615_5 gpc121 (
      {stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_9[12]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[13],stage1_9[36],stage1_8[56]}
   );
   gpc615_5 gpc122 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_9[13]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[14],stage1_9[37],stage1_8[57]}
   );
   gpc615_5 gpc123 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82]},
      {stage0_9[14]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[15],stage1_9[38],stage1_8[58]}
   );
   gpc615_5 gpc124 (
      {stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_9[15]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[16],stage1_9[39],stage1_8[59]}
   );
   gpc615_5 gpc125 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92]},
      {stage0_9[16]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[17],stage1_9[40],stage1_8[60]}
   );
   gpc615_5 gpc126 (
      {stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_9[17]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[18],stage1_9[41],stage1_8[61]}
   );
   gpc615_5 gpc127 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_9[18]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[19],stage1_9[42],stage1_8[62]}
   );
   gpc615_5 gpc128 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_9[19]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[20],stage1_9[43],stage1_8[63]}
   );
   gpc615_5 gpc129 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_9[20]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[21],stage1_9[44],stage1_8[64]}
   );
   gpc615_5 gpc130 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_9[21]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[22],stage1_9[45],stage1_8[65]}
   );
   gpc615_5 gpc131 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[22]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[23],stage1_9[46],stage1_8[66]}
   );
   gpc615_5 gpc132 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[23]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[24],stage1_9[47],stage1_8[67]}
   );
   gpc615_5 gpc133 (
      {stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_9[24]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[25],stage1_9[48],stage1_8[68]}
   );
   gpc615_5 gpc134 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_9[25]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[26],stage1_9[49],stage1_8[69]}
   );
   gpc615_5 gpc135 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142]},
      {stage0_9[26]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[17],stage1_10[27],stage1_9[50],stage1_8[70]}
   );
   gpc615_5 gpc136 (
      {stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147]},
      {stage0_9[27]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[18],stage1_10[28],stage1_9[51],stage1_8[71]}
   );
   gpc615_5 gpc137 (
      {stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152]},
      {stage0_9[28]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[19],stage1_10[29],stage1_9[52],stage1_8[72]}
   );
   gpc615_5 gpc138 (
      {stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_9[29]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[20],stage1_10[30],stage1_9[53],stage1_8[73]}
   );
   gpc615_5 gpc139 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_9[30]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[21],stage1_10[31],stage1_9[54],stage1_8[74]}
   );
   gpc615_5 gpc140 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_9[31]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[22],stage1_10[32],stage1_9[55],stage1_8[75]}
   );
   gpc615_5 gpc141 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172]},
      {stage0_9[32]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[23],stage1_10[33],stage1_9[56],stage1_8[76]}
   );
   gpc615_5 gpc142 (
      {stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_9[33]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[24],stage1_10[34],stage1_9[57],stage1_8[77]}
   );
   gpc615_5 gpc143 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_9[34]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[25],stage1_10[35],stage1_9[58],stage1_8[78]}
   );
   gpc606_5 gpc144 (
      {stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[24],stage1_11[26],stage1_10[36],stage1_9[59]}
   );
   gpc606_5 gpc145 (
      {stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[25],stage1_11[27],stage1_10[37],stage1_9[60]}
   );
   gpc606_5 gpc146 (
      {stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[26],stage1_11[28],stage1_10[38],stage1_9[61]}
   );
   gpc606_5 gpc147 (
      {stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[27],stage1_11[29],stage1_10[39],stage1_9[62]}
   );
   gpc606_5 gpc148 (
      {stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[28],stage1_11[30],stage1_10[40],stage1_9[63]}
   );
   gpc606_5 gpc149 (
      {stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[29],stage1_11[31],stage1_10[41],stage1_9[64]}
   );
   gpc606_5 gpc150 (
      {stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[30],stage1_11[32],stage1_10[42],stage1_9[65]}
   );
   gpc606_5 gpc151 (
      {stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[31],stage1_11[33],stage1_10[43],stage1_9[66]}
   );
   gpc606_5 gpc152 (
      {stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[32],stage1_11[34],stage1_10[44],stage1_9[67]}
   );
   gpc606_5 gpc153 (
      {stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[33],stage1_11[35],stage1_10[45],stage1_9[68]}
   );
   gpc606_5 gpc154 (
      {stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[34],stage1_11[36],stage1_10[46],stage1_9[69]}
   );
   gpc606_5 gpc155 (
      {stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[35],stage1_11[37],stage1_10[47],stage1_9[70]}
   );
   gpc606_5 gpc156 (
      {stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[36],stage1_11[38],stage1_10[48],stage1_9[71]}
   );
   gpc606_5 gpc157 (
      {stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[37],stage1_11[39],stage1_10[49],stage1_9[72]}
   );
   gpc606_5 gpc158 (
      {stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[38],stage1_11[40],stage1_10[50],stage1_9[73]}
   );
   gpc606_5 gpc159 (
      {stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[39],stage1_11[41],stage1_10[51],stage1_9[74]}
   );
   gpc606_5 gpc160 (
      {stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[40],stage1_11[42],stage1_10[52],stage1_9[75]}
   );
   gpc606_5 gpc161 (
      {stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[41],stage1_11[43],stage1_10[53],stage1_9[76]}
   );
   gpc606_5 gpc162 (
      {stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[42],stage1_11[44],stage1_10[54],stage1_9[77]}
   );
   gpc606_5 gpc163 (
      {stage0_9[149], stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[43],stage1_11[45],stage1_10[55],stage1_9[78]}
   );
   gpc606_5 gpc164 (
      {stage0_9[155], stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[44],stage1_11[46],stage1_10[56],stage1_9[79]}
   );
   gpc606_5 gpc165 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[45],stage1_11[47],stage1_10[57],stage1_9[80]}
   );
   gpc606_5 gpc166 (
      {stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[46],stage1_11[48],stage1_10[58],stage1_9[81]}
   );
   gpc606_5 gpc167 (
      {stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[47],stage1_11[49],stage1_10[59],stage1_9[82]}
   );
   gpc606_5 gpc168 (
      {stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[48],stage1_11[50],stage1_10[60],stage1_9[83]}
   );
   gpc615_5 gpc169 (
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148]},
      {stage0_11[150]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[25],stage1_12[49],stage1_11[51],stage1_10[61]}
   );
   gpc615_5 gpc170 (
      {stage0_10[149], stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153]},
      {stage0_11[151]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[26],stage1_12[50],stage1_11[52],stage1_10[62]}
   );
   gpc606_5 gpc171 (
      {stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[27],stage1_12[51],stage1_11[53]}
   );
   gpc606_5 gpc172 (
      {stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[28],stage1_12[52],stage1_11[54]}
   );
   gpc606_5 gpc173 (
      {stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[4],stage1_13[29],stage1_12[53],stage1_11[55]}
   );
   gpc615_5 gpc174 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[12]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[5],stage1_13[30],stage1_12[54],stage1_11[56]}
   );
   gpc615_5 gpc175 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[13]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[6],stage1_13[31],stage1_12[55],stage1_11[57]}
   );
   gpc615_5 gpc176 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[14]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[7],stage1_13[32],stage1_12[56],stage1_11[58]}
   );
   gpc606_5 gpc177 (
      {stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[6],stage1_14[8],stage1_13[33],stage1_12[57]}
   );
   gpc606_5 gpc178 (
      {stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[7],stage1_14[9],stage1_13[34],stage1_12[58]}
   );
   gpc606_5 gpc179 (
      {stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[8],stage1_14[10],stage1_13[35],stage1_12[59]}
   );
   gpc606_5 gpc180 (
      {stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[9],stage1_14[11],stage1_13[36],stage1_12[60]}
   );
   gpc606_5 gpc181 (
      {stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[10],stage1_14[12],stage1_13[37],stage1_12[61]}
   );
   gpc606_5 gpc182 (
      {stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[11],stage1_14[13],stage1_13[38],stage1_12[62]}
   );
   gpc606_5 gpc183 (
      {stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[12],stage1_14[14],stage1_13[39],stage1_12[63]}
   );
   gpc606_5 gpc184 (
      {stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[13],stage1_14[15],stage1_13[40],stage1_12[64]}
   );
   gpc606_5 gpc185 (
      {stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67], stage0_12[68]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[14],stage1_14[16],stage1_13[41],stage1_12[65]}
   );
   gpc606_5 gpc186 (
      {stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73], stage0_12[74]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[15],stage1_14[17],stage1_13[42],stage1_12[66]}
   );
   gpc606_5 gpc187 (
      {stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79], stage0_12[80]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[16],stage1_14[18],stage1_13[43],stage1_12[67]}
   );
   gpc606_5 gpc188 (
      {stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85], stage0_12[86]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[17],stage1_14[19],stage1_13[44],stage1_12[68]}
   );
   gpc606_5 gpc189 (
      {stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91], stage0_12[92]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[18],stage1_14[20],stage1_13[45],stage1_12[69]}
   );
   gpc606_5 gpc190 (
      {stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[19],stage1_14[21],stage1_13[46],stage1_12[70]}
   );
   gpc606_5 gpc191 (
      {stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[20],stage1_14[22],stage1_13[47],stage1_12[71]}
   );
   gpc606_5 gpc192 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[21],stage1_14[23],stage1_13[48],stage1_12[72]}
   );
   gpc606_5 gpc193 (
      {stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[22],stage1_14[24],stage1_13[49],stage1_12[73]}
   );
   gpc606_5 gpc194 (
      {stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[23],stage1_14[25],stage1_13[50],stage1_12[74]}
   );
   gpc615_5 gpc195 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_13[36]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[24],stage1_14[26],stage1_13[51],stage1_12[75]}
   );
   gpc615_5 gpc196 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132]},
      {stage0_13[37]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[25],stage1_14[27],stage1_13[52],stage1_12[76]}
   );
   gpc615_5 gpc197 (
      {stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_13[38]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[26],stage1_14[28],stage1_13[53],stage1_12[77]}
   );
   gpc615_5 gpc198 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142]},
      {stage0_13[39]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[27],stage1_14[29],stage1_13[54],stage1_12[78]}
   );
   gpc615_5 gpc199 (
      {stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_13[40]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[28],stage1_14[30],stage1_13[55],stage1_12[79]}
   );
   gpc615_5 gpc200 (
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152]},
      {stage0_13[41]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[29],stage1_14[31],stage1_13[56],stage1_12[80]}
   );
   gpc615_5 gpc201 (
      {stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157]},
      {stage0_13[42]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[30],stage1_14[32],stage1_13[57],stage1_12[81]}
   );
   gpc615_5 gpc202 (
      {stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161], stage0_12[162]},
      {stage0_13[43]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[31],stage1_14[33],stage1_13[58],stage1_12[82]}
   );
   gpc606_5 gpc203 (
      {stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[26],stage1_15[32],stage1_14[34],stage1_13[59]}
   );
   gpc606_5 gpc204 (
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[27],stage1_15[33],stage1_14[35],stage1_13[60]}
   );
   gpc606_5 gpc205 (
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[28],stage1_15[34],stage1_14[36],stage1_13[61]}
   );
   gpc606_5 gpc206 (
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[29],stage1_15[35],stage1_14[37],stage1_13[62]}
   );
   gpc606_5 gpc207 (
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[30],stage1_15[36],stage1_14[38],stage1_13[63]}
   );
   gpc606_5 gpc208 (
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[31],stage1_15[37],stage1_14[39],stage1_13[64]}
   );
   gpc615_5 gpc209 (
      {stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83], stage0_13[84]},
      {stage0_14[156]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[32],stage1_15[38],stage1_14[40],stage1_13[65]}
   );
   gpc615_5 gpc210 (
      {stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_14[157]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[33],stage1_15[39],stage1_14[41],stage1_13[66]}
   );
   gpc615_5 gpc211 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94]},
      {stage0_14[158]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[34],stage1_15[40],stage1_14[42],stage1_13[67]}
   );
   gpc615_5 gpc212 (
      {stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_14[159]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[35],stage1_15[41],stage1_14[43],stage1_13[68]}
   );
   gpc615_5 gpc213 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104]},
      {stage0_14[160]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[36],stage1_15[42],stage1_14[44],stage1_13[69]}
   );
   gpc615_5 gpc214 (
      {stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109]},
      {stage0_14[161]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[37],stage1_15[43],stage1_14[45],stage1_13[70]}
   );
   gpc615_5 gpc215 (
      {stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114]},
      {stage0_14[162]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[38],stage1_15[44],stage1_14[46],stage1_13[71]}
   );
   gpc615_5 gpc216 (
      {stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_14[163]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[39],stage1_15[45],stage1_14[47],stage1_13[72]}
   );
   gpc615_5 gpc217 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124]},
      {stage0_14[164]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[40],stage1_15[46],stage1_14[48],stage1_13[73]}
   );
   gpc615_5 gpc218 (
      {stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_14[165]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[41],stage1_15[47],stage1_14[49],stage1_13[74]}
   );
   gpc615_5 gpc219 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134]},
      {stage0_14[166]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[42],stage1_15[48],stage1_14[50],stage1_13[75]}
   );
   gpc615_5 gpc220 (
      {stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139]},
      {stage0_14[167]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[43],stage1_15[49],stage1_14[51],stage1_13[76]}
   );
   gpc615_5 gpc221 (
      {stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144]},
      {stage0_14[168]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[44],stage1_15[50],stage1_14[52],stage1_13[77]}
   );
   gpc615_5 gpc222 (
      {stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_14[169]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[45],stage1_15[51],stage1_14[53],stage1_13[78]}
   );
   gpc615_5 gpc223 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154]},
      {stage0_14[170]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[46],stage1_15[52],stage1_14[54],stage1_13[79]}
   );
   gpc615_5 gpc224 (
      {stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_14[171]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[47],stage1_15[53],stage1_14[55],stage1_13[80]}
   );
   gpc615_5 gpc225 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_14[172]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[48],stage1_15[54],stage1_14[56],stage1_13[81]}
   );
   gpc615_5 gpc226 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169]},
      {stage0_14[173]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[49],stage1_15[55],stage1_14[57],stage1_13[82]}
   );
   gpc615_5 gpc227 (
      {stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174]},
      {stage0_14[174]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[50],stage1_15[56],stage1_14[58],stage1_13[83]}
   );
   gpc615_5 gpc228 (
      {stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_14[175]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[51],stage1_15[57],stage1_14[59],stage1_13[84]}
   );
   gpc615_5 gpc229 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184]},
      {stage0_14[176]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[52],stage1_15[58],stage1_14[60],stage1_13[85]}
   );
   gpc1_1 gpc230 (
      {stage0_0[167]},
      {stage1_0[31]}
   );
   gpc1_1 gpc231 (
      {stage0_0[168]},
      {stage1_0[32]}
   );
   gpc1_1 gpc232 (
      {stage0_0[169]},
      {stage1_0[33]}
   );
   gpc1_1 gpc233 (
      {stage0_0[170]},
      {stage1_0[34]}
   );
   gpc1_1 gpc234 (
      {stage0_0[171]},
      {stage1_0[35]}
   );
   gpc1_1 gpc235 (
      {stage0_0[172]},
      {stage1_0[36]}
   );
   gpc1_1 gpc236 (
      {stage0_0[173]},
      {stage1_0[37]}
   );
   gpc1_1 gpc237 (
      {stage0_0[174]},
      {stage1_0[38]}
   );
   gpc1_1 gpc238 (
      {stage0_0[175]},
      {stage1_0[39]}
   );
   gpc1_1 gpc239 (
      {stage0_0[176]},
      {stage1_0[40]}
   );
   gpc1_1 gpc240 (
      {stage0_0[177]},
      {stage1_0[41]}
   );
   gpc1_1 gpc241 (
      {stage0_0[178]},
      {stage1_0[42]}
   );
   gpc1_1 gpc242 (
      {stage0_0[179]},
      {stage1_0[43]}
   );
   gpc1_1 gpc243 (
      {stage0_0[180]},
      {stage1_0[44]}
   );
   gpc1_1 gpc244 (
      {stage0_0[181]},
      {stage1_0[45]}
   );
   gpc1_1 gpc245 (
      {stage0_0[182]},
      {stage1_0[46]}
   );
   gpc1_1 gpc246 (
      {stage0_0[183]},
      {stage1_0[47]}
   );
   gpc1_1 gpc247 (
      {stage0_0[184]},
      {stage1_0[48]}
   );
   gpc1_1 gpc248 (
      {stage0_1[183]},
      {stage1_1[54]}
   );
   gpc1_1 gpc249 (
      {stage0_1[184]},
      {stage1_1[55]}
   );
   gpc1_1 gpc250 (
      {stage0_2[183]},
      {stage1_2[65]}
   );
   gpc1_1 gpc251 (
      {stage0_2[184]},
      {stage1_2[66]}
   );
   gpc1_1 gpc252 (
      {stage0_3[168]},
      {stage1_3[65]}
   );
   gpc1_1 gpc253 (
      {stage0_3[169]},
      {stage1_3[66]}
   );
   gpc1_1 gpc254 (
      {stage0_3[170]},
      {stage1_3[67]}
   );
   gpc1_1 gpc255 (
      {stage0_3[171]},
      {stage1_3[68]}
   );
   gpc1_1 gpc256 (
      {stage0_3[172]},
      {stage1_3[69]}
   );
   gpc1_1 gpc257 (
      {stage0_3[173]},
      {stage1_3[70]}
   );
   gpc1_1 gpc258 (
      {stage0_3[174]},
      {stage1_3[71]}
   );
   gpc1_1 gpc259 (
      {stage0_3[175]},
      {stage1_3[72]}
   );
   gpc1_1 gpc260 (
      {stage0_3[176]},
      {stage1_3[73]}
   );
   gpc1_1 gpc261 (
      {stage0_3[177]},
      {stage1_3[74]}
   );
   gpc1_1 gpc262 (
      {stage0_3[178]},
      {stage1_3[75]}
   );
   gpc1_1 gpc263 (
      {stage0_3[179]},
      {stage1_3[76]}
   );
   gpc1_1 gpc264 (
      {stage0_3[180]},
      {stage1_3[77]}
   );
   gpc1_1 gpc265 (
      {stage0_3[181]},
      {stage1_3[78]}
   );
   gpc1_1 gpc266 (
      {stage0_3[182]},
      {stage1_3[79]}
   );
   gpc1_1 gpc267 (
      {stage0_3[183]},
      {stage1_3[80]}
   );
   gpc1_1 gpc268 (
      {stage0_3[184]},
      {stage1_3[81]}
   );
   gpc1_1 gpc269 (
      {stage0_5[132]},
      {stage1_5[77]}
   );
   gpc1_1 gpc270 (
      {stage0_5[133]},
      {stage1_5[78]}
   );
   gpc1_1 gpc271 (
      {stage0_5[134]},
      {stage1_5[79]}
   );
   gpc1_1 gpc272 (
      {stage0_5[135]},
      {stage1_5[80]}
   );
   gpc1_1 gpc273 (
      {stage0_5[136]},
      {stage1_5[81]}
   );
   gpc1_1 gpc274 (
      {stage0_5[137]},
      {stage1_5[82]}
   );
   gpc1_1 gpc275 (
      {stage0_5[138]},
      {stage1_5[83]}
   );
   gpc1_1 gpc276 (
      {stage0_5[139]},
      {stage1_5[84]}
   );
   gpc1_1 gpc277 (
      {stage0_5[140]},
      {stage1_5[85]}
   );
   gpc1_1 gpc278 (
      {stage0_5[141]},
      {stage1_5[86]}
   );
   gpc1_1 gpc279 (
      {stage0_5[142]},
      {stage1_5[87]}
   );
   gpc1_1 gpc280 (
      {stage0_5[143]},
      {stage1_5[88]}
   );
   gpc1_1 gpc281 (
      {stage0_5[144]},
      {stage1_5[89]}
   );
   gpc1_1 gpc282 (
      {stage0_5[145]},
      {stage1_5[90]}
   );
   gpc1_1 gpc283 (
      {stage0_5[146]},
      {stage1_5[91]}
   );
   gpc1_1 gpc284 (
      {stage0_5[147]},
      {stage1_5[92]}
   );
   gpc1_1 gpc285 (
      {stage0_5[148]},
      {stage1_5[93]}
   );
   gpc1_1 gpc286 (
      {stage0_5[149]},
      {stage1_5[94]}
   );
   gpc1_1 gpc287 (
      {stage0_5[150]},
      {stage1_5[95]}
   );
   gpc1_1 gpc288 (
      {stage0_5[151]},
      {stage1_5[96]}
   );
   gpc1_1 gpc289 (
      {stage0_5[152]},
      {stage1_5[97]}
   );
   gpc1_1 gpc290 (
      {stage0_5[153]},
      {stage1_5[98]}
   );
   gpc1_1 gpc291 (
      {stage0_5[154]},
      {stage1_5[99]}
   );
   gpc1_1 gpc292 (
      {stage0_5[155]},
      {stage1_5[100]}
   );
   gpc1_1 gpc293 (
      {stage0_5[156]},
      {stage1_5[101]}
   );
   gpc1_1 gpc294 (
      {stage0_5[157]},
      {stage1_5[102]}
   );
   gpc1_1 gpc295 (
      {stage0_5[158]},
      {stage1_5[103]}
   );
   gpc1_1 gpc296 (
      {stage0_5[159]},
      {stage1_5[104]}
   );
   gpc1_1 gpc297 (
      {stage0_5[160]},
      {stage1_5[105]}
   );
   gpc1_1 gpc298 (
      {stage0_5[161]},
      {stage1_5[106]}
   );
   gpc1_1 gpc299 (
      {stage0_5[162]},
      {stage1_5[107]}
   );
   gpc1_1 gpc300 (
      {stage0_5[163]},
      {stage1_5[108]}
   );
   gpc1_1 gpc301 (
      {stage0_5[164]},
      {stage1_5[109]}
   );
   gpc1_1 gpc302 (
      {stage0_5[165]},
      {stage1_5[110]}
   );
   gpc1_1 gpc303 (
      {stage0_5[166]},
      {stage1_5[111]}
   );
   gpc1_1 gpc304 (
      {stage0_5[167]},
      {stage1_5[112]}
   );
   gpc1_1 gpc305 (
      {stage0_5[168]},
      {stage1_5[113]}
   );
   gpc1_1 gpc306 (
      {stage0_5[169]},
      {stage1_5[114]}
   );
   gpc1_1 gpc307 (
      {stage0_5[170]},
      {stage1_5[115]}
   );
   gpc1_1 gpc308 (
      {stage0_5[171]},
      {stage1_5[116]}
   );
   gpc1_1 gpc309 (
      {stage0_5[172]},
      {stage1_5[117]}
   );
   gpc1_1 gpc310 (
      {stage0_5[173]},
      {stage1_5[118]}
   );
   gpc1_1 gpc311 (
      {stage0_5[174]},
      {stage1_5[119]}
   );
   gpc1_1 gpc312 (
      {stage0_5[175]},
      {stage1_5[120]}
   );
   gpc1_1 gpc313 (
      {stage0_5[176]},
      {stage1_5[121]}
   );
   gpc1_1 gpc314 (
      {stage0_5[177]},
      {stage1_5[122]}
   );
   gpc1_1 gpc315 (
      {stage0_5[178]},
      {stage1_5[123]}
   );
   gpc1_1 gpc316 (
      {stage0_5[179]},
      {stage1_5[124]}
   );
   gpc1_1 gpc317 (
      {stage0_5[180]},
      {stage1_5[125]}
   );
   gpc1_1 gpc318 (
      {stage0_5[181]},
      {stage1_5[126]}
   );
   gpc1_1 gpc319 (
      {stage0_5[182]},
      {stage1_5[127]}
   );
   gpc1_1 gpc320 (
      {stage0_5[183]},
      {stage1_5[128]}
   );
   gpc1_1 gpc321 (
      {stage0_5[184]},
      {stage1_5[129]}
   );
   gpc1_1 gpc322 (
      {stage0_7[150]},
      {stage1_7[55]}
   );
   gpc1_1 gpc323 (
      {stage0_7[151]},
      {stage1_7[56]}
   );
   gpc1_1 gpc324 (
      {stage0_7[152]},
      {stage1_7[57]}
   );
   gpc1_1 gpc325 (
      {stage0_7[153]},
      {stage1_7[58]}
   );
   gpc1_1 gpc326 (
      {stage0_7[154]},
      {stage1_7[59]}
   );
   gpc1_1 gpc327 (
      {stage0_7[155]},
      {stage1_7[60]}
   );
   gpc1_1 gpc328 (
      {stage0_7[156]},
      {stage1_7[61]}
   );
   gpc1_1 gpc329 (
      {stage0_7[157]},
      {stage1_7[62]}
   );
   gpc1_1 gpc330 (
      {stage0_7[158]},
      {stage1_7[63]}
   );
   gpc1_1 gpc331 (
      {stage0_7[159]},
      {stage1_7[64]}
   );
   gpc1_1 gpc332 (
      {stage0_7[160]},
      {stage1_7[65]}
   );
   gpc1_1 gpc333 (
      {stage0_7[161]},
      {stage1_7[66]}
   );
   gpc1_1 gpc334 (
      {stage0_7[162]},
      {stage1_7[67]}
   );
   gpc1_1 gpc335 (
      {stage0_7[163]},
      {stage1_7[68]}
   );
   gpc1_1 gpc336 (
      {stage0_7[164]},
      {stage1_7[69]}
   );
   gpc1_1 gpc337 (
      {stage0_7[165]},
      {stage1_7[70]}
   );
   gpc1_1 gpc338 (
      {stage0_7[166]},
      {stage1_7[71]}
   );
   gpc1_1 gpc339 (
      {stage0_7[167]},
      {stage1_7[72]}
   );
   gpc1_1 gpc340 (
      {stage0_7[168]},
      {stage1_7[73]}
   );
   gpc1_1 gpc341 (
      {stage0_7[169]},
      {stage1_7[74]}
   );
   gpc1_1 gpc342 (
      {stage0_7[170]},
      {stage1_7[75]}
   );
   gpc1_1 gpc343 (
      {stage0_7[171]},
      {stage1_7[76]}
   );
   gpc1_1 gpc344 (
      {stage0_7[172]},
      {stage1_7[77]}
   );
   gpc1_1 gpc345 (
      {stage0_7[173]},
      {stage1_7[78]}
   );
   gpc1_1 gpc346 (
      {stage0_7[174]},
      {stage1_7[79]}
   );
   gpc1_1 gpc347 (
      {stage0_7[175]},
      {stage1_7[80]}
   );
   gpc1_1 gpc348 (
      {stage0_7[176]},
      {stage1_7[81]}
   );
   gpc1_1 gpc349 (
      {stage0_7[177]},
      {stage1_7[82]}
   );
   gpc1_1 gpc350 (
      {stage0_7[178]},
      {stage1_7[83]}
   );
   gpc1_1 gpc351 (
      {stage0_7[179]},
      {stage1_7[84]}
   );
   gpc1_1 gpc352 (
      {stage0_7[180]},
      {stage1_7[85]}
   );
   gpc1_1 gpc353 (
      {stage0_7[181]},
      {stage1_7[86]}
   );
   gpc1_1 gpc354 (
      {stage0_7[182]},
      {stage1_7[87]}
   );
   gpc1_1 gpc355 (
      {stage0_7[183]},
      {stage1_7[88]}
   );
   gpc1_1 gpc356 (
      {stage0_7[184]},
      {stage1_7[89]}
   );
   gpc1_1 gpc357 (
      {stage0_8[183]},
      {stage1_8[79]}
   );
   gpc1_1 gpc358 (
      {stage0_8[184]},
      {stage1_8[80]}
   );
   gpc1_1 gpc359 (
      {stage0_10[154]},
      {stage1_10[63]}
   );
   gpc1_1 gpc360 (
      {stage0_10[155]},
      {stage1_10[64]}
   );
   gpc1_1 gpc361 (
      {stage0_10[156]},
      {stage1_10[65]}
   );
   gpc1_1 gpc362 (
      {stage0_10[157]},
      {stage1_10[66]}
   );
   gpc1_1 gpc363 (
      {stage0_10[158]},
      {stage1_10[67]}
   );
   gpc1_1 gpc364 (
      {stage0_10[159]},
      {stage1_10[68]}
   );
   gpc1_1 gpc365 (
      {stage0_10[160]},
      {stage1_10[69]}
   );
   gpc1_1 gpc366 (
      {stage0_10[161]},
      {stage1_10[70]}
   );
   gpc1_1 gpc367 (
      {stage0_10[162]},
      {stage1_10[71]}
   );
   gpc1_1 gpc368 (
      {stage0_10[163]},
      {stage1_10[72]}
   );
   gpc1_1 gpc369 (
      {stage0_10[164]},
      {stage1_10[73]}
   );
   gpc1_1 gpc370 (
      {stage0_10[165]},
      {stage1_10[74]}
   );
   gpc1_1 gpc371 (
      {stage0_10[166]},
      {stage1_10[75]}
   );
   gpc1_1 gpc372 (
      {stage0_10[167]},
      {stage1_10[76]}
   );
   gpc1_1 gpc373 (
      {stage0_10[168]},
      {stage1_10[77]}
   );
   gpc1_1 gpc374 (
      {stage0_10[169]},
      {stage1_10[78]}
   );
   gpc1_1 gpc375 (
      {stage0_10[170]},
      {stage1_10[79]}
   );
   gpc1_1 gpc376 (
      {stage0_10[171]},
      {stage1_10[80]}
   );
   gpc1_1 gpc377 (
      {stage0_10[172]},
      {stage1_10[81]}
   );
   gpc1_1 gpc378 (
      {stage0_10[173]},
      {stage1_10[82]}
   );
   gpc1_1 gpc379 (
      {stage0_10[174]},
      {stage1_10[83]}
   );
   gpc1_1 gpc380 (
      {stage0_10[175]},
      {stage1_10[84]}
   );
   gpc1_1 gpc381 (
      {stage0_10[176]},
      {stage1_10[85]}
   );
   gpc1_1 gpc382 (
      {stage0_10[177]},
      {stage1_10[86]}
   );
   gpc1_1 gpc383 (
      {stage0_10[178]},
      {stage1_10[87]}
   );
   gpc1_1 gpc384 (
      {stage0_10[179]},
      {stage1_10[88]}
   );
   gpc1_1 gpc385 (
      {stage0_10[180]},
      {stage1_10[89]}
   );
   gpc1_1 gpc386 (
      {stage0_10[181]},
      {stage1_10[90]}
   );
   gpc1_1 gpc387 (
      {stage0_10[182]},
      {stage1_10[91]}
   );
   gpc1_1 gpc388 (
      {stage0_10[183]},
      {stage1_10[92]}
   );
   gpc1_1 gpc389 (
      {stage0_10[184]},
      {stage1_10[93]}
   );
   gpc1_1 gpc390 (
      {stage0_12[163]},
      {stage1_12[83]}
   );
   gpc1_1 gpc391 (
      {stage0_12[164]},
      {stage1_12[84]}
   );
   gpc1_1 gpc392 (
      {stage0_12[165]},
      {stage1_12[85]}
   );
   gpc1_1 gpc393 (
      {stage0_12[166]},
      {stage1_12[86]}
   );
   gpc1_1 gpc394 (
      {stage0_12[167]},
      {stage1_12[87]}
   );
   gpc1_1 gpc395 (
      {stage0_12[168]},
      {stage1_12[88]}
   );
   gpc1_1 gpc396 (
      {stage0_12[169]},
      {stage1_12[89]}
   );
   gpc1_1 gpc397 (
      {stage0_12[170]},
      {stage1_12[90]}
   );
   gpc1_1 gpc398 (
      {stage0_12[171]},
      {stage1_12[91]}
   );
   gpc1_1 gpc399 (
      {stage0_12[172]},
      {stage1_12[92]}
   );
   gpc1_1 gpc400 (
      {stage0_12[173]},
      {stage1_12[93]}
   );
   gpc1_1 gpc401 (
      {stage0_12[174]},
      {stage1_12[94]}
   );
   gpc1_1 gpc402 (
      {stage0_12[175]},
      {stage1_12[95]}
   );
   gpc1_1 gpc403 (
      {stage0_12[176]},
      {stage1_12[96]}
   );
   gpc1_1 gpc404 (
      {stage0_12[177]},
      {stage1_12[97]}
   );
   gpc1_1 gpc405 (
      {stage0_12[178]},
      {stage1_12[98]}
   );
   gpc1_1 gpc406 (
      {stage0_12[179]},
      {stage1_12[99]}
   );
   gpc1_1 gpc407 (
      {stage0_12[180]},
      {stage1_12[100]}
   );
   gpc1_1 gpc408 (
      {stage0_12[181]},
      {stage1_12[101]}
   );
   gpc1_1 gpc409 (
      {stage0_12[182]},
      {stage1_12[102]}
   );
   gpc1_1 gpc410 (
      {stage0_12[183]},
      {stage1_12[103]}
   );
   gpc1_1 gpc411 (
      {stage0_12[184]},
      {stage1_12[104]}
   );
   gpc1_1 gpc412 (
      {stage0_14[177]},
      {stage1_14[61]}
   );
   gpc1_1 gpc413 (
      {stage0_14[178]},
      {stage1_14[62]}
   );
   gpc1_1 gpc414 (
      {stage0_14[179]},
      {stage1_14[63]}
   );
   gpc1_1 gpc415 (
      {stage0_14[180]},
      {stage1_14[64]}
   );
   gpc1_1 gpc416 (
      {stage0_14[181]},
      {stage1_14[65]}
   );
   gpc1_1 gpc417 (
      {stage0_14[182]},
      {stage1_14[66]}
   );
   gpc1_1 gpc418 (
      {stage0_14[183]},
      {stage1_14[67]}
   );
   gpc1_1 gpc419 (
      {stage0_14[184]},
      {stage1_14[68]}
   );
   gpc1_1 gpc420 (
      {stage0_15[162]},
      {stage1_15[59]}
   );
   gpc1_1 gpc421 (
      {stage0_15[163]},
      {stage1_15[60]}
   );
   gpc1_1 gpc422 (
      {stage0_15[164]},
      {stage1_15[61]}
   );
   gpc1_1 gpc423 (
      {stage0_15[165]},
      {stage1_15[62]}
   );
   gpc1_1 gpc424 (
      {stage0_15[166]},
      {stage1_15[63]}
   );
   gpc1_1 gpc425 (
      {stage0_15[167]},
      {stage1_15[64]}
   );
   gpc1_1 gpc426 (
      {stage0_15[168]},
      {stage1_15[65]}
   );
   gpc1_1 gpc427 (
      {stage0_15[169]},
      {stage1_15[66]}
   );
   gpc1_1 gpc428 (
      {stage0_15[170]},
      {stage1_15[67]}
   );
   gpc1_1 gpc429 (
      {stage0_15[171]},
      {stage1_15[68]}
   );
   gpc1_1 gpc430 (
      {stage0_15[172]},
      {stage1_15[69]}
   );
   gpc1_1 gpc431 (
      {stage0_15[173]},
      {stage1_15[70]}
   );
   gpc1_1 gpc432 (
      {stage0_15[174]},
      {stage1_15[71]}
   );
   gpc1_1 gpc433 (
      {stage0_15[175]},
      {stage1_15[72]}
   );
   gpc1_1 gpc434 (
      {stage0_15[176]},
      {stage1_15[73]}
   );
   gpc1_1 gpc435 (
      {stage0_15[177]},
      {stage1_15[74]}
   );
   gpc1_1 gpc436 (
      {stage0_15[178]},
      {stage1_15[75]}
   );
   gpc1_1 gpc437 (
      {stage0_15[179]},
      {stage1_15[76]}
   );
   gpc1_1 gpc438 (
      {stage0_15[180]},
      {stage1_15[77]}
   );
   gpc1_1 gpc439 (
      {stage0_15[181]},
      {stage1_15[78]}
   );
   gpc1_1 gpc440 (
      {stage0_15[182]},
      {stage1_15[79]}
   );
   gpc1_1 gpc441 (
      {stage0_15[183]},
      {stage1_15[80]}
   );
   gpc1_1 gpc442 (
      {stage0_15[184]},
      {stage1_15[81]}
   );
   gpc1163_5 gpc443 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc444 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc445 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc446 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc447 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc448 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc449 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc450 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc451 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc452 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc453 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc454 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1343_5 gpc455 (
      {stage1_2[32], stage1_2[33], stage1_2[34]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[0], stage1_4[1], stage1_4[2]},
      {stage1_5[0]},
      {stage2_6[0],stage2_5[0],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc456 (
      {stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage1_3[12]},
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage2_6[1],stage2_5[1],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc457 (
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage1_3[13]},
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage2_6[2],stage2_5[2],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc458 (
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_3[14]},
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage2_6[3],stage2_5[3],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc459 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage1_3[15]},
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage2_6[4],stage2_5[4],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc460 (
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_3[16]},
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage2_6[5],stage2_5[5],stage2_4[17],stage2_3[17],stage2_2[17]}
   );
   gpc615_5 gpc461 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[33]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[0],stage2_6[6],stage2_5[6],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc462 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[34]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[1],stage2_6[7],stage2_5[7],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc463 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[35]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[2],stage2_6[8],stage2_5[8],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc464 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[36]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[3],stage2_6[9],stage2_5[9],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc465 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[37]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[4],stage2_6[10],stage2_5[10],stage2_4[22],stage2_3[22]}
   );
   gpc615_5 gpc466 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[38]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[5],stage2_6[11],stage2_5[11],stage2_4[23],stage2_3[23]}
   );
   gpc615_5 gpc467 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[39]},
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage2_7[6],stage2_6[12],stage2_5[12],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc468 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[40]},
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage2_7[7],stage2_6[13],stage2_5[13],stage2_4[25],stage2_3[25]}
   );
   gpc615_5 gpc469 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[41]},
      {stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54]},
      {stage2_7[8],stage2_6[14],stage2_5[14],stage2_4[26],stage2_3[26]}
   );
   gpc615_5 gpc470 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[42]},
      {stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60]},
      {stage2_7[9],stage2_6[15],stage2_5[15],stage2_4[27],stage2_3[27]}
   );
   gpc615_5 gpc471 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[43]},
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage2_7[10],stage2_6[16],stage2_5[16],stage2_4[28],stage2_3[28]}
   );
   gpc615_5 gpc472 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[44]},
      {stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72]},
      {stage2_7[11],stage2_6[17],stage2_5[17],stage2_4[29],stage2_3[29]}
   );
   gpc615_5 gpc473 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[45]},
      {stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78]},
      {stage2_7[12],stage2_6[18],stage2_5[18],stage2_4[30],stage2_3[30]}
   );
   gpc606_5 gpc474 (
      {stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[13],stage2_6[19],stage2_5[19],stage2_4[31]}
   );
   gpc606_5 gpc475 (
      {stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[14],stage2_6[20],stage2_5[20],stage2_4[32]}
   );
   gpc606_5 gpc476 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[15],stage2_6[21],stage2_5[21],stage2_4[33]}
   );
   gpc606_5 gpc477 (
      {stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[16],stage2_6[22],stage2_5[22],stage2_4[34]}
   );
   gpc615_5 gpc478 (
      {stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_5[79]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[17],stage2_6[23],stage2_5[23],stage2_4[35]}
   );
   gpc615_5 gpc479 (
      {stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79]},
      {stage1_5[80]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[18],stage2_6[24],stage2_5[24],stage2_4[36]}
   );
   gpc615_5 gpc480 (
      {stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84]},
      {stage1_5[81]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[19],stage2_6[25],stage2_5[25],stage2_4[37]}
   );
   gpc606_5 gpc481 (
      {stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[7],stage2_7[20],stage2_6[26],stage2_5[26]}
   );
   gpc606_5 gpc482 (
      {stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[8],stage2_7[21],stage2_6[27],stage2_5[27]}
   );
   gpc606_5 gpc483 (
      {stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[9],stage2_7[22],stage2_6[28],stage2_5[28]}
   );
   gpc606_5 gpc484 (
      {stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[10],stage2_7[23],stage2_6[29],stage2_5[29]}
   );
   gpc606_5 gpc485 (
      {stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[11],stage2_7[24],stage2_6[30],stage2_5[30]}
   );
   gpc606_5 gpc486 (
      {stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[12],stage2_7[25],stage2_6[31],stage2_5[31]}
   );
   gpc606_5 gpc487 (
      {stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[13],stage2_7[26],stage2_6[32],stage2_5[32]}
   );
   gpc606_5 gpc488 (
      {stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[14],stage2_7[27],stage2_6[33],stage2_5[33]}
   );
   gpc606_5 gpc489 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[15],stage2_7[28],stage2_6[34]}
   );
   gpc606_5 gpc490 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[16],stage2_7[29],stage2_6[35]}
   );
   gpc615_5 gpc491 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58]},
      {stage1_7[48]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[17],stage2_7[30],stage2_6[36]}
   );
   gpc615_5 gpc492 (
      {stage1_6[59], stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63]},
      {stage1_7[49]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[18],stage2_7[31],stage2_6[37]}
   );
   gpc615_5 gpc493 (
      {stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage1_8[24]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[4],stage2_9[12],stage2_8[19],stage2_7[32]}
   );
   gpc615_5 gpc494 (
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage1_8[25]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[5],stage2_9[13],stage2_8[20],stage2_7[33]}
   );
   gpc615_5 gpc495 (
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64]},
      {stage1_8[26]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[6],stage2_9[14],stage2_8[21],stage2_7[34]}
   );
   gpc615_5 gpc496 (
      {stage1_7[65], stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69]},
      {stage1_8[27]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[7],stage2_9[15],stage2_8[22],stage2_7[35]}
   );
   gpc615_5 gpc497 (
      {stage1_7[70], stage1_7[71], stage1_7[72], stage1_7[73], stage1_7[74]},
      {stage1_8[28]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[8],stage2_9[16],stage2_8[23],stage2_7[36]}
   );
   gpc615_5 gpc498 (
      {stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78], stage1_7[79]},
      {stage1_8[29]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[9],stage2_9[17],stage2_8[24],stage2_7[37]}
   );
   gpc615_5 gpc499 (
      {stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84]},
      {stage1_8[30]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[10],stage2_9[18],stage2_8[25],stage2_7[38]}
   );
   gpc615_5 gpc500 (
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage1_8[31]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[11],stage2_9[19],stage2_8[26],stage2_7[39]}
   );
   gpc606_5 gpc501 (
      {stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[8],stage2_10[12],stage2_9[20],stage2_8[27]}
   );
   gpc606_5 gpc502 (
      {stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[9],stage2_10[13],stage2_9[21],stage2_8[28]}
   );
   gpc606_5 gpc503 (
      {stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[10],stage2_10[14],stage2_9[22],stage2_8[29]}
   );
   gpc606_5 gpc504 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[11],stage2_10[15],stage2_9[23],stage2_8[30]}
   );
   gpc606_5 gpc505 (
      {stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[12],stage2_10[16],stage2_9[24],stage2_8[31]}
   );
   gpc606_5 gpc506 (
      {stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[13],stage2_10[17],stage2_9[25],stage2_8[32]}
   );
   gpc606_5 gpc507 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[6],stage2_11[14],stage2_10[18],stage2_9[26]}
   );
   gpc606_5 gpc508 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[7],stage2_11[15],stage2_10[19],stage2_9[27]}
   );
   gpc606_5 gpc509 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[8],stage2_11[16],stage2_10[20],stage2_9[28]}
   );
   gpc606_5 gpc510 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[9],stage2_11[17],stage2_10[21],stage2_9[29]}
   );
   gpc606_5 gpc511 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[10],stage2_11[18],stage2_10[22],stage2_9[30]}
   );
   gpc606_5 gpc512 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[11],stage2_11[19],stage2_10[23],stage2_9[31]}
   );
   gpc606_5 gpc513 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[6],stage2_12[12],stage2_11[20],stage2_10[24]}
   );
   gpc606_5 gpc514 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[7],stage2_12[13],stage2_11[21],stage2_10[25]}
   );
   gpc615_5 gpc515 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52]},
      {stage1_11[36]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[8],stage2_12[14],stage2_11[22],stage2_10[26]}
   );
   gpc615_5 gpc516 (
      {stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57]},
      {stage1_11[37]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[9],stage2_12[15],stage2_11[23],stage2_10[27]}
   );
   gpc615_5 gpc517 (
      {stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62]},
      {stage1_11[38]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[10],stage2_12[16],stage2_11[24],stage2_10[28]}
   );
   gpc615_5 gpc518 (
      {stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67]},
      {stage1_11[39]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[11],stage2_12[17],stage2_11[25],stage2_10[29]}
   );
   gpc615_5 gpc519 (
      {stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72]},
      {stage1_11[40]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[12],stage2_12[18],stage2_11[26],stage2_10[30]}
   );
   gpc615_5 gpc520 (
      {stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage1_11[41]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[13],stage2_12[19],stage2_11[27],stage2_10[31]}
   );
   gpc615_5 gpc521 (
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82]},
      {stage1_11[42]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[14],stage2_12[20],stage2_11[28],stage2_10[32]}
   );
   gpc615_5 gpc522 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87]},
      {stage1_11[43]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[15],stage2_12[21],stage2_11[29],stage2_10[33]}
   );
   gpc615_5 gpc523 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[60]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[10],stage2_13[16],stage2_12[22],stage2_11[30]}
   );
   gpc615_5 gpc524 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[61]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[11],stage2_13[17],stage2_12[23],stage2_11[31]}
   );
   gpc615_5 gpc525 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[62]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[12],stage2_13[18],stage2_12[24],stage2_11[32]}
   );
   gpc606_5 gpc526 (
      {stage1_12[63], stage1_12[64], stage1_12[65], stage1_12[66], stage1_12[67], stage1_12[68]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[3],stage2_14[13],stage2_13[19],stage2_12[25]}
   );
   gpc606_5 gpc527 (
      {stage1_12[69], stage1_12[70], stage1_12[71], stage1_12[72], stage1_12[73], stage1_12[74]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[4],stage2_14[14],stage2_13[20],stage2_12[26]}
   );
   gpc606_5 gpc528 (
      {stage1_12[75], stage1_12[76], stage1_12[77], stage1_12[78], stage1_12[79], stage1_12[80]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[5],stage2_14[15],stage2_13[21],stage2_12[27]}
   );
   gpc606_5 gpc529 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[6],stage2_14[16],stage2_13[22]}
   );
   gpc606_5 gpc530 (
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[7],stage2_14[17],stage2_13[23]}
   );
   gpc606_5 gpc531 (
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[8],stage2_14[18],stage2_13[24]}
   );
   gpc606_5 gpc532 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[6],stage2_15[9],stage2_14[19],stage2_13[25]}
   );
   gpc606_5 gpc533 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[7],stage2_15[10],stage2_14[20],stage2_13[26]}
   );
   gpc606_5 gpc534 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[8],stage2_15[11],stage2_14[21],stage2_13[27]}
   );
   gpc606_5 gpc535 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[9],stage2_15[12],stage2_14[22],stage2_13[28]}
   );
   gpc606_5 gpc536 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[10],stage2_15[13],stage2_14[23],stage2_13[29]}
   );
   gpc606_5 gpc537 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[11],stage2_15[14],stage2_14[24],stage2_13[30]}
   );
   gpc606_5 gpc538 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[12],stage2_15[15],stage2_14[25],stage2_13[31]}
   );
   gpc606_5 gpc539 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[10],stage2_16[13],stage2_15[16],stage2_14[26]}
   );
   gpc606_5 gpc540 (
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[11],stage2_16[14],stage2_15[17],stage2_14[27]}
   );
   gpc606_5 gpc541 (
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[12],stage2_16[15],stage2_15[18],stage2_14[28]}
   );
   gpc606_5 gpc542 (
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[13],stage2_16[16],stage2_15[19],stage2_14[29]}
   );
   gpc606_5 gpc543 (
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[14],stage2_16[17],stage2_15[20],stage2_14[30]}
   );
   gpc606_5 gpc544 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[15],stage2_16[18],stage2_15[21],stage2_14[31]}
   );
   gpc606_5 gpc545 (
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[16],stage2_16[19],stage2_15[22],stage2_14[32]}
   );
   gpc606_5 gpc546 (
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[17],stage2_16[20],stage2_15[23],stage2_14[33]}
   );
   gpc606_5 gpc547 (
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[8],stage2_17[18],stage2_16[21],stage2_15[24]}
   );
   gpc606_5 gpc548 (
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[9],stage2_17[19],stage2_16[22],stage2_15[25]}
   );
   gpc615_5 gpc549 (
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76]},
      {stage1_16[48]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[10],stage2_17[20],stage2_16[23],stage2_15[26]}
   );
   gpc615_5 gpc550 (
      {stage1_15[77], stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81]},
      {stage1_16[49]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[11],stage2_17[21],stage2_16[24],stage2_15[27]}
   );
   gpc1_1 gpc551 (
      {stage1_0[48]},
      {stage2_0[12]}
   );
   gpc1_1 gpc552 (
      {stage1_1[48]},
      {stage2_1[12]}
   );
   gpc1_1 gpc553 (
      {stage1_1[49]},
      {stage2_1[13]}
   );
   gpc1_1 gpc554 (
      {stage1_1[50]},
      {stage2_1[14]}
   );
   gpc1_1 gpc555 (
      {stage1_1[51]},
      {stage2_1[15]}
   );
   gpc1_1 gpc556 (
      {stage1_1[52]},
      {stage2_1[16]}
   );
   gpc1_1 gpc557 (
      {stage1_1[53]},
      {stage2_1[17]}
   );
   gpc1_1 gpc558 (
      {stage1_1[54]},
      {stage2_1[18]}
   );
   gpc1_1 gpc559 (
      {stage1_1[55]},
      {stage2_1[19]}
   );
   gpc1_1 gpc560 (
      {stage1_2[60]},
      {stage2_2[18]}
   );
   gpc1_1 gpc561 (
      {stage1_2[61]},
      {stage2_2[19]}
   );
   gpc1_1 gpc562 (
      {stage1_2[62]},
      {stage2_2[20]}
   );
   gpc1_1 gpc563 (
      {stage1_2[63]},
      {stage2_2[21]}
   );
   gpc1_1 gpc564 (
      {stage1_2[64]},
      {stage2_2[22]}
   );
   gpc1_1 gpc565 (
      {stage1_2[65]},
      {stage2_2[23]}
   );
   gpc1_1 gpc566 (
      {stage1_2[66]},
      {stage2_2[24]}
   );
   gpc1_1 gpc567 (
      {stage1_8[68]},
      {stage2_8[33]}
   );
   gpc1_1 gpc568 (
      {stage1_8[69]},
      {stage2_8[34]}
   );
   gpc1_1 gpc569 (
      {stage1_8[70]},
      {stage2_8[35]}
   );
   gpc1_1 gpc570 (
      {stage1_8[71]},
      {stage2_8[36]}
   );
   gpc1_1 gpc571 (
      {stage1_8[72]},
      {stage2_8[37]}
   );
   gpc1_1 gpc572 (
      {stage1_8[73]},
      {stage2_8[38]}
   );
   gpc1_1 gpc573 (
      {stage1_8[74]},
      {stage2_8[39]}
   );
   gpc1_1 gpc574 (
      {stage1_8[75]},
      {stage2_8[40]}
   );
   gpc1_1 gpc575 (
      {stage1_8[76]},
      {stage2_8[41]}
   );
   gpc1_1 gpc576 (
      {stage1_8[77]},
      {stage2_8[42]}
   );
   gpc1_1 gpc577 (
      {stage1_8[78]},
      {stage2_8[43]}
   );
   gpc1_1 gpc578 (
      {stage1_8[79]},
      {stage2_8[44]}
   );
   gpc1_1 gpc579 (
      {stage1_8[80]},
      {stage2_8[45]}
   );
   gpc1_1 gpc580 (
      {stage1_10[88]},
      {stage2_10[34]}
   );
   gpc1_1 gpc581 (
      {stage1_10[89]},
      {stage2_10[35]}
   );
   gpc1_1 gpc582 (
      {stage1_10[90]},
      {stage2_10[36]}
   );
   gpc1_1 gpc583 (
      {stage1_10[91]},
      {stage2_10[37]}
   );
   gpc1_1 gpc584 (
      {stage1_10[92]},
      {stage2_10[38]}
   );
   gpc1_1 gpc585 (
      {stage1_10[93]},
      {stage2_10[39]}
   );
   gpc1_1 gpc586 (
      {stage1_12[81]},
      {stage2_12[28]}
   );
   gpc1_1 gpc587 (
      {stage1_12[82]},
      {stage2_12[29]}
   );
   gpc1_1 gpc588 (
      {stage1_12[83]},
      {stage2_12[30]}
   );
   gpc1_1 gpc589 (
      {stage1_12[84]},
      {stage2_12[31]}
   );
   gpc1_1 gpc590 (
      {stage1_12[85]},
      {stage2_12[32]}
   );
   gpc1_1 gpc591 (
      {stage1_12[86]},
      {stage2_12[33]}
   );
   gpc1_1 gpc592 (
      {stage1_12[87]},
      {stage2_12[34]}
   );
   gpc1_1 gpc593 (
      {stage1_12[88]},
      {stage2_12[35]}
   );
   gpc1_1 gpc594 (
      {stage1_12[89]},
      {stage2_12[36]}
   );
   gpc1_1 gpc595 (
      {stage1_12[90]},
      {stage2_12[37]}
   );
   gpc1_1 gpc596 (
      {stage1_12[91]},
      {stage2_12[38]}
   );
   gpc1_1 gpc597 (
      {stage1_12[92]},
      {stage2_12[39]}
   );
   gpc1_1 gpc598 (
      {stage1_12[93]},
      {stage2_12[40]}
   );
   gpc1_1 gpc599 (
      {stage1_12[94]},
      {stage2_12[41]}
   );
   gpc1_1 gpc600 (
      {stage1_12[95]},
      {stage2_12[42]}
   );
   gpc1_1 gpc601 (
      {stage1_12[96]},
      {stage2_12[43]}
   );
   gpc1_1 gpc602 (
      {stage1_12[97]},
      {stage2_12[44]}
   );
   gpc1_1 gpc603 (
      {stage1_12[98]},
      {stage2_12[45]}
   );
   gpc1_1 gpc604 (
      {stage1_12[99]},
      {stage2_12[46]}
   );
   gpc1_1 gpc605 (
      {stage1_12[100]},
      {stage2_12[47]}
   );
   gpc1_1 gpc606 (
      {stage1_12[101]},
      {stage2_12[48]}
   );
   gpc1_1 gpc607 (
      {stage1_12[102]},
      {stage2_12[49]}
   );
   gpc1_1 gpc608 (
      {stage1_12[103]},
      {stage2_12[50]}
   );
   gpc1_1 gpc609 (
      {stage1_12[104]},
      {stage2_12[51]}
   );
   gpc1_1 gpc610 (
      {stage1_13[78]},
      {stage2_13[32]}
   );
   gpc1_1 gpc611 (
      {stage1_13[79]},
      {stage2_13[33]}
   );
   gpc1_1 gpc612 (
      {stage1_13[80]},
      {stage2_13[34]}
   );
   gpc1_1 gpc613 (
      {stage1_13[81]},
      {stage2_13[35]}
   );
   gpc1_1 gpc614 (
      {stage1_13[82]},
      {stage2_13[36]}
   );
   gpc1_1 gpc615 (
      {stage1_13[83]},
      {stage2_13[37]}
   );
   gpc1_1 gpc616 (
      {stage1_13[84]},
      {stage2_13[38]}
   );
   gpc1_1 gpc617 (
      {stage1_13[85]},
      {stage2_13[39]}
   );
   gpc1_1 gpc618 (
      {stage1_14[66]},
      {stage2_14[34]}
   );
   gpc1_1 gpc619 (
      {stage1_14[67]},
      {stage2_14[35]}
   );
   gpc1_1 gpc620 (
      {stage1_14[68]},
      {stage2_14[36]}
   );
   gpc1_1 gpc621 (
      {stage1_16[50]},
      {stage2_16[25]}
   );
   gpc1_1 gpc622 (
      {stage1_16[51]},
      {stage2_16[26]}
   );
   gpc1_1 gpc623 (
      {stage1_16[52]},
      {stage2_16[27]}
   );
   gpc1_1 gpc624 (
      {stage1_17[24]},
      {stage2_17[22]}
   );
   gpc1_1 gpc625 (
      {stage1_17[25]},
      {stage2_17[23]}
   );
   gpc1_1 gpc626 (
      {stage1_17[26]},
      {stage2_17[24]}
   );
   gpc1163_5 gpc627 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc628 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7]},
      {stage2_1[6]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc629 (
      {stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11], stage2_1[12]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc630 (
      {stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17], stage2_1[18]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc631 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc632 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage2_3[13]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[3],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc1163_5 gpc633 (
      {stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc1163_5 gpc634 (
      {stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[5],stage3_4[7],stage3_3[7]}
   );
   gpc615_5 gpc635 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage2_4[24]},
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage3_7[2],stage3_6[4],stage3_5[6],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc636 (
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage2_4[25]},
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12], stage2_5[13]},
      {stage3_7[3],stage3_6[5],stage3_5[7],stage3_4[9],stage3_3[9]}
   );
   gpc606_5 gpc637 (
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7]},
      {stage3_8[0],stage3_7[4],stage3_6[6],stage3_5[8],stage3_4[10]}
   );
   gpc606_5 gpc638 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13]},
      {stage3_8[1],stage3_7[5],stage3_6[7],stage3_5[9],stage3_4[11]}
   );
   gpc606_5 gpc639 (
      {stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18], stage2_5[19]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[6],stage3_6[8],stage3_5[10]}
   );
   gpc606_5 gpc640 (
      {stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24], stage2_5[25]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[7],stage3_6[9],stage3_5[11]}
   );
   gpc606_5 gpc641 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[4],stage3_7[8],stage3_6[10],stage3_5[12]}
   );
   gpc606_5 gpc642 (
      {stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[5],stage3_7[9],stage3_6[11]}
   );
   gpc606_5 gpc643 (
      {stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[4],stage3_8[6],stage3_7[10],stage3_6[12]}
   );
   gpc606_5 gpc644 (
      {stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30], stage2_6[31]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[5],stage3_8[7],stage3_7[11],stage3_6[13]}
   );
   gpc615_5 gpc645 (
      {stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35], stage2_6[36]},
      {stage2_7[18]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[6],stage3_8[8],stage3_7[12],stage3_6[14]}
   );
   gpc615_5 gpc646 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[24]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[4],stage3_9[7],stage3_8[9],stage3_7[13]}
   );
   gpc615_5 gpc647 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[25]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[5],stage3_9[8],stage3_8[10],stage3_7[14]}
   );
   gpc615_5 gpc648 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[26]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[6],stage3_9[9],stage3_8[11],stage3_7[15]}
   );
   gpc615_5 gpc649 (
      {stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31]},
      {stage2_9[18]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[3],stage3_10[7],stage3_9[10],stage3_8[12]}
   );
   gpc615_5 gpc650 (
      {stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_9[19]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[4],stage3_10[8],stage3_9[11],stage3_8[13]}
   );
   gpc615_5 gpc651 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage2_9[20]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[5],stage3_10[9],stage3_9[12],stage3_8[14]}
   );
   gpc606_5 gpc652 (
      {stage2_9[21], stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[6],stage3_10[10],stage3_9[13]}
   );
   gpc615_5 gpc653 (
      {stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30], stage2_9[31]},
      {stage2_10[18]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[7],stage3_10[11],stage3_9[14]}
   );
   gpc615_5 gpc654 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[12]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[2],stage3_12[5],stage3_11[8],stage3_10[12]}
   );
   gpc615_5 gpc655 (
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28]},
      {stage2_11[13]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[3],stage3_12[6],stage3_11[9],stage3_10[13]}
   );
   gpc615_5 gpc656 (
      {stage2_10[29], stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33]},
      {stage2_11[14]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[4],stage3_12[7],stage3_11[10],stage3_10[14]}
   );
   gpc615_5 gpc657 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[5],stage3_12[8],stage3_11[11]}
   );
   gpc615_5 gpc658 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[6],stage3_12[9],stage3_11[12]}
   );
   gpc615_5 gpc659 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_12[20]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[7],stage3_12[10],stage3_11[13]}
   );
   gpc606_5 gpc660 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[6],stage3_13[8],stage3_12[11]}
   );
   gpc606_5 gpc661 (
      {stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31], stage2_12[32]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[4],stage3_14[7],stage3_13[9],stage3_12[12]}
   );
   gpc606_5 gpc662 (
      {stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37], stage2_12[38]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[5],stage3_14[8],stage3_13[10],stage3_12[13]}
   );
   gpc606_5 gpc663 (
      {stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43], stage2_12[44]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[6],stage3_14[9],stage3_13[11],stage3_12[14]}
   );
   gpc606_5 gpc664 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[7],stage3_14[10],stage3_13[12]}
   );
   gpc606_5 gpc665 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[5],stage3_15[8],stage3_14[11],stage3_13[13]}
   );
   gpc606_5 gpc666 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[6],stage3_15[9],stage3_14[12],stage3_13[14]}
   );
   gpc606_5 gpc667 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[7],stage3_15[10],stage3_14[13]}
   );
   gpc606_5 gpc668 (
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[4],stage3_16[8],stage3_15[11],stage3_14[14]}
   );
   gpc615_5 gpc669 (
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22]},
      {stage2_16[12]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[5],stage3_16[9],stage3_15[12]}
   );
   gpc615_5 gpc670 (
      {stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_16[13]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[3],stage3_17[6],stage3_16[10],stage3_15[13]}
   );
   gpc606_5 gpc671 (
      {stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17], stage2_16[18], stage2_16[19]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[4],stage3_17[7],stage3_16[11]}
   );
   gpc606_5 gpc672 (
      {stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23], stage2_16[24], stage2_16[25]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[3],stage3_18[5],stage3_17[8],stage3_16[12]}
   );
   gpc1_1 gpc673 (
      {stage2_0[8]},
      {stage3_0[2]}
   );
   gpc1_1 gpc674 (
      {stage2_0[9]},
      {stage3_0[3]}
   );
   gpc1_1 gpc675 (
      {stage2_0[10]},
      {stage3_0[4]}
   );
   gpc1_1 gpc676 (
      {stage2_0[11]},
      {stage3_0[5]}
   );
   gpc1_1 gpc677 (
      {stage2_0[12]},
      {stage3_0[6]}
   );
   gpc1_1 gpc678 (
      {stage2_1[19]},
      {stage3_1[4]}
   );
   gpc1_1 gpc679 (
      {stage2_2[18]},
      {stage3_2[6]}
   );
   gpc1_1 gpc680 (
      {stage2_2[19]},
      {stage3_2[7]}
   );
   gpc1_1 gpc681 (
      {stage2_2[20]},
      {stage3_2[8]}
   );
   gpc1_1 gpc682 (
      {stage2_2[21]},
      {stage3_2[9]}
   );
   gpc1_1 gpc683 (
      {stage2_2[22]},
      {stage3_2[10]}
   );
   gpc1_1 gpc684 (
      {stage2_2[23]},
      {stage3_2[11]}
   );
   gpc1_1 gpc685 (
      {stage2_2[24]},
      {stage3_2[12]}
   );
   gpc1_1 gpc686 (
      {stage2_3[30]},
      {stage3_3[10]}
   );
   gpc1_1 gpc687 (
      {stage2_5[32]},
      {stage3_5[13]}
   );
   gpc1_1 gpc688 (
      {stage2_5[33]},
      {stage3_5[14]}
   );
   gpc1_1 gpc689 (
      {stage2_6[37]},
      {stage3_6[15]}
   );
   gpc1_1 gpc690 (
      {stage2_7[34]},
      {stage3_7[16]}
   );
   gpc1_1 gpc691 (
      {stage2_7[35]},
      {stage3_7[17]}
   );
   gpc1_1 gpc692 (
      {stage2_7[36]},
      {stage3_7[18]}
   );
   gpc1_1 gpc693 (
      {stage2_7[37]},
      {stage3_7[19]}
   );
   gpc1_1 gpc694 (
      {stage2_7[38]},
      {stage3_7[20]}
   );
   gpc1_1 gpc695 (
      {stage2_7[39]},
      {stage3_7[21]}
   );
   gpc1_1 gpc696 (
      {stage2_8[42]},
      {stage3_8[15]}
   );
   gpc1_1 gpc697 (
      {stage2_8[43]},
      {stage3_8[16]}
   );
   gpc1_1 gpc698 (
      {stage2_8[44]},
      {stage3_8[17]}
   );
   gpc1_1 gpc699 (
      {stage2_8[45]},
      {stage3_8[18]}
   );
   gpc1_1 gpc700 (
      {stage2_10[34]},
      {stage3_10[15]}
   );
   gpc1_1 gpc701 (
      {stage2_10[35]},
      {stage3_10[16]}
   );
   gpc1_1 gpc702 (
      {stage2_10[36]},
      {stage3_10[17]}
   );
   gpc1_1 gpc703 (
      {stage2_10[37]},
      {stage3_10[18]}
   );
   gpc1_1 gpc704 (
      {stage2_10[38]},
      {stage3_10[19]}
   );
   gpc1_1 gpc705 (
      {stage2_10[39]},
      {stage3_10[20]}
   );
   gpc1_1 gpc706 (
      {stage2_11[30]},
      {stage3_11[14]}
   );
   gpc1_1 gpc707 (
      {stage2_11[31]},
      {stage3_11[15]}
   );
   gpc1_1 gpc708 (
      {stage2_11[32]},
      {stage3_11[16]}
   );
   gpc1_1 gpc709 (
      {stage2_12[45]},
      {stage3_12[15]}
   );
   gpc1_1 gpc710 (
      {stage2_12[46]},
      {stage3_12[16]}
   );
   gpc1_1 gpc711 (
      {stage2_12[47]},
      {stage3_12[17]}
   );
   gpc1_1 gpc712 (
      {stage2_12[48]},
      {stage3_12[18]}
   );
   gpc1_1 gpc713 (
      {stage2_12[49]},
      {stage3_12[19]}
   );
   gpc1_1 gpc714 (
      {stage2_12[50]},
      {stage3_12[20]}
   );
   gpc1_1 gpc715 (
      {stage2_12[51]},
      {stage3_12[21]}
   );
   gpc1_1 gpc716 (
      {stage2_13[36]},
      {stage3_13[15]}
   );
   gpc1_1 gpc717 (
      {stage2_13[37]},
      {stage3_13[16]}
   );
   gpc1_1 gpc718 (
      {stage2_13[38]},
      {stage3_13[17]}
   );
   gpc1_1 gpc719 (
      {stage2_13[39]},
      {stage3_13[18]}
   );
   gpc1_1 gpc720 (
      {stage2_14[36]},
      {stage3_14[15]}
   );
   gpc1_1 gpc721 (
      {stage2_16[26]},
      {stage3_16[13]}
   );
   gpc1_1 gpc722 (
      {stage2_16[27]},
      {stage3_16[14]}
   );
   gpc1_1 gpc723 (
      {stage2_17[12]},
      {stage3_17[9]}
   );
   gpc1_1 gpc724 (
      {stage2_17[13]},
      {stage3_17[10]}
   );
   gpc1_1 gpc725 (
      {stage2_17[14]},
      {stage3_17[11]}
   );
   gpc1_1 gpc726 (
      {stage2_17[15]},
      {stage3_17[12]}
   );
   gpc1_1 gpc727 (
      {stage2_17[16]},
      {stage3_17[13]}
   );
   gpc1_1 gpc728 (
      {stage2_17[17]},
      {stage3_17[14]}
   );
   gpc1_1 gpc729 (
      {stage2_17[18]},
      {stage3_17[15]}
   );
   gpc1_1 gpc730 (
      {stage2_17[19]},
      {stage3_17[16]}
   );
   gpc1_1 gpc731 (
      {stage2_17[20]},
      {stage3_17[17]}
   );
   gpc1_1 gpc732 (
      {stage2_17[21]},
      {stage3_17[18]}
   );
   gpc1_1 gpc733 (
      {stage2_17[22]},
      {stage3_17[19]}
   );
   gpc1_1 gpc734 (
      {stage2_17[23]},
      {stage3_17[20]}
   );
   gpc1_1 gpc735 (
      {stage2_17[24]},
      {stage3_17[21]}
   );
   gpc1_1 gpc736 (
      {stage2_19[0]},
      {stage3_19[4]}
   );
   gpc1_1 gpc737 (
      {stage2_19[1]},
      {stage3_19[5]}
   );
   gpc1_1 gpc738 (
      {stage2_19[2]},
      {stage3_19[6]}
   );
   gpc1_1 gpc739 (
      {stage2_19[3]},
      {stage3_19[7]}
   );
   gpc606_5 gpc740 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc741 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc615_5 gpc742 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc743 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[6]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc744 (
      {stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[3],stage4_5[3]}
   );
   gpc615_5 gpc745 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[2],stage4_7[3],stage4_6[4]}
   );
   gpc615_5 gpc746 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[3],stage4_7[4],stage4_6[5]}
   );
   gpc615_5 gpc747 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12]},
      {stage3_8[12]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[2],stage4_9[3],stage4_8[4],stage4_7[5]}
   );
   gpc615_5 gpc748 (
      {stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage3_8[13]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[3],stage4_9[4],stage4_8[5],stage4_7[6]}
   );
   gpc615_5 gpc749 (
      {stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17], stage3_8[18]},
      {stage3_9[12]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[2],stage4_10[4],stage4_9[5],stage4_8[6]}
   );
   gpc2135_5 gpc750 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10]},
      {stage3_11[0], stage3_11[1], stage3_11[2]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[3],stage4_10[5]}
   );
   gpc615_5 gpc751 (
      {stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15]},
      {stage3_11[3]},
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage4_14[1],stage4_13[1],stage4_12[2],stage4_11[4],stage4_10[6]}
   );
   gpc615_5 gpc752 (
      {stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19], stage3_10[20]},
      {stage3_11[4]},
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage4_14[2],stage4_13[2],stage4_12[3],stage4_11[5],stage4_10[7]}
   );
   gpc615_5 gpc753 (
      {stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage3_12[13]},
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage4_15[0],stage4_14[3],stage4_13[3],stage4_12[4],stage4_11[6]}
   );
   gpc606_5 gpc754 (
      {stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18], stage3_12[19]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[4],stage4_13[4],stage4_12[5]}
   );
   gpc1325_5 gpc755 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12]},
      {stage3_14[6], stage3_14[7]},
      {stage3_15[0], stage3_15[1], stage3_15[2]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[5],stage4_13[5]}
   );
   gpc1325_5 gpc756 (
      {stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_14[8], stage3_14[9]},
      {stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage3_16[1]},
      {stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[6],stage4_13[6]}
   );
   gpc606_5 gpc757 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6], stage3_16[7]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[7]}
   );
   gpc1163_5 gpc758 (
      {stage3_15[6], stage3_15[7], stage3_15[8]},
      {stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[5]}
   );
   gpc615_5 gpc759 (
      {stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13]},
      {stage3_16[14]},
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage4_19[1],stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[6]}
   );
   gpc117_4 gpc760 (
      {stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11], stage3_17[12], stage3_17[13]},
      {stage3_18[1]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[2],stage4_18[3],stage4_17[5]}
   );
   gpc606_5 gpc761 (
      {stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17], stage3_17[18], stage3_17[19]},
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage4_21[0],stage4_20[1],stage4_19[3],stage4_18[4],stage4_17[6]}
   );
   gpc1_1 gpc762 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc763 (
      {stage3_1[0]},
      {stage4_1[1]}
   );
   gpc1_1 gpc764 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc765 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc766 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc767 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc768 (
      {stage3_2[11]},
      {stage4_2[2]}
   );
   gpc1_1 gpc769 (
      {stage3_2[12]},
      {stage4_2[3]}
   );
   gpc1_1 gpc770 (
      {stage3_3[6]},
      {stage4_3[3]}
   );
   gpc1_1 gpc771 (
      {stage3_3[7]},
      {stage4_3[4]}
   );
   gpc1_1 gpc772 (
      {stage3_3[8]},
      {stage4_3[5]}
   );
   gpc1_1 gpc773 (
      {stage3_3[9]},
      {stage4_3[6]}
   );
   gpc1_1 gpc774 (
      {stage3_3[10]},
      {stage4_3[7]}
   );
   gpc1_1 gpc775 (
      {stage3_5[13]},
      {stage4_5[4]}
   );
   gpc1_1 gpc776 (
      {stage3_5[14]},
      {stage4_5[5]}
   );
   gpc1_1 gpc777 (
      {stage3_7[18]},
      {stage4_7[7]}
   );
   gpc1_1 gpc778 (
      {stage3_7[19]},
      {stage4_7[8]}
   );
   gpc1_1 gpc779 (
      {stage3_7[20]},
      {stage4_7[9]}
   );
   gpc1_1 gpc780 (
      {stage3_7[21]},
      {stage4_7[10]}
   );
   gpc1_1 gpc781 (
      {stage3_9[13]},
      {stage4_9[6]}
   );
   gpc1_1 gpc782 (
      {stage3_9[14]},
      {stage4_9[7]}
   );
   gpc1_1 gpc783 (
      {stage3_11[10]},
      {stage4_11[7]}
   );
   gpc1_1 gpc784 (
      {stage3_11[11]},
      {stage4_11[8]}
   );
   gpc1_1 gpc785 (
      {stage3_11[12]},
      {stage4_11[9]}
   );
   gpc1_1 gpc786 (
      {stage3_11[13]},
      {stage4_11[10]}
   );
   gpc1_1 gpc787 (
      {stage3_11[14]},
      {stage4_11[11]}
   );
   gpc1_1 gpc788 (
      {stage3_11[15]},
      {stage4_11[12]}
   );
   gpc1_1 gpc789 (
      {stage3_11[16]},
      {stage4_11[13]}
   );
   gpc1_1 gpc790 (
      {stage3_12[20]},
      {stage4_12[6]}
   );
   gpc1_1 gpc791 (
      {stage3_12[21]},
      {stage4_12[7]}
   );
   gpc1_1 gpc792 (
      {stage3_13[18]},
      {stage4_13[7]}
   );
   gpc1_1 gpc793 (
      {stage3_17[20]},
      {stage4_17[7]}
   );
   gpc1_1 gpc794 (
      {stage3_17[21]},
      {stage4_17[8]}
   );
   gpc1_1 gpc795 (
      {stage3_18[2]},
      {stage4_18[5]}
   );
   gpc1_1 gpc796 (
      {stage3_18[3]},
      {stage4_18[6]}
   );
   gpc1_1 gpc797 (
      {stage3_18[4]},
      {stage4_18[7]}
   );
   gpc1_1 gpc798 (
      {stage3_18[5]},
      {stage4_18[8]}
   );
   gpc1_1 gpc799 (
      {stage3_19[7]},
      {stage4_19[4]}
   );
   gpc1_1 gpc800 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc1_1 gpc801 (
      {stage3_20[1]},
      {stage4_20[3]}
   );
   gpc2135_5 gpc802 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc7_3 gpc803 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6], stage4_3[7]},
      {stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1343_5 gpc804 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0], stage4_8[1], stage4_8[2]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0]}
   );
   gpc1343_5 gpc805 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc1343_5 gpc806 (
      {stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc1343_5 gpc807 (
      {stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3],stage5_9[3]}
   );
   gpc117_4 gpc808 (
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12]},
      {stage4_12[2]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[2]}
   );
   gpc15_3 gpc809 (
      {stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage4_13[1]},
      {stage5_14[1],stage5_13[3],stage5_12[3]}
   );
   gpc615_5 gpc810 (
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[4]}
   );
   gpc606_5 gpc811 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5], stage4_14[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[3]}
   );
   gpc2135_5 gpc812 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4]},
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1]},
      {stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[2]}
   );
   gpc2135_5 gpc813 (
      {stage4_17[5], stage4_17[6], stage4_17[7], stage4_17[8], 1'b0},
      {stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[1]},
      {stage4_20[2], stage4_20[3]},
      {stage5_21[1],stage5_20[1],stage5_19[1],stage5_18[2],stage5_17[3]}
   );
   gpc1163_5 gpc814 (
      {stage4_18[6], stage4_18[7], stage4_18[8]},
      {stage4_19[2], stage4_19[3], stage4_19[4], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[2],stage5_20[2],stage5_19[2],stage5_18[3]}
   );
   gpc1_1 gpc815 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc816 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc817 (
      {stage4_1[5]},
      {stage5_1[1]}
   );
   gpc1_1 gpc818 (
      {stage4_2[3]},
      {stage5_2[1]}
   );
   gpc1_1 gpc819 (
      {stage4_4[2]},
      {stage5_4[2]}
   );
   gpc1_1 gpc820 (
      {stage4_4[3]},
      {stage5_4[3]}
   );
   gpc1_1 gpc821 (
      {stage4_5[0]},
      {stage5_5[2]}
   );
   gpc1_1 gpc822 (
      {stage4_5[1]},
      {stage5_5[3]}
   );
   gpc1_1 gpc823 (
      {stage4_5[2]},
      {stage5_5[4]}
   );
   gpc1_1 gpc824 (
      {stage4_5[3]},
      {stage5_5[5]}
   );
   gpc1_1 gpc825 (
      {stage4_5[4]},
      {stage5_5[6]}
   );
   gpc1_1 gpc826 (
      {stage4_5[5]},
      {stage5_5[7]}
   );
   gpc1_1 gpc827 (
      {stage4_7[8]},
      {stage5_7[2]}
   );
   gpc1_1 gpc828 (
      {stage4_7[9]},
      {stage5_7[3]}
   );
   gpc1_1 gpc829 (
      {stage4_7[10]},
      {stage5_7[4]}
   );
   gpc1_1 gpc830 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc831 (
      {stage4_11[13]},
      {stage5_11[3]}
   );
   gpc1_1 gpc832 (
      {stage4_13[7]},
      {stage5_13[5]}
   );
   gpc1_1 gpc833 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc834 (
      {stage4_15[6]},
      {stage5_15[2]}
   );
   gpc223_4 gpc835 (
      {stage5_4[0], stage5_4[1], stage5_4[2]},
      {stage5_5[0], stage5_5[1]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0]}
   );
   gpc606_5 gpc836 (
      {stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5], stage5_5[6], stage5_5[7]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], 1'b0},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc837 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc1343_5 gpc838 (
      {stage5_11[1], stage5_11[2], stage5_11[3]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3]},
      {stage5_13[0], stage5_13[1], stage5_13[2]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1343_5 gpc839 (
      {stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc2135_5 gpc840 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], 1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2]},
      {stage5_19[0]},
      {stage5_20[0], stage5_20[1]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1]}
   );
   gpc1343_5 gpc841 (
      {stage5_19[1], stage5_19[2], 1'b0},
      {stage5_20[2], 1'b0, 1'b0, 1'b0},
      {stage5_21[0], stage5_21[1], stage5_21[2]},
      {stage5_22[0]},
      {stage6_23[0],stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1]}
   );
   gpc1_1 gpc842 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc843 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc844 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc845 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc846 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc847 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc848 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc849 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc850 (
      {stage5_4[3]},
      {stage6_4[1]}
   );
   gpc1_1 gpc851 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc852 (
      {stage5_16[1]},
      {stage6_16[1]}
   );
   gpc1_1 gpc853 (
      {stage5_18[3]},
      {stage6_18[1]}
   );
endmodule
module rowadder2_1_24(input [23:0] src0, input [23:0] src1, output [24:0] dst0);
    wire [23:0] gene;
    wire [23:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    assign dst0 = {carryout[23], out[23:0]};
endmodule


module comp2_1test_185_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    reg [15:0] src128;
    reg [15:0] src129;
    reg [15:0] src130;
    reg [15:0] src131;
    reg [15:0] src132;
    reg [15:0] src133;
    reg [15:0] src134;
    reg [15:0] src135;
    reg [15:0] src136;
    reg [15:0] src137;
    reg [15:0] src138;
    reg [15:0] src139;
    reg [15:0] src140;
    reg [15:0] src141;
    reg [15:0] src142;
    reg [15:0] src143;
    reg [15:0] src144;
    reg [15:0] src145;
    reg [15:0] src146;
    reg [15:0] src147;
    reg [15:0] src148;
    reg [15:0] src149;
    reg [15:0] src150;
    reg [15:0] src151;
    reg [15:0] src152;
    reg [15:0] src153;
    reg [15:0] src154;
    reg [15:0] src155;
    reg [15:0] src156;
    reg [15:0] src157;
    reg [15:0] src158;
    reg [15:0] src159;
    reg [15:0] src160;
    reg [15:0] src161;
    reg [15:0] src162;
    reg [15:0] src163;
    reg [15:0] src164;
    reg [15:0] src165;
    reg [15:0] src166;
    reg [15:0] src167;
    reg [15:0] src168;
    reg [15:0] src169;
    reg [15:0] src170;
    reg [15:0] src171;
    reg [15:0] src172;
    reg [15:0] src173;
    reg [15:0] src174;
    reg [15:0] src175;
    reg [15:0] src176;
    reg [15:0] src177;
    reg [15:0] src178;
    reg [15:0] src179;
    reg [15:0] src180;
    reg [15:0] src181;
    reg [15:0] src182;
    reg [15:0] src183;
    reg [15:0] src184;
    reg [23:0] exp;
    wire [23:0] dst;
    assign test = dst == exp;
    compressor2_1_185_16 compressor2_1_185_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .src128(src128),
        .src129(src129),
        .src130(src130),
        .src131(src131),
        .src132(src132),
        .src133(src133),
        .src134(src134),
        .src135(src135),
        .src136(src136),
        .src137(src137),
        .src138(src138),
        .src139(src139),
        .src140(src140),
        .src141(src141),
        .src142(src142),
        .src143(src143),
        .src144(src144),
        .src145(src145),
        .src146(src146),
        .src147(src147),
        .src148(src148),
        .src149(src149),
        .src150(src150),
        .src151(src151),
        .src152(src152),
        .src153(src153),
        .src154(src154),
        .src155(src155),
        .src156(src156),
        .src157(src157),
        .src158(src158),
        .src159(src159),
        .src160(src160),
        .src161(src161),
        .src162(src162),
        .src163(src163),
        .src164(src164),
        .src165(src165),
        .src166(src166),
        .src167(src167),
        .src168(src168),
        .src169(src169),
        .src170(src170),
        .src171(src171),
        .src172(src172),
        .src173(src173),
        .src174(src174),
        .src175(src175),
        .src176(src176),
        .src177(src177),
        .src178(src178),
        .src179(src179),
        .src180(src180),
        .src181(src181),
        .src182(src182),
        .src183(src183),
        .src184(src184),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, src128, src129, src130, src131, src132, src133, src134, src135, src136, src137, src138, src139, src140, src141, src142, src143, src144, src145, src146, src147, src148, src149, src150, src151, src152, src153, src154, src155, src156, src157, src158, src159, src160, src161, src162, src163, src164, src165, src166, src167, src168, src169, src170, src171, src172, src173, src174, src175, src176, src177, src178, src179, src180, src181, src182, src183, src184, dst, exp, test);
        src0 <= 16'ha071;
        src1 <= 16'h9d8c;
        src2 <= 16'h4f75;
        src3 <= 16'h1250;
        src4 <= 16'he7fb;
        src5 <= 16'h1ca0;
        src6 <= 16'hb74f;
        src7 <= 16'hbfd;
        src8 <= 16'h8c0a;
        src9 <= 16'he497;
        src10 <= 16'hcb34;
        src11 <= 16'hbc48;
        src12 <= 16'h4997;
        src13 <= 16'h31f;
        src14 <= 16'hdbbc;
        src15 <= 16'hd7db;
        src16 <= 16'h47d1;
        src17 <= 16'h151f;
        src18 <= 16'h1846;
        src19 <= 16'h21c4;
        src20 <= 16'h9b8b;
        src21 <= 16'hf3cf;
        src22 <= 16'hf925;
        src23 <= 16'h3d8f;
        src24 <= 16'h6f1b;
        src25 <= 16'h860d;
        src26 <= 16'hab03;
        src27 <= 16'hd71f;
        src28 <= 16'h9bfb;
        src29 <= 16'hba26;
        src30 <= 16'hc535;
        src31 <= 16'hf7a3;
        src32 <= 16'h56a8;
        src33 <= 16'hca82;
        src34 <= 16'h13b1;
        src35 <= 16'he28a;
        src36 <= 16'h3cd2;
        src37 <= 16'hdb24;
        src38 <= 16'h2b10;
        src39 <= 16'hf8bd;
        src40 <= 16'h77ac;
        src41 <= 16'h4d78;
        src42 <= 16'hbbda;
        src43 <= 16'h6fe0;
        src44 <= 16'hea7f;
        src45 <= 16'ha554;
        src46 <= 16'hc104;
        src47 <= 16'hba40;
        src48 <= 16'h7e7d;
        src49 <= 16'hf8f8;
        src50 <= 16'hf3f1;
        src51 <= 16'hd81b;
        src52 <= 16'ha689;
        src53 <= 16'h24ea;
        src54 <= 16'hc9b9;
        src55 <= 16'h1ad4;
        src56 <= 16'h7b09;
        src57 <= 16'hc29b;
        src58 <= 16'hdae4;
        src59 <= 16'hc1a6;
        src60 <= 16'hac9;
        src61 <= 16'hde6;
        src62 <= 16'h89c6;
        src63 <= 16'h8094;
        src64 <= 16'hac6;
        src65 <= 16'hd003;
        src66 <= 16'hb837;
        src67 <= 16'h5ce3;
        src68 <= 16'hdf1e;
        src69 <= 16'hb6b2;
        src70 <= 16'h77a8;
        src71 <= 16'h438b;
        src72 <= 16'hfadf;
        src73 <= 16'h6dd5;
        src74 <= 16'h38c8;
        src75 <= 16'h6a87;
        src76 <= 16'hdbb5;
        src77 <= 16'h9855;
        src78 <= 16'hdc11;
        src79 <= 16'hdd8d;
        src80 <= 16'h2230;
        src81 <= 16'hdd16;
        src82 <= 16'h7e50;
        src83 <= 16'hd3e2;
        src84 <= 16'h85be;
        src85 <= 16'h423d;
        src86 <= 16'hc564;
        src87 <= 16'h3103;
        src88 <= 16'h14fa;
        src89 <= 16'h3766;
        src90 <= 16'hfd9;
        src91 <= 16'h512e;
        src92 <= 16'h340a;
        src93 <= 16'h42d9;
        src94 <= 16'h554f;
        src95 <= 16'hd01e;
        src96 <= 16'hbbe2;
        src97 <= 16'he1e5;
        src98 <= 16'hac0b;
        src99 <= 16'h8dae;
        src100 <= 16'ha93c;
        src101 <= 16'h236f;
        src102 <= 16'hb9cf;
        src103 <= 16'h5719;
        src104 <= 16'h424e;
        src105 <= 16'h6fc1;
        src106 <= 16'h7ac3;
        src107 <= 16'h7e64;
        src108 <= 16'h5042;
        src109 <= 16'h1fa4;
        src110 <= 16'h8ccf;
        src111 <= 16'h638d;
        src112 <= 16'hca16;
        src113 <= 16'h4595;
        src114 <= 16'h9482;
        src115 <= 16'he77d;
        src116 <= 16'h8a57;
        src117 <= 16'h29a0;
        src118 <= 16'h2e01;
        src119 <= 16'he309;
        src120 <= 16'h3c4;
        src121 <= 16'h908d;
        src122 <= 16'hf57a;
        src123 <= 16'hc28e;
        src124 <= 16'hf9b6;
        src125 <= 16'h1cf9;
        src126 <= 16'h22f4;
        src127 <= 16'h624;
        src128 <= 16'haa3f;
        src129 <= 16'h5ca8;
        src130 <= 16'h1756;
        src131 <= 16'h3a38;
        src132 <= 16'h4c01;
        src133 <= 16'h25aa;
        src134 <= 16'h7404;
        src135 <= 16'h4f1;
        src136 <= 16'hf354;
        src137 <= 16'hae7;
        src138 <= 16'h3f6b;
        src139 <= 16'h97f9;
        src140 <= 16'h7342;
        src141 <= 16'hc44a;
        src142 <= 16'he14d;
        src143 <= 16'h441;
        src144 <= 16'h6b03;
        src145 <= 16'hb2b4;
        src146 <= 16'h55d;
        src147 <= 16'h7a5d;
        src148 <= 16'h5c02;
        src149 <= 16'h5462;
        src150 <= 16'hd2ff;
        src151 <= 16'h86d1;
        src152 <= 16'hae0;
        src153 <= 16'h83d3;
        src154 <= 16'h5551;
        src155 <= 16'h8bf2;
        src156 <= 16'h879c;
        src157 <= 16'h8815;
        src158 <= 16'h9a64;
        src159 <= 16'h3c12;
        src160 <= 16'h9686;
        src161 <= 16'hd478;
        src162 <= 16'h70fb;
        src163 <= 16'h982c;
        src164 <= 16'hb1c7;
        src165 <= 16'hb646;
        src166 <= 16'hc483;
        src167 <= 16'hdffc;
        src168 <= 16'h8a96;
        src169 <= 16'hecf3;
        src170 <= 16'h486;
        src171 <= 16'h6d6b;
        src172 <= 16'h181f;
        src173 <= 16'h4eb4;
        src174 <= 16'h77b4;
        src175 <= 16'h131e;
        src176 <= 16'ha608;
        src177 <= 16'hfdc8;
        src178 <= 16'hc33a;
        src179 <= 16'hba3c;
        src180 <= 16'h5aba;
        src181 <= 16'h6afa;
        src182 <= 16'h643d;
        src183 <= 16'hafd7;
        src184 <= 16'h92ff;
        exp <= 24'h5e1618;
        #1
        src0 <= 16'h3aba;
        src1 <= 16'h142b;
        src2 <= 16'h87c9;
        src3 <= 16'hfd25;
        src4 <= 16'h6c57;
        src5 <= 16'h12b9;
        src6 <= 16'hf9c5;
        src7 <= 16'h8d0;
        src8 <= 16'hb641;
        src9 <= 16'h2d97;
        src10 <= 16'h6858;
        src11 <= 16'h5f0a;
        src12 <= 16'h7b1d;
        src13 <= 16'hc55b;
        src14 <= 16'h4a3d;
        src15 <= 16'hdf4e;
        src16 <= 16'h7971;
        src17 <= 16'h8a5f;
        src18 <= 16'h7953;
        src19 <= 16'h1b27;
        src20 <= 16'h4a9a;
        src21 <= 16'h7216;
        src22 <= 16'h5512;
        src23 <= 16'h25e7;
        src24 <= 16'hc5e2;
        src25 <= 16'h503e;
        src26 <= 16'hc60a;
        src27 <= 16'h2adc;
        src28 <= 16'hf8a0;
        src29 <= 16'hd62e;
        src30 <= 16'h8434;
        src31 <= 16'he5b1;
        src32 <= 16'hda18;
        src33 <= 16'h2236;
        src34 <= 16'hff00;
        src35 <= 16'h597b;
        src36 <= 16'hd5fc;
        src37 <= 16'h34b;
        src38 <= 16'h4a9c;
        src39 <= 16'hfda5;
        src40 <= 16'hce59;
        src41 <= 16'h97e;
        src42 <= 16'h8cd2;
        src43 <= 16'h64d7;
        src44 <= 16'h28a2;
        src45 <= 16'h6175;
        src46 <= 16'h73d3;
        src47 <= 16'hbff6;
        src48 <= 16'he7b1;
        src49 <= 16'hd868;
        src50 <= 16'h47a3;
        src51 <= 16'h98d3;
        src52 <= 16'h338a;
        src53 <= 16'had9e;
        src54 <= 16'h243c;
        src55 <= 16'hd38d;
        src56 <= 16'h6f77;
        src57 <= 16'h1834;
        src58 <= 16'h3649;
        src59 <= 16'hc799;
        src60 <= 16'hdbc1;
        src61 <= 16'h54db;
        src62 <= 16'h4c7d;
        src63 <= 16'h85cd;
        src64 <= 16'h966c;
        src65 <= 16'hed11;
        src66 <= 16'ha41d;
        src67 <= 16'hc200;
        src68 <= 16'h67e3;
        src69 <= 16'hc06a;
        src70 <= 16'h459e;
        src71 <= 16'hca4b;
        src72 <= 16'hd83b;
        src73 <= 16'h1ac4;
        src74 <= 16'h8a20;
        src75 <= 16'h9ad8;
        src76 <= 16'hdab6;
        src77 <= 16'hd377;
        src78 <= 16'hecbb;
        src79 <= 16'h6449;
        src80 <= 16'h15c4;
        src81 <= 16'h77b4;
        src82 <= 16'hd74b;
        src83 <= 16'h1254;
        src84 <= 16'h19be;
        src85 <= 16'hee30;
        src86 <= 16'hccac;
        src87 <= 16'h47f8;
        src88 <= 16'h87d8;
        src89 <= 16'ha99a;
        src90 <= 16'h52b1;
        src91 <= 16'h3502;
        src92 <= 16'h251;
        src93 <= 16'hf191;
        src94 <= 16'hb00;
        src95 <= 16'he759;
        src96 <= 16'hc789;
        src97 <= 16'hfb80;
        src98 <= 16'ha3ed;
        src99 <= 16'h6c64;
        src100 <= 16'h2221;
        src101 <= 16'hc93c;
        src102 <= 16'hbad8;
        src103 <= 16'h14a7;
        src104 <= 16'h4cbd;
        src105 <= 16'h2e3f;
        src106 <= 16'h9ff5;
        src107 <= 16'h4daa;
        src108 <= 16'hfec;
        src109 <= 16'h4567;
        src110 <= 16'hbda3;
        src111 <= 16'hcda5;
        src112 <= 16'hee39;
        src113 <= 16'hff5d;
        src114 <= 16'h4c77;
        src115 <= 16'h985b;
        src116 <= 16'ha9ae;
        src117 <= 16'h5f52;
        src118 <= 16'h6147;
        src119 <= 16'h52c4;
        src120 <= 16'h44f4;
        src121 <= 16'hb373;
        src122 <= 16'hefab;
        src123 <= 16'h8174;
        src124 <= 16'h31f5;
        src125 <= 16'h95cd;
        src126 <= 16'h31f7;
        src127 <= 16'h497;
        src128 <= 16'hbdc6;
        src129 <= 16'he178;
        src130 <= 16'h7c16;
        src131 <= 16'h1722;
        src132 <= 16'hab14;
        src133 <= 16'h9ddf;
        src134 <= 16'hfff7;
        src135 <= 16'h2661;
        src136 <= 16'he7da;
        src137 <= 16'h3203;
        src138 <= 16'h21be;
        src139 <= 16'h4600;
        src140 <= 16'h625e;
        src141 <= 16'h13e7;
        src142 <= 16'h6519;
        src143 <= 16'h6ce2;
        src144 <= 16'had03;
        src145 <= 16'h9fbb;
        src146 <= 16'h4223;
        src147 <= 16'h322b;
        src148 <= 16'h666c;
        src149 <= 16'h5d3c;
        src150 <= 16'h58d4;
        src151 <= 16'hb0df;
        src152 <= 16'h5ca2;
        src153 <= 16'hb142;
        src154 <= 16'heda8;
        src155 <= 16'h7e7d;
        src156 <= 16'h148d;
        src157 <= 16'hed47;
        src158 <= 16'h2a4d;
        src159 <= 16'h1372;
        src160 <= 16'h2eb6;
        src161 <= 16'he70b;
        src162 <= 16'h65fb;
        src163 <= 16'hd9b6;
        src164 <= 16'h2b81;
        src165 <= 16'h40d0;
        src166 <= 16'h9763;
        src167 <= 16'h6bf6;
        src168 <= 16'h24f5;
        src169 <= 16'he8d2;
        src170 <= 16'h36de;
        src171 <= 16'h6de7;
        src172 <= 16'h470e;
        src173 <= 16'he527;
        src174 <= 16'hd29e;
        src175 <= 16'h85d3;
        src176 <= 16'ha2fe;
        src177 <= 16'hdb1b;
        src178 <= 16'h7e2f;
        src179 <= 16'h6650;
        src180 <= 16'hcf28;
        src181 <= 16'h6b39;
        src182 <= 16'h47e9;
        src183 <= 16'hf02f;
        src184 <= 16'h90f0;
        exp <= 24'h5ccaa9;
        #1
        src0 <= 16'h2a74;
        src1 <= 16'he24e;
        src2 <= 16'h6cee;
        src3 <= 16'hedd2;
        src4 <= 16'h4457;
        src5 <= 16'h2bb4;
        src6 <= 16'h8ecd;
        src7 <= 16'h34f4;
        src8 <= 16'h867b;
        src9 <= 16'he176;
        src10 <= 16'h4891;
        src11 <= 16'hdd6d;
        src12 <= 16'h96b9;
        src13 <= 16'h4578;
        src14 <= 16'he7d4;
        src15 <= 16'hb857;
        src16 <= 16'h433f;
        src17 <= 16'hf635;
        src18 <= 16'h8e1e;
        src19 <= 16'h2cbe;
        src20 <= 16'hc106;
        src21 <= 16'h4c83;
        src22 <= 16'h6c37;
        src23 <= 16'ha528;
        src24 <= 16'h4485;
        src25 <= 16'hf2da;
        src26 <= 16'h5cf1;
        src27 <= 16'hf6b6;
        src28 <= 16'h8581;
        src29 <= 16'h77c4;
        src30 <= 16'hd8c9;
        src31 <= 16'h3ee2;
        src32 <= 16'h3503;
        src33 <= 16'h71c0;
        src34 <= 16'h9fd0;
        src35 <= 16'h6641;
        src36 <= 16'hf145;
        src37 <= 16'h4760;
        src38 <= 16'h93b4;
        src39 <= 16'h805;
        src40 <= 16'h66b6;
        src41 <= 16'h6600;
        src42 <= 16'h68f8;
        src43 <= 16'h413f;
        src44 <= 16'h98d1;
        src45 <= 16'h3fbd;
        src46 <= 16'hd7c6;
        src47 <= 16'hdbc1;
        src48 <= 16'h8cc7;
        src49 <= 16'h91c5;
        src50 <= 16'h8a24;
        src51 <= 16'h19c0;
        src52 <= 16'hb88e;
        src53 <= 16'haa0e;
        src54 <= 16'hed78;
        src55 <= 16'h334a;
        src56 <= 16'h85b5;
        src57 <= 16'h2c47;
        src58 <= 16'he0d6;
        src59 <= 16'h1f63;
        src60 <= 16'h6e00;
        src61 <= 16'h9c20;
        src62 <= 16'hd908;
        src63 <= 16'h1ed8;
        src64 <= 16'h4d64;
        src65 <= 16'hf753;
        src66 <= 16'he374;
        src67 <= 16'h73e1;
        src68 <= 16'hdad0;
        src69 <= 16'h3f47;
        src70 <= 16'hc576;
        src71 <= 16'hefa2;
        src72 <= 16'hb191;
        src73 <= 16'hea4f;
        src74 <= 16'h909;
        src75 <= 16'h7c26;
        src76 <= 16'h75e3;
        src77 <= 16'h5bd;
        src78 <= 16'hafd8;
        src79 <= 16'hbd02;
        src80 <= 16'hf224;
        src81 <= 16'hff9f;
        src82 <= 16'ha04b;
        src83 <= 16'hee3d;
        src84 <= 16'h5bfe;
        src85 <= 16'hc64c;
        src86 <= 16'hb0fa;
        src87 <= 16'hd9b5;
        src88 <= 16'he199;
        src89 <= 16'h8008;
        src90 <= 16'h4ade;
        src91 <= 16'h31c3;
        src92 <= 16'h1b40;
        src93 <= 16'h83ab;
        src94 <= 16'hb25e;
        src95 <= 16'hd1df;
        src96 <= 16'h9519;
        src97 <= 16'hfe5f;
        src98 <= 16'ha5cc;
        src99 <= 16'h7e16;
        src100 <= 16'h3e7a;
        src101 <= 16'h3247;
        src102 <= 16'h39fb;
        src103 <= 16'hab77;
        src104 <= 16'h6b3a;
        src105 <= 16'h546;
        src106 <= 16'hb2f;
        src107 <= 16'h77ac;
        src108 <= 16'h518c;
        src109 <= 16'h75a5;
        src110 <= 16'h4eaf;
        src111 <= 16'h337;
        src112 <= 16'h37ed;
        src113 <= 16'hdf64;
        src114 <= 16'hd07a;
        src115 <= 16'hff10;
        src116 <= 16'h3ddb;
        src117 <= 16'hff0e;
        src118 <= 16'h1afc;
        src119 <= 16'h6794;
        src120 <= 16'h58f7;
        src121 <= 16'h66e0;
        src122 <= 16'hf01b;
        src123 <= 16'h7d2;
        src124 <= 16'h55ae;
        src125 <= 16'h2ed3;
        src126 <= 16'h2882;
        src127 <= 16'h12df;
        src128 <= 16'hd583;
        src129 <= 16'h7dab;
        src130 <= 16'hc95f;
        src131 <= 16'h13fd;
        src132 <= 16'h9763;
        src133 <= 16'hb570;
        src134 <= 16'h4b6b;
        src135 <= 16'h9b10;
        src136 <= 16'hd27;
        src137 <= 16'h396c;
        src138 <= 16'h46dc;
        src139 <= 16'h82fe;
        src140 <= 16'ha050;
        src141 <= 16'h8b2d;
        src142 <= 16'h9876;
        src143 <= 16'h35f9;
        src144 <= 16'hb959;
        src145 <= 16'hbb8a;
        src146 <= 16'hedb3;
        src147 <= 16'h9ef5;
        src148 <= 16'h2724;
        src149 <= 16'h2620;
        src150 <= 16'hde0a;
        src151 <= 16'h6ff1;
        src152 <= 16'h6cfc;
        src153 <= 16'hd766;
        src154 <= 16'h54fa;
        src155 <= 16'hfa79;
        src156 <= 16'ha207;
        src157 <= 16'he476;
        src158 <= 16'h9ee;
        src159 <= 16'h9297;
        src160 <= 16'h2f4d;
        src161 <= 16'hf00b;
        src162 <= 16'h9f56;
        src163 <= 16'h338a;
        src164 <= 16'he238;
        src165 <= 16'h4a99;
        src166 <= 16'h7b77;
        src167 <= 16'h724a;
        src168 <= 16'h9d84;
        src169 <= 16'h1ef7;
        src170 <= 16'h8eae;
        src171 <= 16'ha4be;
        src172 <= 16'h24a2;
        src173 <= 16'h95e5;
        src174 <= 16'hab64;
        src175 <= 16'h3464;
        src176 <= 16'ha843;
        src177 <= 16'h90d4;
        src178 <= 16'h9e60;
        src179 <= 16'hdbc0;
        src180 <= 16'hce01;
        src181 <= 16'h3eeb;
        src182 <= 16'h1c20;
        src183 <= 16'heb23;
        src184 <= 16'hdf58;
        exp <= 24'h5fb1f9;
        #1
        src0 <= 16'h2282;
        src1 <= 16'h35e0;
        src2 <= 16'h7755;
        src3 <= 16'h79a3;
        src4 <= 16'h3606;
        src5 <= 16'h930a;
        src6 <= 16'h3b0f;
        src7 <= 16'hc931;
        src8 <= 16'h5b18;
        src9 <= 16'he11c;
        src10 <= 16'h35bb;
        src11 <= 16'hfb0d;
        src12 <= 16'ha54a;
        src13 <= 16'h30af;
        src14 <= 16'h2b84;
        src15 <= 16'h80d1;
        src16 <= 16'hefd5;
        src17 <= 16'hd4b1;
        src18 <= 16'h7207;
        src19 <= 16'h9a9b;
        src20 <= 16'h5b0c;
        src21 <= 16'ha1ce;
        src22 <= 16'h5cd2;
        src23 <= 16'h9fae;
        src24 <= 16'h5c02;
        src25 <= 16'he146;
        src26 <= 16'hf973;
        src27 <= 16'hb9ab;
        src28 <= 16'h1d8d;
        src29 <= 16'h1b03;
        src30 <= 16'hfb62;
        src31 <= 16'hd8b3;
        src32 <= 16'h3d94;
        src33 <= 16'h2bd2;
        src34 <= 16'h66e0;
        src35 <= 16'hde42;
        src36 <= 16'he29a;
        src37 <= 16'h5370;
        src38 <= 16'hbfa2;
        src39 <= 16'h4781;
        src40 <= 16'h87f7;
        src41 <= 16'hc36b;
        src42 <= 16'h5f6f;
        src43 <= 16'he91e;
        src44 <= 16'h8fd1;
        src45 <= 16'h23d9;
        src46 <= 16'h5341;
        src47 <= 16'hadbb;
        src48 <= 16'h4d95;
        src49 <= 16'h556c;
        src50 <= 16'hc18c;
        src51 <= 16'ha9ae;
        src52 <= 16'h97e7;
        src53 <= 16'h95a9;
        src54 <= 16'h55b8;
        src55 <= 16'h30c0;
        src56 <= 16'he13a;
        src57 <= 16'h88aa;
        src58 <= 16'hc4e3;
        src59 <= 16'h4bff;
        src60 <= 16'h3bdc;
        src61 <= 16'h8534;
        src62 <= 16'h1195;
        src63 <= 16'h78f;
        src64 <= 16'h1316;
        src65 <= 16'h7823;
        src66 <= 16'hccf6;
        src67 <= 16'ha7e;
        src68 <= 16'h67e2;
        src69 <= 16'hf84f;
        src70 <= 16'h1137;
        src71 <= 16'hcb0f;
        src72 <= 16'hd416;
        src73 <= 16'h156f;
        src74 <= 16'hb4bb;
        src75 <= 16'hf0d6;
        src76 <= 16'ha460;
        src77 <= 16'h1b8;
        src78 <= 16'hd089;
        src79 <= 16'h5105;
        src80 <= 16'h6afb;
        src81 <= 16'ha52a;
        src82 <= 16'h5051;
        src83 <= 16'h6346;
        src84 <= 16'hf763;
        src85 <= 16'h4d1f;
        src86 <= 16'h474b;
        src87 <= 16'h1c97;
        src88 <= 16'h4c36;
        src89 <= 16'h4d58;
        src90 <= 16'hd5d0;
        src91 <= 16'hfd3e;
        src92 <= 16'hef16;
        src93 <= 16'h5a92;
        src94 <= 16'hc916;
        src95 <= 16'h1218;
        src96 <= 16'hde06;
        src97 <= 16'h1e03;
        src98 <= 16'hc0f9;
        src99 <= 16'hb549;
        src100 <= 16'hf7da;
        src101 <= 16'h226a;
        src102 <= 16'h79c7;
        src103 <= 16'h3cf3;
        src104 <= 16'h8364;
        src105 <= 16'hafd4;
        src106 <= 16'h949c;
        src107 <= 16'he98b;
        src108 <= 16'hb87c;
        src109 <= 16'h18ed;
        src110 <= 16'h769c;
        src111 <= 16'h8e1d;
        src112 <= 16'h75ac;
        src113 <= 16'h51cb;
        src114 <= 16'he9d8;
        src115 <= 16'h35a;
        src116 <= 16'h5897;
        src117 <= 16'hb71;
        src118 <= 16'h7e20;
        src119 <= 16'h1557;
        src120 <= 16'h9885;
        src121 <= 16'hc2c2;
        src122 <= 16'hd291;
        src123 <= 16'h93a;
        src124 <= 16'h744b;
        src125 <= 16'ha8a8;
        src126 <= 16'hd953;
        src127 <= 16'h900f;
        src128 <= 16'h2a92;
        src129 <= 16'h1eae;
        src130 <= 16'hc861;
        src131 <= 16'h7ce;
        src132 <= 16'h5d2c;
        src133 <= 16'h1c18;
        src134 <= 16'ha37f;
        src135 <= 16'h864a;
        src136 <= 16'h7cd3;
        src137 <= 16'h7716;
        src138 <= 16'h8496;
        src139 <= 16'h880b;
        src140 <= 16'hd9a0;
        src141 <= 16'he602;
        src142 <= 16'hbda4;
        src143 <= 16'h24d0;
        src144 <= 16'h4630;
        src145 <= 16'h939d;
        src146 <= 16'hfdb4;
        src147 <= 16'h5906;
        src148 <= 16'h6cb0;
        src149 <= 16'h2016;
        src150 <= 16'h5ec1;
        src151 <= 16'h2975;
        src152 <= 16'hca6c;
        src153 <= 16'hb901;
        src154 <= 16'h2d52;
        src155 <= 16'h791;
        src156 <= 16'hc383;
        src157 <= 16'ha462;
        src158 <= 16'hcb76;
        src159 <= 16'hae13;
        src160 <= 16'h768c;
        src161 <= 16'hc24d;
        src162 <= 16'hbda4;
        src163 <= 16'ha4bc;
        src164 <= 16'hd314;
        src165 <= 16'h172f;
        src166 <= 16'h80d8;
        src167 <= 16'had03;
        src168 <= 16'hc2a6;
        src169 <= 16'hb24b;
        src170 <= 16'h6978;
        src171 <= 16'h5bad;
        src172 <= 16'h1e36;
        src173 <= 16'h348a;
        src174 <= 16'ha2d9;
        src175 <= 16'h3150;
        src176 <= 16'h802f;
        src177 <= 16'he4f1;
        src178 <= 16'h3b23;
        src179 <= 16'h5e9b;
        src180 <= 16'hf937;
        src181 <= 16'h34c1;
        src182 <= 16'hf897;
        src183 <= 16'h507e;
        src184 <= 16'h3f31;
        exp <= 24'h5c48a2;
        #1
        src0 <= 16'h9950;
        src1 <= 16'hae96;
        src2 <= 16'h75e9;
        src3 <= 16'h2113;
        src4 <= 16'h35e5;
        src5 <= 16'h48d;
        src6 <= 16'h181a;
        src7 <= 16'h5c30;
        src8 <= 16'hccc5;
        src9 <= 16'h6e3d;
        src10 <= 16'h9f23;
        src11 <= 16'hb716;
        src12 <= 16'he7e;
        src13 <= 16'h217b;
        src14 <= 16'hbd8b;
        src15 <= 16'hc288;
        src16 <= 16'h8b7e;
        src17 <= 16'h3247;
        src18 <= 16'h67b8;
        src19 <= 16'hdea;
        src20 <= 16'h6d4c;
        src21 <= 16'h8826;
        src22 <= 16'h1b0c;
        src23 <= 16'h1ba4;
        src24 <= 16'h34ec;
        src25 <= 16'h9124;
        src26 <= 16'h1e21;
        src27 <= 16'ha3d4;
        src28 <= 16'hebe6;
        src29 <= 16'h2168;
        src30 <= 16'ha326;
        src31 <= 16'h419f;
        src32 <= 16'hef53;
        src33 <= 16'h61eb;
        src34 <= 16'h60cf;
        src35 <= 16'hbd59;
        src36 <= 16'h1480;
        src37 <= 16'haada;
        src38 <= 16'h805d;
        src39 <= 16'h3eec;
        src40 <= 16'h64ed;
        src41 <= 16'hcac5;
        src42 <= 16'h3e5e;
        src43 <= 16'hc505;
        src44 <= 16'h7cbf;
        src45 <= 16'hd879;
        src46 <= 16'h54e2;
        src47 <= 16'hbb71;
        src48 <= 16'h84f8;
        src49 <= 16'h1053;
        src50 <= 16'hd5a3;
        src51 <= 16'h6224;
        src52 <= 16'h8e23;
        src53 <= 16'h720f;
        src54 <= 16'ha21e;
        src55 <= 16'hce64;
        src56 <= 16'h4661;
        src57 <= 16'h9ea8;
        src58 <= 16'hd9f0;
        src59 <= 16'h3aac;
        src60 <= 16'h3d2d;
        src61 <= 16'h7c52;
        src62 <= 16'hf13;
        src63 <= 16'h84bc;
        src64 <= 16'hd00e;
        src65 <= 16'hd825;
        src66 <= 16'hade4;
        src67 <= 16'hae4d;
        src68 <= 16'h6613;
        src69 <= 16'h5992;
        src70 <= 16'hd8eb;
        src71 <= 16'hf354;
        src72 <= 16'h48ce;
        src73 <= 16'h6071;
        src74 <= 16'h40f4;
        src75 <= 16'h48bd;
        src76 <= 16'h9ec3;
        src77 <= 16'hb652;
        src78 <= 16'ha7b3;
        src79 <= 16'h3f5b;
        src80 <= 16'ha56f;
        src81 <= 16'h7524;
        src82 <= 16'h5b00;
        src83 <= 16'h48cc;
        src84 <= 16'h8702;
        src85 <= 16'h2a30;
        src86 <= 16'heaeb;
        src87 <= 16'h4bf;
        src88 <= 16'he8b0;
        src89 <= 16'h5428;
        src90 <= 16'h8de0;
        src91 <= 16'h119d;
        src92 <= 16'hb710;
        src93 <= 16'h8b82;
        src94 <= 16'h69d2;
        src95 <= 16'h6070;
        src96 <= 16'h2d10;
        src97 <= 16'h5e3d;
        src98 <= 16'h89a8;
        src99 <= 16'h4af9;
        src100 <= 16'hc902;
        src101 <= 16'h73b7;
        src102 <= 16'hb30e;
        src103 <= 16'h2d00;
        src104 <= 16'ha493;
        src105 <= 16'h9815;
        src106 <= 16'h8d0f;
        src107 <= 16'h5f04;
        src108 <= 16'h5e9b;
        src109 <= 16'h5161;
        src110 <= 16'hf3af;
        src111 <= 16'h424c;
        src112 <= 16'hc09;
        src113 <= 16'ha93d;
        src114 <= 16'h5400;
        src115 <= 16'h465d;
        src116 <= 16'hb8e7;
        src117 <= 16'hbe84;
        src118 <= 16'h5d40;
        src119 <= 16'h6ed;
        src120 <= 16'h5e7a;
        src121 <= 16'hea45;
        src122 <= 16'h4583;
        src123 <= 16'h53d7;
        src124 <= 16'h5904;
        src125 <= 16'h99bb;
        src126 <= 16'hafe0;
        src127 <= 16'h881a;
        src128 <= 16'h3176;
        src129 <= 16'h3ec9;
        src130 <= 16'h8105;
        src131 <= 16'hd7c5;
        src132 <= 16'hbcd5;
        src133 <= 16'he0c1;
        src134 <= 16'h6398;
        src135 <= 16'hd1b0;
        src136 <= 16'he0cb;
        src137 <= 16'h6415;
        src138 <= 16'hcc5f;
        src139 <= 16'hab50;
        src140 <= 16'h3a60;
        src141 <= 16'hed49;
        src142 <= 16'h859;
        src143 <= 16'hf1e3;
        src144 <= 16'h163a;
        src145 <= 16'hd7d5;
        src146 <= 16'ha84d;
        src147 <= 16'he49;
        src148 <= 16'h4cec;
        src149 <= 16'h7be9;
        src150 <= 16'h7479;
        src151 <= 16'h9cfd;
        src152 <= 16'hb13e;
        src153 <= 16'h3df8;
        src154 <= 16'h7909;
        src155 <= 16'h8492;
        src156 <= 16'hce52;
        src157 <= 16'h1230;
        src158 <= 16'hba86;
        src159 <= 16'he47;
        src160 <= 16'hce1e;
        src161 <= 16'hc804;
        src162 <= 16'h5540;
        src163 <= 16'h7216;
        src164 <= 16'ha56d;
        src165 <= 16'h9351;
        src166 <= 16'h41ab;
        src167 <= 16'h2f24;
        src168 <= 16'h6c79;
        src169 <= 16'hb568;
        src170 <= 16'hc667;
        src171 <= 16'h76ed;
        src172 <= 16'hc1ed;
        src173 <= 16'hb194;
        src174 <= 16'h15cd;
        src175 <= 16'ha2c2;
        src176 <= 16'h6de7;
        src177 <= 16'hb4ad;
        src178 <= 16'hbb1c;
        src179 <= 16'h581e;
        src180 <= 16'h5e1d;
        src181 <= 16'hf7b6;
        src182 <= 16'he62b;
        src183 <= 16'hc40b;
        src184 <= 16'had19;
        exp <= 24'h5ac3c0;
        #1
        src0 <= 16'h321a;
        src1 <= 16'h70fd;
        src2 <= 16'h996d;
        src3 <= 16'ha3a5;
        src4 <= 16'hc38e;
        src5 <= 16'hc126;
        src6 <= 16'h198b;
        src7 <= 16'ha45d;
        src8 <= 16'h2a67;
        src9 <= 16'h9d78;
        src10 <= 16'h7677;
        src11 <= 16'h4a1b;
        src12 <= 16'he98;
        src13 <= 16'h41c2;
        src14 <= 16'h4a4f;
        src15 <= 16'hfe28;
        src16 <= 16'hf881;
        src17 <= 16'h8816;
        src18 <= 16'h181d;
        src19 <= 16'h2b76;
        src20 <= 16'hdb5b;
        src21 <= 16'h73c5;
        src22 <= 16'h48c9;
        src23 <= 16'ha740;
        src24 <= 16'h3278;
        src25 <= 16'h2663;
        src26 <= 16'h41db;
        src27 <= 16'hd763;
        src28 <= 16'hb281;
        src29 <= 16'heb86;
        src30 <= 16'h8057;
        src31 <= 16'h57a5;
        src32 <= 16'hadd6;
        src33 <= 16'h1cc4;
        src34 <= 16'hfcca;
        src35 <= 16'he41e;
        src36 <= 16'h7c6c;
        src37 <= 16'hfc9a;
        src38 <= 16'hbd56;
        src39 <= 16'hb676;
        src40 <= 16'h9970;
        src41 <= 16'ha64c;
        src42 <= 16'h734a;
        src43 <= 16'h905c;
        src44 <= 16'hc83b;
        src45 <= 16'h1ad6;
        src46 <= 16'h3663;
        src47 <= 16'h7b0b;
        src48 <= 16'h2c22;
        src49 <= 16'h6973;
        src50 <= 16'hc6d;
        src51 <= 16'h31cb;
        src52 <= 16'h3499;
        src53 <= 16'heff2;
        src54 <= 16'h8031;
        src55 <= 16'he391;
        src56 <= 16'h5fa4;
        src57 <= 16'hc314;
        src58 <= 16'h4764;
        src59 <= 16'h39b3;
        src60 <= 16'h3c6c;
        src61 <= 16'h277f;
        src62 <= 16'h8a72;
        src63 <= 16'hb97e;
        src64 <= 16'h2fce;
        src65 <= 16'h270c;
        src66 <= 16'had2c;
        src67 <= 16'h7675;
        src68 <= 16'hf05e;
        src69 <= 16'ha5d6;
        src70 <= 16'h1aa9;
        src71 <= 16'h6324;
        src72 <= 16'h5843;
        src73 <= 16'h8748;
        src74 <= 16'hac97;
        src75 <= 16'hd482;
        src76 <= 16'h55de;
        src77 <= 16'h7682;
        src78 <= 16'h505b;
        src79 <= 16'h75d6;
        src80 <= 16'ha635;
        src81 <= 16'h57ac;
        src82 <= 16'h7c8c;
        src83 <= 16'h7435;
        src84 <= 16'h9b49;
        src85 <= 16'ha955;
        src86 <= 16'hf9dd;
        src87 <= 16'h44fc;
        src88 <= 16'h75bd;
        src89 <= 16'h93e9;
        src90 <= 16'h7082;
        src91 <= 16'h70ba;
        src92 <= 16'h5acf;
        src93 <= 16'h846;
        src94 <= 16'h452;
        src95 <= 16'h78af;
        src96 <= 16'h639e;
        src97 <= 16'hed5;
        src98 <= 16'h1ffa;
        src99 <= 16'h9f65;
        src100 <= 16'hd77c;
        src101 <= 16'hc952;
        src102 <= 16'hc5df;
        src103 <= 16'hd6eb;
        src104 <= 16'hae35;
        src105 <= 16'he7f6;
        src106 <= 16'h5ffd;
        src107 <= 16'haabc;
        src108 <= 16'hbfc;
        src109 <= 16'h725c;
        src110 <= 16'hc779;
        src111 <= 16'hee68;
        src112 <= 16'hd46a;
        src113 <= 16'he3ab;
        src114 <= 16'h1779;
        src115 <= 16'hb069;
        src116 <= 16'he75b;
        src117 <= 16'h30fe;
        src118 <= 16'h500e;
        src119 <= 16'h3482;
        src120 <= 16'h4130;
        src121 <= 16'h576e;
        src122 <= 16'hf705;
        src123 <= 16'h2a2a;
        src124 <= 16'h2532;
        src125 <= 16'hbd4;
        src126 <= 16'hd30b;
        src127 <= 16'h976f;
        src128 <= 16'h6a0;
        src129 <= 16'hd76a;
        src130 <= 16'he524;
        src131 <= 16'h5f96;
        src132 <= 16'h59fe;
        src133 <= 16'h44a1;
        src134 <= 16'h211a;
        src135 <= 16'h2a69;
        src136 <= 16'he6f7;
        src137 <= 16'h144;
        src138 <= 16'h6fb2;
        src139 <= 16'he22c;
        src140 <= 16'h9bab;
        src141 <= 16'h5097;
        src142 <= 16'h3514;
        src143 <= 16'hc982;
        src144 <= 16'h18f9;
        src145 <= 16'h9df2;
        src146 <= 16'hf783;
        src147 <= 16'hf12b;
        src148 <= 16'he640;
        src149 <= 16'h70fc;
        src150 <= 16'had8c;
        src151 <= 16'h4e53;
        src152 <= 16'h5cf9;
        src153 <= 16'hbf64;
        src154 <= 16'h113b;
        src155 <= 16'he90;
        src156 <= 16'hd908;
        src157 <= 16'hadb3;
        src158 <= 16'h4745;
        src159 <= 16'h6a6b;
        src160 <= 16'h61f3;
        src161 <= 16'h9298;
        src162 <= 16'h309e;
        src163 <= 16'hfd34;
        src164 <= 16'hc91b;
        src165 <= 16'hf073;
        src166 <= 16'h7a5c;
        src167 <= 16'hdb7c;
        src168 <= 16'h50ec;
        src169 <= 16'h6798;
        src170 <= 16'hd93b;
        src171 <= 16'h39b5;
        src172 <= 16'h791;
        src173 <= 16'h6567;
        src174 <= 16'h5c9d;
        src175 <= 16'h7dd5;
        src176 <= 16'h570b;
        src177 <= 16'he914;
        src178 <= 16'h1d61;
        src179 <= 16'h8569;
        src180 <= 16'h7db7;
        src181 <= 16'h1082;
        src182 <= 16'h242;
        src183 <= 16'h2606;
        src184 <= 16'h451e;
        exp <= 24'h59792c;
        #1
        src0 <= 16'h1395;
        src1 <= 16'hc5d8;
        src2 <= 16'h9ab3;
        src3 <= 16'hff2e;
        src4 <= 16'h50ad;
        src5 <= 16'hc324;
        src6 <= 16'h22df;
        src7 <= 16'h490e;
        src8 <= 16'hbfa2;
        src9 <= 16'h1ba3;
        src10 <= 16'h563c;
        src11 <= 16'hdc17;
        src12 <= 16'ha97a;
        src13 <= 16'hf4fc;
        src14 <= 16'h8001;
        src15 <= 16'hcaa1;
        src16 <= 16'h99fe;
        src17 <= 16'h36da;
        src18 <= 16'h236a;
        src19 <= 16'heefb;
        src20 <= 16'hace;
        src21 <= 16'hedb0;
        src22 <= 16'hacc2;
        src23 <= 16'h777b;
        src24 <= 16'hd7f2;
        src25 <= 16'hc2e5;
        src26 <= 16'h662;
        src27 <= 16'hd80f;
        src28 <= 16'h79b0;
        src29 <= 16'h7f88;
        src30 <= 16'hfd64;
        src31 <= 16'h89ae;
        src32 <= 16'hb486;
        src33 <= 16'h85d5;
        src34 <= 16'h6b58;
        src35 <= 16'h224a;
        src36 <= 16'he409;
        src37 <= 16'had3d;
        src38 <= 16'hdab7;
        src39 <= 16'he504;
        src40 <= 16'hf69f;
        src41 <= 16'h24b1;
        src42 <= 16'h1377;
        src43 <= 16'ha85f;
        src44 <= 16'h5f90;
        src45 <= 16'h544f;
        src46 <= 16'hf265;
        src47 <= 16'hd660;
        src48 <= 16'hf3d5;
        src49 <= 16'h737e;
        src50 <= 16'h8a4e;
        src51 <= 16'hf1b8;
        src52 <= 16'h6605;
        src53 <= 16'hae04;
        src54 <= 16'h5fab;
        src55 <= 16'hc71d;
        src56 <= 16'h7c5;
        src57 <= 16'hac60;
        src58 <= 16'h7c59;
        src59 <= 16'hb371;
        src60 <= 16'h2f59;
        src61 <= 16'h289;
        src62 <= 16'h291d;
        src63 <= 16'he893;
        src64 <= 16'hd58e;
        src65 <= 16'h295;
        src66 <= 16'ha257;
        src67 <= 16'h2c52;
        src68 <= 16'hf289;
        src69 <= 16'h95c0;
        src70 <= 16'h666;
        src71 <= 16'h255e;
        src72 <= 16'hfbf;
        src73 <= 16'h1d56;
        src74 <= 16'h866d;
        src75 <= 16'h65be;
        src76 <= 16'h9c36;
        src77 <= 16'h8974;
        src78 <= 16'hd48b;
        src79 <= 16'h2646;
        src80 <= 16'hde42;
        src81 <= 16'h72f;
        src82 <= 16'h5816;
        src83 <= 16'h7a6b;
        src84 <= 16'h64db;
        src85 <= 16'h381a;
        src86 <= 16'heb7f;
        src87 <= 16'ha6bb;
        src88 <= 16'h5a12;
        src89 <= 16'he664;
        src90 <= 16'h8b23;
        src91 <= 16'h91a5;
        src92 <= 16'hbc3e;
        src93 <= 16'hbba4;
        src94 <= 16'h2be;
        src95 <= 16'hd0;
        src96 <= 16'hf48f;
        src97 <= 16'hf9f2;
        src98 <= 16'h59ca;
        src99 <= 16'h9a47;
        src100 <= 16'h4c29;
        src101 <= 16'h4c43;
        src102 <= 16'h7401;
        src103 <= 16'he502;
        src104 <= 16'h97f3;
        src105 <= 16'he416;
        src106 <= 16'h726d;
        src107 <= 16'hf10a;
        src108 <= 16'hb2e1;
        src109 <= 16'h874b;
        src110 <= 16'hb1a3;
        src111 <= 16'he50e;
        src112 <= 16'he1ba;
        src113 <= 16'h9a61;
        src114 <= 16'hac42;
        src115 <= 16'h77b1;
        src116 <= 16'haa80;
        src117 <= 16'ha41e;
        src118 <= 16'hef05;
        src119 <= 16'h894;
        src120 <= 16'hf63b;
        src121 <= 16'hd363;
        src122 <= 16'ha9de;
        src123 <= 16'h2115;
        src124 <= 16'hcf33;
        src125 <= 16'h24d1;
        src126 <= 16'h7c1b;
        src127 <= 16'h6930;
        src128 <= 16'h8c18;
        src129 <= 16'hab59;
        src130 <= 16'h6b6a;
        src131 <= 16'h13c8;
        src132 <= 16'h563e;
        src133 <= 16'h1473;
        src134 <= 16'hf69f;
        src135 <= 16'h55b7;
        src136 <= 16'h4167;
        src137 <= 16'hec3c;
        src138 <= 16'he9f;
        src139 <= 16'h1c2e;
        src140 <= 16'hf8bf;
        src141 <= 16'heae6;
        src142 <= 16'h52da;
        src143 <= 16'h9a6a;
        src144 <= 16'he07c;
        src145 <= 16'h2ee8;
        src146 <= 16'h359e;
        src147 <= 16'h1fb0;
        src148 <= 16'hb3c;
        src149 <= 16'h7b7;
        src150 <= 16'h5a09;
        src151 <= 16'h240e;
        src152 <= 16'h9228;
        src153 <= 16'he982;
        src154 <= 16'h74d7;
        src155 <= 16'h1a2f;
        src156 <= 16'hfdda;
        src157 <= 16'he8fe;
        src158 <= 16'h37ea;
        src159 <= 16'hd2a6;
        src160 <= 16'hdc34;
        src161 <= 16'hfec;
        src162 <= 16'h2b49;
        src163 <= 16'h4192;
        src164 <= 16'h4bb2;
        src165 <= 16'ha559;
        src166 <= 16'hbd19;
        src167 <= 16'h3334;
        src168 <= 16'h312e;
        src169 <= 16'hf6c6;
        src170 <= 16'h7f9e;
        src171 <= 16'h82db;
        src172 <= 16'h5282;
        src173 <= 16'ha27b;
        src174 <= 16'hab45;
        src175 <= 16'h3b4d;
        src176 <= 16'h1497;
        src177 <= 16'h99c1;
        src178 <= 16'h8616;
        src179 <= 16'h5b0b;
        src180 <= 16'hdf50;
        src181 <= 16'h9235;
        src182 <= 16'hca44;
        src183 <= 16'hf8b9;
        src184 <= 16'hc584;
        exp <= 24'h611544;
        #1
        src0 <= 16'ha427;
        src1 <= 16'h2281;
        src2 <= 16'hc8b3;
        src3 <= 16'h68e2;
        src4 <= 16'h1198;
        src5 <= 16'h121f;
        src6 <= 16'h1998;
        src7 <= 16'hc470;
        src8 <= 16'h9556;
        src9 <= 16'h5e66;
        src10 <= 16'ha0e7;
        src11 <= 16'h9201;
        src12 <= 16'h5cf3;
        src13 <= 16'hd3f7;
        src14 <= 16'h21c4;
        src15 <= 16'h82ec;
        src16 <= 16'h2c9d;
        src17 <= 16'h3651;
        src18 <= 16'h8652;
        src19 <= 16'h26b1;
        src20 <= 16'h7004;
        src21 <= 16'h9d97;
        src22 <= 16'hbc88;
        src23 <= 16'hd3d0;
        src24 <= 16'h1580;
        src25 <= 16'h3b43;
        src26 <= 16'h1ed4;
        src27 <= 16'hae92;
        src28 <= 16'h8f3f;
        src29 <= 16'h7f71;
        src30 <= 16'hb9d0;
        src31 <= 16'h1f10;
        src32 <= 16'h2d86;
        src33 <= 16'h1b34;
        src34 <= 16'h3fcc;
        src35 <= 16'h4cbe;
        src36 <= 16'h4258;
        src37 <= 16'h133e;
        src38 <= 16'h9a9d;
        src39 <= 16'hde99;
        src40 <= 16'h1ac3;
        src41 <= 16'h7baa;
        src42 <= 16'ha515;
        src43 <= 16'h31fc;
        src44 <= 16'h3e0a;
        src45 <= 16'hc6da;
        src46 <= 16'h7f7d;
        src47 <= 16'h46a9;
        src48 <= 16'hc3da;
        src49 <= 16'h24d1;
        src50 <= 16'h5c8d;
        src51 <= 16'h97a4;
        src52 <= 16'hbe79;
        src53 <= 16'h96b3;
        src54 <= 16'he2e0;
        src55 <= 16'h12ef;
        src56 <= 16'h6f4c;
        src57 <= 16'h8ad5;
        src58 <= 16'h7ae0;
        src59 <= 16'h831;
        src60 <= 16'hd0f4;
        src61 <= 16'hbea8;
        src62 <= 16'h91b0;
        src63 <= 16'h2da7;
        src64 <= 16'hd553;
        src65 <= 16'h88;
        src66 <= 16'h5b5e;
        src67 <= 16'h8847;
        src68 <= 16'h561c;
        src69 <= 16'h2a15;
        src70 <= 16'hbf03;
        src71 <= 16'h5ec2;
        src72 <= 16'hb2b7;
        src73 <= 16'h987f;
        src74 <= 16'h910;
        src75 <= 16'hf3c1;
        src76 <= 16'he39f;
        src77 <= 16'hd048;
        src78 <= 16'h38de;
        src79 <= 16'h7c8;
        src80 <= 16'h394a;
        src81 <= 16'h225;
        src82 <= 16'hbfc6;
        src83 <= 16'h4db3;
        src84 <= 16'h64c2;
        src85 <= 16'h8e16;
        src86 <= 16'h76ef;
        src87 <= 16'h6f57;
        src88 <= 16'h9c9a;
        src89 <= 16'hdcc4;
        src90 <= 16'h5654;
        src91 <= 16'he761;
        src92 <= 16'habce;
        src93 <= 16'he0e;
        src94 <= 16'h6930;
        src95 <= 16'h7be5;
        src96 <= 16'hef75;
        src97 <= 16'h3a4d;
        src98 <= 16'h4518;
        src99 <= 16'hff4f;
        src100 <= 16'h94d9;
        src101 <= 16'ha69c;
        src102 <= 16'h4fe2;
        src103 <= 16'h73fb;
        src104 <= 16'h59ba;
        src105 <= 16'hbb3d;
        src106 <= 16'h2379;
        src107 <= 16'hfdf4;
        src108 <= 16'h2ecc;
        src109 <= 16'h59da;
        src110 <= 16'hc94c;
        src111 <= 16'h5710;
        src112 <= 16'hfb92;
        src113 <= 16'h882b;
        src114 <= 16'h6210;
        src115 <= 16'hc8bd;
        src116 <= 16'h6ea1;
        src117 <= 16'hdcf2;
        src118 <= 16'h753e;
        src119 <= 16'hff68;
        src120 <= 16'h24ca;
        src121 <= 16'hacfb;
        src122 <= 16'hd781;
        src123 <= 16'h8deb;
        src124 <= 16'h5805;
        src125 <= 16'h5513;
        src126 <= 16'h1def;
        src127 <= 16'h9ee8;
        src128 <= 16'h314a;
        src129 <= 16'h2b2c;
        src130 <= 16'h8a88;
        src131 <= 16'h99c;
        src132 <= 16'h5110;
        src133 <= 16'h190f;
        src134 <= 16'h2abe;
        src135 <= 16'h4d6c;
        src136 <= 16'hf4d0;
        src137 <= 16'hcb17;
        src138 <= 16'h9aa;
        src139 <= 16'h2b93;
        src140 <= 16'h5a7d;
        src141 <= 16'hd2ea;
        src142 <= 16'hd357;
        src143 <= 16'hb50a;
        src144 <= 16'h9cd9;
        src145 <= 16'hebd7;
        src146 <= 16'h821a;
        src147 <= 16'hf666;
        src148 <= 16'h23b0;
        src149 <= 16'h91c;
        src150 <= 16'h6285;
        src151 <= 16'hae3c;
        src152 <= 16'h5df9;
        src153 <= 16'h7d55;
        src154 <= 16'hbdd3;
        src155 <= 16'h88df;
        src156 <= 16'h7e59;
        src157 <= 16'h5ad1;
        src158 <= 16'h3144;
        src159 <= 16'hd17c;
        src160 <= 16'h54e;
        src161 <= 16'hbfcc;
        src162 <= 16'hd3f1;
        src163 <= 16'hfc17;
        src164 <= 16'h7f5b;
        src165 <= 16'h1f64;
        src166 <= 16'h7a71;
        src167 <= 16'h9ea1;
        src168 <= 16'hd86f;
        src169 <= 16'h4dfa;
        src170 <= 16'hdc1f;
        src171 <= 16'h761d;
        src172 <= 16'h7efb;
        src173 <= 16'h4148;
        src174 <= 16'h3020;
        src175 <= 16'h4bdf;
        src176 <= 16'hec5;
        src177 <= 16'h6753;
        src178 <= 16'h641e;
        src179 <= 16'h6cdf;
        src180 <= 16'h125d;
        src181 <= 16'hb876;
        src182 <= 16'haf4c;
        src183 <= 16'hbb59;
        src184 <= 16'h2e87;
        exp <= 24'h564aa7;
        #1
        src0 <= 16'h9dfb;
        src1 <= 16'h9594;
        src2 <= 16'hd8e7;
        src3 <= 16'he5b3;
        src4 <= 16'h5a00;
        src5 <= 16'he584;
        src6 <= 16'habc9;
        src7 <= 16'h2364;
        src8 <= 16'h5fb5;
        src9 <= 16'h70f4;
        src10 <= 16'hc6c2;
        src11 <= 16'ha387;
        src12 <= 16'h354b;
        src13 <= 16'ha229;
        src14 <= 16'h1b6c;
        src15 <= 16'h7db4;
        src16 <= 16'h62e6;
        src17 <= 16'h9c19;
        src18 <= 16'h912d;
        src19 <= 16'heefc;
        src20 <= 16'h7fe3;
        src21 <= 16'hfc51;
        src22 <= 16'hb5a0;
        src23 <= 16'h536d;
        src24 <= 16'hbfb4;
        src25 <= 16'hf888;
        src26 <= 16'h2b1b;
        src27 <= 16'h3790;
        src28 <= 16'h7482;
        src29 <= 16'h64a0;
        src30 <= 16'hd75d;
        src31 <= 16'h645a;
        src32 <= 16'hbd46;
        src33 <= 16'h2542;
        src34 <= 16'ha0b6;
        src35 <= 16'h24da;
        src36 <= 16'hc2ff;
        src37 <= 16'h9d75;
        src38 <= 16'h5a27;
        src39 <= 16'h2204;
        src40 <= 16'h2df;
        src41 <= 16'hcd61;
        src42 <= 16'h383c;
        src43 <= 16'hbc6e;
        src44 <= 16'hca61;
        src45 <= 16'h3e81;
        src46 <= 16'hd4ec;
        src47 <= 16'hf274;
        src48 <= 16'hb670;
        src49 <= 16'hc204;
        src50 <= 16'h3fc2;
        src51 <= 16'h1908;
        src52 <= 16'hcc12;
        src53 <= 16'hbb57;
        src54 <= 16'hffee;
        src55 <= 16'h64bb;
        src56 <= 16'h32f4;
        src57 <= 16'h55d0;
        src58 <= 16'hfc09;
        src59 <= 16'h60c4;
        src60 <= 16'ha21a;
        src61 <= 16'h62fa;
        src62 <= 16'h7b76;
        src63 <= 16'h8175;
        src64 <= 16'h27af;
        src65 <= 16'hbead;
        src66 <= 16'h106f;
        src67 <= 16'hf39e;
        src68 <= 16'hc087;
        src69 <= 16'h6734;
        src70 <= 16'h7a8f;
        src71 <= 16'h6400;
        src72 <= 16'h6a40;
        src73 <= 16'h2f9c;
        src74 <= 16'h6e3c;
        src75 <= 16'hc175;
        src76 <= 16'h6825;
        src77 <= 16'h7fe2;
        src78 <= 16'h3a04;
        src79 <= 16'h6228;
        src80 <= 16'hf168;
        src81 <= 16'hebd;
        src82 <= 16'habc6;
        src83 <= 16'h5583;
        src84 <= 16'h36ee;
        src85 <= 16'h6abe;
        src86 <= 16'hc295;
        src87 <= 16'h1090;
        src88 <= 16'hdfc1;
        src89 <= 16'h992e;
        src90 <= 16'h405f;
        src91 <= 16'h3115;
        src92 <= 16'hbbac;
        src93 <= 16'hec4a;
        src94 <= 16'heb96;
        src95 <= 16'h6ea3;
        src96 <= 16'h1066;
        src97 <= 16'hcc21;
        src98 <= 16'h77a7;
        src99 <= 16'h362;
        src100 <= 16'h4796;
        src101 <= 16'ha465;
        src102 <= 16'hefca;
        src103 <= 16'hbde8;
        src104 <= 16'hcf94;
        src105 <= 16'hcb1a;
        src106 <= 16'h2d33;
        src107 <= 16'h5af1;
        src108 <= 16'h86bb;
        src109 <= 16'h8a6f;
        src110 <= 16'h4ad2;
        src111 <= 16'h48f7;
        src112 <= 16'h617c;
        src113 <= 16'h4663;
        src114 <= 16'h5331;
        src115 <= 16'ha717;
        src116 <= 16'h548c;
        src117 <= 16'hbf50;
        src118 <= 16'h6937;
        src119 <= 16'h432;
        src120 <= 16'habe1;
        src121 <= 16'ha6ec;
        src122 <= 16'h2d5a;
        src123 <= 16'hd69a;
        src124 <= 16'h3888;
        src125 <= 16'hc490;
        src126 <= 16'h3d89;
        src127 <= 16'h3759;
        src128 <= 16'h20dd;
        src129 <= 16'hc2c;
        src130 <= 16'h403f;
        src131 <= 16'hbf11;
        src132 <= 16'h5e5a;
        src133 <= 16'h6845;
        src134 <= 16'he791;
        src135 <= 16'h553;
        src136 <= 16'h8d20;
        src137 <= 16'h2f63;
        src138 <= 16'hc969;
        src139 <= 16'h2819;
        src140 <= 16'h2ca6;
        src141 <= 16'hb192;
        src142 <= 16'hf633;
        src143 <= 16'he487;
        src144 <= 16'h7833;
        src145 <= 16'hed0c;
        src146 <= 16'habec;
        src147 <= 16'h50f;
        src148 <= 16'h2b20;
        src149 <= 16'he5d5;
        src150 <= 16'h5177;
        src151 <= 16'hb69e;
        src152 <= 16'h46d6;
        src153 <= 16'h7070;
        src154 <= 16'h423b;
        src155 <= 16'hf1d8;
        src156 <= 16'h1829;
        src157 <= 16'h9654;
        src158 <= 16'h7c7;
        src159 <= 16'hb8c8;
        src160 <= 16'h9b82;
        src161 <= 16'h87d0;
        src162 <= 16'h7f14;
        src163 <= 16'hf2b0;
        src164 <= 16'h90a2;
        src165 <= 16'h1823;
        src166 <= 16'h4f80;
        src167 <= 16'hb792;
        src168 <= 16'h1f44;
        src169 <= 16'h2c86;
        src170 <= 16'hf0b6;
        src171 <= 16'h9f99;
        src172 <= 16'hcab9;
        src173 <= 16'hbdc;
        src174 <= 16'h19a;
        src175 <= 16'h756a;
        src176 <= 16'h3a95;
        src177 <= 16'h6514;
        src178 <= 16'h55b9;
        src179 <= 16'h1a4c;
        src180 <= 16'h960e;
        src181 <= 16'hf14c;
        src182 <= 16'h1d3;
        src183 <= 16'ha82c;
        src184 <= 16'h8bcd;
        exp <= 24'h5af1a8;
        #1
        src0 <= 16'h1c32;
        src1 <= 16'h716e;
        src2 <= 16'hfd8;
        src3 <= 16'h77a5;
        src4 <= 16'h80c5;
        src5 <= 16'h4679;
        src6 <= 16'h680d;
        src7 <= 16'hdd9d;
        src8 <= 16'h83e5;
        src9 <= 16'h6f17;
        src10 <= 16'hc74d;
        src11 <= 16'hcc16;
        src12 <= 16'h76cf;
        src13 <= 16'h7b8c;
        src14 <= 16'hf932;
        src15 <= 16'h5532;
        src16 <= 16'h27c7;
        src17 <= 16'h40df;
        src18 <= 16'h69d6;
        src19 <= 16'h72f5;
        src20 <= 16'hdc58;
        src21 <= 16'h5c15;
        src22 <= 16'h4305;
        src23 <= 16'h498b;
        src24 <= 16'hed68;
        src25 <= 16'had75;
        src26 <= 16'h72d4;
        src27 <= 16'h8b03;
        src28 <= 16'h9283;
        src29 <= 16'h1803;
        src30 <= 16'ha61b;
        src31 <= 16'h7b84;
        src32 <= 16'h64e4;
        src33 <= 16'h9999;
        src34 <= 16'he51f;
        src35 <= 16'h2b17;
        src36 <= 16'h42cc;
        src37 <= 16'ha673;
        src38 <= 16'hca23;
        src39 <= 16'h637f;
        src40 <= 16'h6605;
        src41 <= 16'ha4c2;
        src42 <= 16'hc47a;
        src43 <= 16'h8791;
        src44 <= 16'haad0;
        src45 <= 16'h439;
        src46 <= 16'h137c;
        src47 <= 16'he563;
        src48 <= 16'he045;
        src49 <= 16'hb65d;
        src50 <= 16'hcc0c;
        src51 <= 16'h6099;
        src52 <= 16'h3a9b;
        src53 <= 16'h8663;
        src54 <= 16'h851b;
        src55 <= 16'h7471;
        src56 <= 16'h732;
        src57 <= 16'hc72f;
        src58 <= 16'h6f84;
        src59 <= 16'hc412;
        src60 <= 16'hc29;
        src61 <= 16'h437c;
        src62 <= 16'he68c;
        src63 <= 16'he316;
        src64 <= 16'hd518;
        src65 <= 16'h577f;
        src66 <= 16'h352c;
        src67 <= 16'h9c55;
        src68 <= 16'h7e24;
        src69 <= 16'h9ce6;
        src70 <= 16'hdd76;
        src71 <= 16'h4363;
        src72 <= 16'hb419;
        src73 <= 16'hc7ad;
        src74 <= 16'h5616;
        src75 <= 16'hfdff;
        src76 <= 16'h16d8;
        src77 <= 16'h70a;
        src78 <= 16'hea8f;
        src79 <= 16'h1225;
        src80 <= 16'hb43f;
        src81 <= 16'h35d6;
        src82 <= 16'h3c00;
        src83 <= 16'h28e5;
        src84 <= 16'h6bba;
        src85 <= 16'h81ac;
        src86 <= 16'h9a90;
        src87 <= 16'ha906;
        src88 <= 16'h7c40;
        src89 <= 16'h597f;
        src90 <= 16'h916f;
        src91 <= 16'hed37;
        src92 <= 16'h9e6d;
        src93 <= 16'he973;
        src94 <= 16'h8c24;
        src95 <= 16'h4b67;
        src96 <= 16'h6e21;
        src97 <= 16'ha4dd;
        src98 <= 16'h230c;
        src99 <= 16'h4b10;
        src100 <= 16'hf064;
        src101 <= 16'h8c68;
        src102 <= 16'ha556;
        src103 <= 16'h1b24;
        src104 <= 16'h14e7;
        src105 <= 16'hc33c;
        src106 <= 16'hed47;
        src107 <= 16'h6bd1;
        src108 <= 16'hcaea;
        src109 <= 16'h7d32;
        src110 <= 16'h78de;
        src111 <= 16'h67bb;
        src112 <= 16'h8797;
        src113 <= 16'hed43;
        src114 <= 16'he569;
        src115 <= 16'h4cf8;
        src116 <= 16'hd12d;
        src117 <= 16'ha1e7;
        src118 <= 16'hacf4;
        src119 <= 16'h76e1;
        src120 <= 16'hc67b;
        src121 <= 16'h6bd0;
        src122 <= 16'hbf0c;
        src123 <= 16'h84ab;
        src124 <= 16'he527;
        src125 <= 16'h8cbd;
        src126 <= 16'h8871;
        src127 <= 16'hddc5;
        src128 <= 16'h9a9f;
        src129 <= 16'h3030;
        src130 <= 16'h8fdc;
        src131 <= 16'h376b;
        src132 <= 16'hbb69;
        src133 <= 16'hc605;
        src134 <= 16'h1daa;
        src135 <= 16'h410b;
        src136 <= 16'hece3;
        src137 <= 16'hf692;
        src138 <= 16'had0d;
        src139 <= 16'h44d7;
        src140 <= 16'h973c;
        src141 <= 16'h9dbf;
        src142 <= 16'h1f8d;
        src143 <= 16'haf3b;
        src144 <= 16'h7543;
        src145 <= 16'he32;
        src146 <= 16'h342;
        src147 <= 16'hbefa;
        src148 <= 16'h9a33;
        src149 <= 16'hd24a;
        src150 <= 16'h2ca6;
        src151 <= 16'hef40;
        src152 <= 16'hafe8;
        src153 <= 16'h1ccd;
        src154 <= 16'h83d3;
        src155 <= 16'hcaf8;
        src156 <= 16'h1128;
        src157 <= 16'haa84;
        src158 <= 16'ha6fa;
        src159 <= 16'hd802;
        src160 <= 16'hf99c;
        src161 <= 16'h23c;
        src162 <= 16'hb727;
        src163 <= 16'h17ec;
        src164 <= 16'hdad9;
        src165 <= 16'h15bd;
        src166 <= 16'h120c;
        src167 <= 16'hf54f;
        src168 <= 16'ha4ee;
        src169 <= 16'h589f;
        src170 <= 16'h75ee;
        src171 <= 16'h9f3d;
        src172 <= 16'hcf07;
        src173 <= 16'he47b;
        src174 <= 16'hdb2b;
        src175 <= 16'h79e7;
        src176 <= 16'hd25a;
        src177 <= 16'h5eaa;
        src178 <= 16'h791;
        src179 <= 16'h7511;
        src180 <= 16'hf02b;
        src181 <= 16'h1267;
        src182 <= 16'h44a3;
        src183 <= 16'hb30b;
        src184 <= 16'h90c4;
        exp <= 24'h6098ec;
        #1
        src0 <= 16'h30ca;
        src1 <= 16'hab42;
        src2 <= 16'h8e46;
        src3 <= 16'hc80b;
        src4 <= 16'hc46a;
        src5 <= 16'hf5f9;
        src6 <= 16'h3d99;
        src7 <= 16'hfad;
        src8 <= 16'h4fb4;
        src9 <= 16'hae81;
        src10 <= 16'he6a1;
        src11 <= 16'hdb51;
        src12 <= 16'h4d0a;
        src13 <= 16'h1b41;
        src14 <= 16'h7aeb;
        src15 <= 16'haf0b;
        src16 <= 16'hd669;
        src17 <= 16'h212e;
        src18 <= 16'h8bba;
        src19 <= 16'h7b45;
        src20 <= 16'h2f13;
        src21 <= 16'h764;
        src22 <= 16'h589a;
        src23 <= 16'h77ea;
        src24 <= 16'hf326;
        src25 <= 16'h97ff;
        src26 <= 16'h7c9c;
        src27 <= 16'h9981;
        src28 <= 16'hbd80;
        src29 <= 16'h1308;
        src30 <= 16'h88c;
        src31 <= 16'h7fce;
        src32 <= 16'hbb6f;
        src33 <= 16'h846f;
        src34 <= 16'hfc98;
        src35 <= 16'h480c;
        src36 <= 16'h8b06;
        src37 <= 16'haf1c;
        src38 <= 16'haa90;
        src39 <= 16'hd255;
        src40 <= 16'h7b38;
        src41 <= 16'h32a7;
        src42 <= 16'h23d0;
        src43 <= 16'he0a6;
        src44 <= 16'hf897;
        src45 <= 16'h1e8b;
        src46 <= 16'h4185;
        src47 <= 16'h68a1;
        src48 <= 16'hb090;
        src49 <= 16'h35a6;
        src50 <= 16'h9f11;
        src51 <= 16'h7da8;
        src52 <= 16'hb2bf;
        src53 <= 16'hdd4a;
        src54 <= 16'hd265;
        src55 <= 16'hdad9;
        src56 <= 16'ha0c5;
        src57 <= 16'h4542;
        src58 <= 16'h1a88;
        src59 <= 16'hd7d;
        src60 <= 16'he322;
        src61 <= 16'h47a2;
        src62 <= 16'h48e;
        src63 <= 16'h8c0b;
        src64 <= 16'he198;
        src65 <= 16'hb6d6;
        src66 <= 16'h676b;
        src67 <= 16'h32d5;
        src68 <= 16'h177;
        src69 <= 16'h4141;
        src70 <= 16'h10cb;
        src71 <= 16'hc1e7;
        src72 <= 16'he219;
        src73 <= 16'h87e7;
        src74 <= 16'hf589;
        src75 <= 16'h13ea;
        src76 <= 16'h5e51;
        src77 <= 16'hcc86;
        src78 <= 16'hae7c;
        src79 <= 16'h2a1f;
        src80 <= 16'h2b99;
        src81 <= 16'hdf;
        src82 <= 16'h602b;
        src83 <= 16'h9027;
        src84 <= 16'hfae4;
        src85 <= 16'hc840;
        src86 <= 16'he010;
        src87 <= 16'hba32;
        src88 <= 16'h3e23;
        src89 <= 16'hf515;
        src90 <= 16'hbcf1;
        src91 <= 16'h4ba5;
        src92 <= 16'he87b;
        src93 <= 16'h7488;
        src94 <= 16'he8ad;
        src95 <= 16'hcd53;
        src96 <= 16'h6c46;
        src97 <= 16'hbb98;
        src98 <= 16'h7131;
        src99 <= 16'h8ac9;
        src100 <= 16'he4bc;
        src101 <= 16'h4643;
        src102 <= 16'hac4c;
        src103 <= 16'h1184;
        src104 <= 16'hf9b2;
        src105 <= 16'heca0;
        src106 <= 16'h62af;
        src107 <= 16'heb0a;
        src108 <= 16'hebd9;
        src109 <= 16'h1682;
        src110 <= 16'h69fc;
        src111 <= 16'h372e;
        src112 <= 16'h2533;
        src113 <= 16'h4c0c;
        src114 <= 16'h800d;
        src115 <= 16'he91e;
        src116 <= 16'hc4f9;
        src117 <= 16'hae93;
        src118 <= 16'ha76d;
        src119 <= 16'hf349;
        src120 <= 16'hf818;
        src121 <= 16'heab5;
        src122 <= 16'h2727;
        src123 <= 16'h350b;
        src124 <= 16'hffbd;
        src125 <= 16'hece2;
        src126 <= 16'hca77;
        src127 <= 16'h42f4;
        src128 <= 16'h6601;
        src129 <= 16'h1fc6;
        src130 <= 16'h2fd4;
        src131 <= 16'h719c;
        src132 <= 16'h5c8e;
        src133 <= 16'h6285;
        src134 <= 16'hd703;
        src135 <= 16'h46d4;
        src136 <= 16'h4217;
        src137 <= 16'h408f;
        src138 <= 16'h2e8e;
        src139 <= 16'hb4ba;
        src140 <= 16'h9470;
        src141 <= 16'h2e74;
        src142 <= 16'h374d;
        src143 <= 16'hcf41;
        src144 <= 16'h7cc9;
        src145 <= 16'h15d6;
        src146 <= 16'h842a;
        src147 <= 16'h82c0;
        src148 <= 16'hc226;
        src149 <= 16'h9d3e;
        src150 <= 16'hc1f;
        src151 <= 16'h10f6;
        src152 <= 16'he8a;
        src153 <= 16'hcffa;
        src154 <= 16'h1311;
        src155 <= 16'h3c75;
        src156 <= 16'hb43a;
        src157 <= 16'h42d9;
        src158 <= 16'he0c6;
        src159 <= 16'h7666;
        src160 <= 16'h6f17;
        src161 <= 16'h5fd;
        src162 <= 16'h9b3;
        src163 <= 16'h4bb4;
        src164 <= 16'h7eab;
        src165 <= 16'h5bb;
        src166 <= 16'h5cd0;
        src167 <= 16'h332a;
        src168 <= 16'h6d28;
        src169 <= 16'he05d;
        src170 <= 16'h418a;
        src171 <= 16'h3cb;
        src172 <= 16'hbed9;
        src173 <= 16'h8123;
        src174 <= 16'h1cb;
        src175 <= 16'hc0dd;
        src176 <= 16'hc04b;
        src177 <= 16'hbeb6;
        src178 <= 16'h669;
        src179 <= 16'h8ac8;
        src180 <= 16'he021;
        src181 <= 16'hbfb2;
        src182 <= 16'hec2;
        src183 <= 16'hc835;
        src184 <= 16'h9f4f;
        exp <= 24'h5c3342;
        #1
        src0 <= 16'h9355;
        src1 <= 16'ha1c4;
        src2 <= 16'hf82b;
        src3 <= 16'hbee3;
        src4 <= 16'h33fc;
        src5 <= 16'hb3c5;
        src6 <= 16'h41ec;
        src7 <= 16'h88f6;
        src8 <= 16'he996;
        src9 <= 16'hf075;
        src10 <= 16'h9f5c;
        src11 <= 16'h1921;
        src12 <= 16'he3ec;
        src13 <= 16'h7629;
        src14 <= 16'h501b;
        src15 <= 16'hc15c;
        src16 <= 16'h14dc;
        src17 <= 16'h64c3;
        src18 <= 16'hae83;
        src19 <= 16'hbfc7;
        src20 <= 16'h355b;
        src21 <= 16'h283c;
        src22 <= 16'h2567;
        src23 <= 16'h43a1;
        src24 <= 16'h6008;
        src25 <= 16'h4d3a;
        src26 <= 16'hf60a;
        src27 <= 16'h90a4;
        src28 <= 16'hdcd4;
        src29 <= 16'h8a69;
        src30 <= 16'hfb35;
        src31 <= 16'h865e;
        src32 <= 16'h8b34;
        src33 <= 16'h98a7;
        src34 <= 16'h8be3;
        src35 <= 16'h1f2a;
        src36 <= 16'ha097;
        src37 <= 16'hb80e;
        src38 <= 16'h7552;
        src39 <= 16'h260a;
        src40 <= 16'h1858;
        src41 <= 16'h898c;
        src42 <= 16'haa73;
        src43 <= 16'hd08d;
        src44 <= 16'ha37d;
        src45 <= 16'h2a6b;
        src46 <= 16'hcbba;
        src47 <= 16'h6281;
        src48 <= 16'h4e42;
        src49 <= 16'h9bff;
        src50 <= 16'h862d;
        src51 <= 16'ha4b;
        src52 <= 16'h6462;
        src53 <= 16'ha938;
        src54 <= 16'ha81a;
        src55 <= 16'hd42d;
        src56 <= 16'h4df8;
        src57 <= 16'h6712;
        src58 <= 16'he073;
        src59 <= 16'h1cda;
        src60 <= 16'h3812;
        src61 <= 16'hdb55;
        src62 <= 16'hce72;
        src63 <= 16'h5733;
        src64 <= 16'h86ec;
        src65 <= 16'h5a0d;
        src66 <= 16'hf0d9;
        src67 <= 16'hf1d9;
        src68 <= 16'h7ded;
        src69 <= 16'h2848;
        src70 <= 16'hcd60;
        src71 <= 16'h5ff5;
        src72 <= 16'h94dc;
        src73 <= 16'h7e29;
        src74 <= 16'hbb9f;
        src75 <= 16'h5a37;
        src76 <= 16'h1cc;
        src77 <= 16'h48ab;
        src78 <= 16'h32ff;
        src79 <= 16'ha8f6;
        src80 <= 16'h36e3;
        src81 <= 16'hf1b;
        src82 <= 16'hf9a8;
        src83 <= 16'h9d11;
        src84 <= 16'h7582;
        src85 <= 16'h85ee;
        src86 <= 16'h7c5c;
        src87 <= 16'hcaa8;
        src88 <= 16'h129b;
        src89 <= 16'h6e7b;
        src90 <= 16'h1e18;
        src91 <= 16'h5e24;
        src92 <= 16'h8142;
        src93 <= 16'h6c25;
        src94 <= 16'h24d1;
        src95 <= 16'hec1f;
        src96 <= 16'h6b80;
        src97 <= 16'h9e8c;
        src98 <= 16'h2089;
        src99 <= 16'h9f59;
        src100 <= 16'hd47e;
        src101 <= 16'hf99;
        src102 <= 16'hfbc7;
        src103 <= 16'h9413;
        src104 <= 16'h5365;
        src105 <= 16'hc86;
        src106 <= 16'h65e8;
        src107 <= 16'h59bb;
        src108 <= 16'h88b8;
        src109 <= 16'h4811;
        src110 <= 16'hd500;
        src111 <= 16'ha0ff;
        src112 <= 16'h280d;
        src113 <= 16'h3077;
        src114 <= 16'hefe;
        src115 <= 16'h10dc;
        src116 <= 16'hcef5;
        src117 <= 16'h18f7;
        src118 <= 16'hc1b8;
        src119 <= 16'h3419;
        src120 <= 16'h144c;
        src121 <= 16'heec2;
        src122 <= 16'ha73a;
        src123 <= 16'hbae8;
        src124 <= 16'h2540;
        src125 <= 16'h59cd;
        src126 <= 16'hbddb;
        src127 <= 16'h4bc9;
        src128 <= 16'h6806;
        src129 <= 16'haec5;
        src130 <= 16'h6a14;
        src131 <= 16'h18cf;
        src132 <= 16'hf5da;
        src133 <= 16'h520a;
        src134 <= 16'h1de3;
        src135 <= 16'h3e6b;
        src136 <= 16'h6b73;
        src137 <= 16'ha16e;
        src138 <= 16'h2409;
        src139 <= 16'h2a5b;
        src140 <= 16'ha1d0;
        src141 <= 16'hf735;
        src142 <= 16'h6df8;
        src143 <= 16'hdbc7;
        src144 <= 16'hdcde;
        src145 <= 16'h187d;
        src146 <= 16'hedd7;
        src147 <= 16'h79e;
        src148 <= 16'h25d8;
        src149 <= 16'hff16;
        src150 <= 16'h9c4f;
        src151 <= 16'hb3ce;
        src152 <= 16'h6f3f;
        src153 <= 16'he298;
        src154 <= 16'h1f2b;
        src155 <= 16'h1693;
        src156 <= 16'h7b44;
        src157 <= 16'he32a;
        src158 <= 16'h42cd;
        src159 <= 16'hfd8a;
        src160 <= 16'h642d;
        src161 <= 16'hf9b6;
        src162 <= 16'hb175;
        src163 <= 16'h4613;
        src164 <= 16'h2bcf;
        src165 <= 16'h61bd;
        src166 <= 16'h468b;
        src167 <= 16'h2d04;
        src168 <= 16'h11f0;
        src169 <= 16'h1c;
        src170 <= 16'h4aab;
        src171 <= 16'hffee;
        src172 <= 16'h12e7;
        src173 <= 16'hdcf;
        src174 <= 16'h4144;
        src175 <= 16'h9578;
        src176 <= 16'h41c0;
        src177 <= 16'h8e7b;
        src178 <= 16'h9c9d;
        src179 <= 16'hf1b2;
        src180 <= 16'h9af4;
        src181 <= 16'h8c0f;
        src182 <= 16'h6909;
        src183 <= 16'h3342;
        src184 <= 16'hb9fd;
        exp <= 24'h58a624;
        #1
        src0 <= 16'hf4eb;
        src1 <= 16'h5ec;
        src2 <= 16'ha21e;
        src3 <= 16'h7b3c;
        src4 <= 16'h9c96;
        src5 <= 16'hfc35;
        src6 <= 16'h240;
        src7 <= 16'h9ee8;
        src8 <= 16'h58ca;
        src9 <= 16'hfc30;
        src10 <= 16'h842f;
        src11 <= 16'h5d84;
        src12 <= 16'hca88;
        src13 <= 16'h1436;
        src14 <= 16'hac63;
        src15 <= 16'hd7cf;
        src16 <= 16'h8732;
        src17 <= 16'hcb35;
        src18 <= 16'hc59e;
        src19 <= 16'hfd31;
        src20 <= 16'h597a;
        src21 <= 16'hc595;
        src22 <= 16'hd027;
        src23 <= 16'h6154;
        src24 <= 16'h7966;
        src25 <= 16'h12ce;
        src26 <= 16'hc246;
        src27 <= 16'hf048;
        src28 <= 16'h1dd8;
        src29 <= 16'he679;
        src30 <= 16'he571;
        src31 <= 16'h864a;
        src32 <= 16'h1774;
        src33 <= 16'hcb6;
        src34 <= 16'h9aea;
        src35 <= 16'hc008;
        src36 <= 16'h3902;
        src37 <= 16'h5f7c;
        src38 <= 16'h476c;
        src39 <= 16'h65c6;
        src40 <= 16'h2f0d;
        src41 <= 16'hd25a;
        src42 <= 16'h8e3d;
        src43 <= 16'h3760;
        src44 <= 16'h1c55;
        src45 <= 16'ha441;
        src46 <= 16'h2307;
        src47 <= 16'h60c8;
        src48 <= 16'h182;
        src49 <= 16'hfe20;
        src50 <= 16'h8cf4;
        src51 <= 16'ha831;
        src52 <= 16'h5345;
        src53 <= 16'hdd76;
        src54 <= 16'h6edd;
        src55 <= 16'h68a9;
        src56 <= 16'h3bdb;
        src57 <= 16'h8215;
        src58 <= 16'h9a0e;
        src59 <= 16'he09e;
        src60 <= 16'h2c21;
        src61 <= 16'hc1da;
        src62 <= 16'hcdab;
        src63 <= 16'h5b9c;
        src64 <= 16'he1f5;
        src65 <= 16'haf71;
        src66 <= 16'hb586;
        src67 <= 16'h5db0;
        src68 <= 16'h2a19;
        src69 <= 16'hd6c1;
        src70 <= 16'h121d;
        src71 <= 16'hdbfc;
        src72 <= 16'ha361;
        src73 <= 16'h30c5;
        src74 <= 16'h75c0;
        src75 <= 16'h864b;
        src76 <= 16'hfbbd;
        src77 <= 16'ha0bf;
        src78 <= 16'h606c;
        src79 <= 16'h8013;
        src80 <= 16'h6145;
        src81 <= 16'hc41;
        src82 <= 16'h30a1;
        src83 <= 16'h7819;
        src84 <= 16'h4a05;
        src85 <= 16'h527d;
        src86 <= 16'h8d74;
        src87 <= 16'h3c65;
        src88 <= 16'hd860;
        src89 <= 16'h8d41;
        src90 <= 16'he555;
        src91 <= 16'h724c;
        src92 <= 16'h4dfd;
        src93 <= 16'h575b;
        src94 <= 16'h42eb;
        src95 <= 16'he8d6;
        src96 <= 16'hb016;
        src97 <= 16'h829b;
        src98 <= 16'h653f;
        src99 <= 16'h2c53;
        src100 <= 16'h8e34;
        src101 <= 16'hd335;
        src102 <= 16'ha894;
        src103 <= 16'h9ce7;
        src104 <= 16'hb311;
        src105 <= 16'h783f;
        src106 <= 16'h1720;
        src107 <= 16'hce7d;
        src108 <= 16'h47b2;
        src109 <= 16'hc389;
        src110 <= 16'h13fa;
        src111 <= 16'ha5ef;
        src112 <= 16'h35fd;
        src113 <= 16'hc9d5;
        src114 <= 16'h9135;
        src115 <= 16'h1bdd;
        src116 <= 16'h344;
        src117 <= 16'h4fc4;
        src118 <= 16'hd602;
        src119 <= 16'h42a3;
        src120 <= 16'h450e;
        src121 <= 16'hb87e;
        src122 <= 16'h7589;
        src123 <= 16'h2f74;
        src124 <= 16'h8215;
        src125 <= 16'h55b5;
        src126 <= 16'h1bf5;
        src127 <= 16'h880a;
        src128 <= 16'h4b73;
        src129 <= 16'h5352;
        src130 <= 16'hea51;
        src131 <= 16'ha44d;
        src132 <= 16'hc1d0;
        src133 <= 16'hd823;
        src134 <= 16'he0dd;
        src135 <= 16'hd667;
        src136 <= 16'h7ff4;
        src137 <= 16'h43b1;
        src138 <= 16'h67c6;
        src139 <= 16'h514b;
        src140 <= 16'hae09;
        src141 <= 16'h191f;
        src142 <= 16'h933;
        src143 <= 16'h54c8;
        src144 <= 16'h9876;
        src145 <= 16'hc4db;
        src146 <= 16'h88fb;
        src147 <= 16'h96ac;
        src148 <= 16'hbc05;
        src149 <= 16'h40e;
        src150 <= 16'hab0a;
        src151 <= 16'h8b96;
        src152 <= 16'h9b96;
        src153 <= 16'h5de;
        src154 <= 16'h5af5;
        src155 <= 16'h368b;
        src156 <= 16'h96d4;
        src157 <= 16'h8460;
        src158 <= 16'hc51a;
        src159 <= 16'h45ef;
        src160 <= 16'hf65c;
        src161 <= 16'h32d0;
        src162 <= 16'hcb5f;
        src163 <= 16'haefa;
        src164 <= 16'h835e;
        src165 <= 16'hf3e7;
        src166 <= 16'hf22;
        src167 <= 16'h8a30;
        src168 <= 16'hcd90;
        src169 <= 16'hf04b;
        src170 <= 16'hcd73;
        src171 <= 16'h1e4;
        src172 <= 16'h20c2;
        src173 <= 16'hbfb8;
        src174 <= 16'h90b9;
        src175 <= 16'hbc1;
        src176 <= 16'h276f;
        src177 <= 16'h59eb;
        src178 <= 16'hc153;
        src179 <= 16'he1ec;
        src180 <= 16'h61e6;
        src181 <= 16'h8c4f;
        src182 <= 16'h5736;
        src183 <= 16'h4ff0;
        src184 <= 16'hb964;
        exp <= 24'h5ce01f;
        #1
        src0 <= 16'h8be5;
        src1 <= 16'h6de3;
        src2 <= 16'hdddd;
        src3 <= 16'h7439;
        src4 <= 16'hee74;
        src5 <= 16'h9e5d;
        src6 <= 16'h8502;
        src7 <= 16'hd989;
        src8 <= 16'hb93d;
        src9 <= 16'ha630;
        src10 <= 16'h2aaf;
        src11 <= 16'heab9;
        src12 <= 16'hdbfd;
        src13 <= 16'h9f14;
        src14 <= 16'h5646;
        src15 <= 16'ha930;
        src16 <= 16'hba09;
        src17 <= 16'h752d;
        src18 <= 16'he2ad;
        src19 <= 16'h4791;
        src20 <= 16'h1df5;
        src21 <= 16'he1b2;
        src22 <= 16'hc2af;
        src23 <= 16'h6a89;
        src24 <= 16'hbe64;
        src25 <= 16'h828b;
        src26 <= 16'h61bc;
        src27 <= 16'heef0;
        src28 <= 16'h519b;
        src29 <= 16'h411d;
        src30 <= 16'h5713;
        src31 <= 16'h9229;
        src32 <= 16'h4f9a;
        src33 <= 16'h2cdc;
        src34 <= 16'hc76c;
        src35 <= 16'hc05a;
        src36 <= 16'h87c4;
        src37 <= 16'h6806;
        src38 <= 16'h8270;
        src39 <= 16'hc2b4;
        src40 <= 16'h5055;
        src41 <= 16'h53c9;
        src42 <= 16'h220c;
        src43 <= 16'h9380;
        src44 <= 16'h421b;
        src45 <= 16'h537f;
        src46 <= 16'hab5c;
        src47 <= 16'h9421;
        src48 <= 16'h4594;
        src49 <= 16'h3bd2;
        src50 <= 16'h423;
        src51 <= 16'hb39a;
        src52 <= 16'h1781;
        src53 <= 16'hbde6;
        src54 <= 16'h6606;
        src55 <= 16'h467e;
        src56 <= 16'hfc1e;
        src57 <= 16'hf4db;
        src58 <= 16'he33c;
        src59 <= 16'h6243;
        src60 <= 16'hc1e5;
        src61 <= 16'h797c;
        src62 <= 16'h22ee;
        src63 <= 16'hbb47;
        src64 <= 16'had9d;
        src65 <= 16'h215c;
        src66 <= 16'h1d05;
        src67 <= 16'h364;
        src68 <= 16'h779d;
        src69 <= 16'hdbad;
        src70 <= 16'h8c8a;
        src71 <= 16'h7d5d;
        src72 <= 16'hde70;
        src73 <= 16'h1e4b;
        src74 <= 16'h3132;
        src75 <= 16'ha2f1;
        src76 <= 16'hb40a;
        src77 <= 16'h3420;
        src78 <= 16'h1096;
        src79 <= 16'h9f80;
        src80 <= 16'h5c0;
        src81 <= 16'h7291;
        src82 <= 16'h6a0d;
        src83 <= 16'hc4b1;
        src84 <= 16'h4a34;
        src85 <= 16'hf031;
        src86 <= 16'h3c39;
        src87 <= 16'hba71;
        src88 <= 16'h67b;
        src89 <= 16'h6fc;
        src90 <= 16'h6683;
        src91 <= 16'h866;
        src92 <= 16'h462c;
        src93 <= 16'hf701;
        src94 <= 16'h95f9;
        src95 <= 16'h7167;
        src96 <= 16'h6754;
        src97 <= 16'hbf4a;
        src98 <= 16'hd4be;
        src99 <= 16'h2ef5;
        src100 <= 16'hb9b2;
        src101 <= 16'h2e97;
        src102 <= 16'h9514;
        src103 <= 16'h6ce4;
        src104 <= 16'h3ce0;
        src105 <= 16'hc041;
        src106 <= 16'h1f6a;
        src107 <= 16'h18a2;
        src108 <= 16'h6565;
        src109 <= 16'h122c;
        src110 <= 16'h2705;
        src111 <= 16'h2d0a;
        src112 <= 16'h4973;
        src113 <= 16'h2051;
        src114 <= 16'h550f;
        src115 <= 16'hde5a;
        src116 <= 16'h433b;
        src117 <= 16'h7b9f;
        src118 <= 16'he3d5;
        src119 <= 16'h71bc;
        src120 <= 16'h58b4;
        src121 <= 16'h1d19;
        src122 <= 16'hf9fe;
        src123 <= 16'h6c8;
        src124 <= 16'h5e8;
        src125 <= 16'h6298;
        src126 <= 16'h39ef;
        src127 <= 16'he18f;
        src128 <= 16'h5d95;
        src129 <= 16'h6511;
        src130 <= 16'h3932;
        src131 <= 16'h70af;
        src132 <= 16'h7b5a;
        src133 <= 16'h765c;
        src134 <= 16'h3197;
        src135 <= 16'h8ceb;
        src136 <= 16'h128;
        src137 <= 16'h9ab4;
        src138 <= 16'h4bd5;
        src139 <= 16'hdb89;
        src140 <= 16'hcf5a;
        src141 <= 16'h5e46;
        src142 <= 16'h7520;
        src143 <= 16'h9a7c;
        src144 <= 16'h7e98;
        src145 <= 16'hdddc;
        src146 <= 16'hcbb;
        src147 <= 16'h6dd3;
        src148 <= 16'h856d;
        src149 <= 16'h3452;
        src150 <= 16'h7196;
        src151 <= 16'h146d;
        src152 <= 16'h8d23;
        src153 <= 16'h1b12;
        src154 <= 16'h2a78;
        src155 <= 16'h7a1f;
        src156 <= 16'h9b40;
        src157 <= 16'h897e;
        src158 <= 16'h347b;
        src159 <= 16'hbfb5;
        src160 <= 16'h718e;
        src161 <= 16'h2a52;
        src162 <= 16'h6be0;
        src163 <= 16'h8ad8;
        src164 <= 16'hb82;
        src165 <= 16'hd794;
        src166 <= 16'h130;
        src167 <= 16'hc9cd;
        src168 <= 16'h122;
        src169 <= 16'h67e3;
        src170 <= 16'hc1dc;
        src171 <= 16'h1e43;
        src172 <= 16'h81a7;
        src173 <= 16'h5415;
        src174 <= 16'h5b3c;
        src175 <= 16'h156f;
        src176 <= 16'hf09f;
        src177 <= 16'hc548;
        src178 <= 16'h41d2;
        src179 <= 16'hfd20;
        src180 <= 16'h6a44;
        src181 <= 16'hb751;
        src182 <= 16'hc996;
        src183 <= 16'hec05;
        src184 <= 16'h88c8;
        exp <= 24'h55fc7d;
        #1
        src0 <= 16'h4a28;
        src1 <= 16'h1903;
        src2 <= 16'h3086;
        src3 <= 16'h5d1d;
        src4 <= 16'hb7ba;
        src5 <= 16'h1cfa;
        src6 <= 16'h8cb2;
        src7 <= 16'h68a9;
        src8 <= 16'he9b5;
        src9 <= 16'h8c88;
        src10 <= 16'hd049;
        src11 <= 16'h4ca7;
        src12 <= 16'h1eec;
        src13 <= 16'ha2f1;
        src14 <= 16'hd8ae;
        src15 <= 16'h1673;
        src16 <= 16'h6bdd;
        src17 <= 16'he494;
        src18 <= 16'h74e3;
        src19 <= 16'h62d4;
        src20 <= 16'h9852;
        src21 <= 16'h4418;
        src22 <= 16'hb389;
        src23 <= 16'h2469;
        src24 <= 16'he489;
        src25 <= 16'h9933;
        src26 <= 16'hc7d0;
        src27 <= 16'h2267;
        src28 <= 16'hb61c;
        src29 <= 16'h358a;
        src30 <= 16'h1388;
        src31 <= 16'h78aa;
        src32 <= 16'he143;
        src33 <= 16'h167f;
        src34 <= 16'h1beb;
        src35 <= 16'h3ce8;
        src36 <= 16'h7408;
        src37 <= 16'hae39;
        src38 <= 16'h828;
        src39 <= 16'h8035;
        src40 <= 16'h546f;
        src41 <= 16'h3894;
        src42 <= 16'hc60d;
        src43 <= 16'hb6ab;
        src44 <= 16'h72ab;
        src45 <= 16'h8c44;
        src46 <= 16'haee4;
        src47 <= 16'hcd00;
        src48 <= 16'h45e1;
        src49 <= 16'hab5f;
        src50 <= 16'hdcf2;
        src51 <= 16'h9eac;
        src52 <= 16'h9930;
        src53 <= 16'hf3d0;
        src54 <= 16'ha90b;
        src55 <= 16'h7631;
        src56 <= 16'h2d7c;
        src57 <= 16'hd3f3;
        src58 <= 16'hd3bc;
        src59 <= 16'hbe16;
        src60 <= 16'h952f;
        src61 <= 16'hc000;
        src62 <= 16'ha3d2;
        src63 <= 16'ha34b;
        src64 <= 16'hdcb0;
        src65 <= 16'h1c02;
        src66 <= 16'hefeb;
        src67 <= 16'hdbe5;
        src68 <= 16'hea55;
        src69 <= 16'hcf3;
        src70 <= 16'h8814;
        src71 <= 16'h75da;
        src72 <= 16'hefe8;
        src73 <= 16'h215;
        src74 <= 16'h1e79;
        src75 <= 16'h835f;
        src76 <= 16'hec12;
        src77 <= 16'hf6f;
        src78 <= 16'h7acf;
        src79 <= 16'h4ae;
        src80 <= 16'h8a1;
        src81 <= 16'h3c72;
        src82 <= 16'hbc73;
        src83 <= 16'he356;
        src84 <= 16'hd27;
        src85 <= 16'hcfdc;
        src86 <= 16'h38db;
        src87 <= 16'hdbb6;
        src88 <= 16'h7cb;
        src89 <= 16'h49d2;
        src90 <= 16'h4766;
        src91 <= 16'h5249;
        src92 <= 16'ha34b;
        src93 <= 16'h654f;
        src94 <= 16'h2620;
        src95 <= 16'hfa67;
        src96 <= 16'h5879;
        src97 <= 16'h2ba6;
        src98 <= 16'hcbc0;
        src99 <= 16'h73bf;
        src100 <= 16'h6089;
        src101 <= 16'h5cce;
        src102 <= 16'he63e;
        src103 <= 16'h60d3;
        src104 <= 16'hdb75;
        src105 <= 16'ha579;
        src106 <= 16'h8de8;
        src107 <= 16'h3d27;
        src108 <= 16'hefd6;
        src109 <= 16'h4b9;
        src110 <= 16'hf9de;
        src111 <= 16'hc923;
        src112 <= 16'h2f40;
        src113 <= 16'hb7fa;
        src114 <= 16'hf057;
        src115 <= 16'h30b8;
        src116 <= 16'h7ca6;
        src117 <= 16'ha154;
        src118 <= 16'hf96c;
        src119 <= 16'h5fc4;
        src120 <= 16'he3d1;
        src121 <= 16'hfb48;
        src122 <= 16'he8b0;
        src123 <= 16'h90ea;
        src124 <= 16'hdfda;
        src125 <= 16'h87d0;
        src126 <= 16'h7fbc;
        src127 <= 16'haacf;
        src128 <= 16'hf8ed;
        src129 <= 16'h8d43;
        src130 <= 16'h3f4f;
        src131 <= 16'h9dc;
        src132 <= 16'h1c02;
        src133 <= 16'h65a6;
        src134 <= 16'h1be7;
        src135 <= 16'hf17;
        src136 <= 16'h3153;
        src137 <= 16'hf95f;
        src138 <= 16'h621b;
        src139 <= 16'h8c40;
        src140 <= 16'h5206;
        src141 <= 16'h7d84;
        src142 <= 16'hce9;
        src143 <= 16'haa18;
        src144 <= 16'hc408;
        src145 <= 16'h6678;
        src146 <= 16'h3b5d;
        src147 <= 16'ha37a;
        src148 <= 16'h72dd;
        src149 <= 16'h8e6f;
        src150 <= 16'h2c97;
        src151 <= 16'hf155;
        src152 <= 16'hc08;
        src153 <= 16'hc9cb;
        src154 <= 16'he8cc;
        src155 <= 16'h8752;
        src156 <= 16'h10c0;
        src157 <= 16'hc16c;
        src158 <= 16'hcf8e;
        src159 <= 16'h5324;
        src160 <= 16'hc1ee;
        src161 <= 16'h52d6;
        src162 <= 16'hb6fd;
        src163 <= 16'hc7f6;
        src164 <= 16'hbc47;
        src165 <= 16'h9c3c;
        src166 <= 16'h440a;
        src167 <= 16'hc119;
        src168 <= 16'h33aa;
        src169 <= 16'h7180;
        src170 <= 16'h7e35;
        src171 <= 16'h5ff8;
        src172 <= 16'h7ce3;
        src173 <= 16'h8a92;
        src174 <= 16'h5841;
        src175 <= 16'h1569;
        src176 <= 16'h6e9f;
        src177 <= 16'h391;
        src178 <= 16'hd446;
        src179 <= 16'hf662;
        src180 <= 16'h3125;
        src181 <= 16'h9f2b;
        src182 <= 16'h5c86;
        src183 <= 16'hfcf5;
        src184 <= 16'hf4dc;
        exp <= 24'h5e315e;
        #1
        src0 <= 16'h3455;
        src1 <= 16'he91c;
        src2 <= 16'h254b;
        src3 <= 16'ha5af;
        src4 <= 16'ha7d1;
        src5 <= 16'h342;
        src6 <= 16'h7029;
        src7 <= 16'h17a2;
        src8 <= 16'h2670;
        src9 <= 16'h6f84;
        src10 <= 16'h97c9;
        src11 <= 16'h12de;
        src12 <= 16'h91d7;
        src13 <= 16'hbe00;
        src14 <= 16'h5814;
        src15 <= 16'h720b;
        src16 <= 16'h64c8;
        src17 <= 16'hf495;
        src18 <= 16'h2a1c;
        src19 <= 16'h976a;
        src20 <= 16'ha7c1;
        src21 <= 16'h8d8c;
        src22 <= 16'ha7a7;
        src23 <= 16'h7bde;
        src24 <= 16'h3222;
        src25 <= 16'h41e2;
        src26 <= 16'hc9b6;
        src27 <= 16'h4d19;
        src28 <= 16'h178;
        src29 <= 16'h8321;
        src30 <= 16'h47a0;
        src31 <= 16'h8d27;
        src32 <= 16'h2af8;
        src33 <= 16'h866f;
        src34 <= 16'h3140;
        src35 <= 16'hbd02;
        src36 <= 16'hb02e;
        src37 <= 16'h8646;
        src38 <= 16'h3be8;
        src39 <= 16'h4276;
        src40 <= 16'ha9fb;
        src41 <= 16'h3d0f;
        src42 <= 16'h2a85;
        src43 <= 16'h75f6;
        src44 <= 16'h1073;
        src45 <= 16'h2319;
        src46 <= 16'h1369;
        src47 <= 16'h3a41;
        src48 <= 16'h44e8;
        src49 <= 16'h124c;
        src50 <= 16'he0f3;
        src51 <= 16'hea92;
        src52 <= 16'hf289;
        src53 <= 16'h9372;
        src54 <= 16'h6064;
        src55 <= 16'h2f5d;
        src56 <= 16'h24f2;
        src57 <= 16'h66f7;
        src58 <= 16'h6752;
        src59 <= 16'h92ae;
        src60 <= 16'hf756;
        src61 <= 16'h8df3;
        src62 <= 16'h5281;
        src63 <= 16'h2886;
        src64 <= 16'h9f79;
        src65 <= 16'h2ed4;
        src66 <= 16'ha0b8;
        src67 <= 16'h78a8;
        src68 <= 16'hcafc;
        src69 <= 16'h6e05;
        src70 <= 16'h61e2;
        src71 <= 16'hc875;
        src72 <= 16'h5eb0;
        src73 <= 16'h5b7e;
        src74 <= 16'h733a;
        src75 <= 16'hf3ed;
        src76 <= 16'h6b6f;
        src77 <= 16'he1a0;
        src78 <= 16'h1629;
        src79 <= 16'h917d;
        src80 <= 16'hb985;
        src81 <= 16'h1d20;
        src82 <= 16'h9c89;
        src83 <= 16'h698b;
        src84 <= 16'h573d;
        src85 <= 16'hca25;
        src86 <= 16'ha8d9;
        src87 <= 16'h2134;
        src88 <= 16'hab9f;
        src89 <= 16'hc4f2;
        src90 <= 16'h6830;
        src91 <= 16'h9bf2;
        src92 <= 16'ha6c;
        src93 <= 16'h1483;
        src94 <= 16'h2995;
        src95 <= 16'h7f45;
        src96 <= 16'h1cde;
        src97 <= 16'h29e2;
        src98 <= 16'h163f;
        src99 <= 16'h996;
        src100 <= 16'ha0e4;
        src101 <= 16'h25e0;
        src102 <= 16'h3cc6;
        src103 <= 16'h92c8;
        src104 <= 16'hf531;
        src105 <= 16'h573d;
        src106 <= 16'h6532;
        src107 <= 16'h133b;
        src108 <= 16'had04;
        src109 <= 16'h26c4;
        src110 <= 16'hff28;
        src111 <= 16'h108f;
        src112 <= 16'hd3c0;
        src113 <= 16'hf091;
        src114 <= 16'h4e48;
        src115 <= 16'h5dbc;
        src116 <= 16'h86d5;
        src117 <= 16'h878f;
        src118 <= 16'he1ed;
        src119 <= 16'h805;
        src120 <= 16'h7500;
        src121 <= 16'h82c1;
        src122 <= 16'h5d80;
        src123 <= 16'h2df9;
        src124 <= 16'h2ce3;
        src125 <= 16'h2aea;
        src126 <= 16'hc7bc;
        src127 <= 16'hcaef;
        src128 <= 16'h1778;
        src129 <= 16'h3e54;
        src130 <= 16'heb68;
        src131 <= 16'h9b1f;
        src132 <= 16'hc4ea;
        src133 <= 16'hadfa;
        src134 <= 16'hd6dc;
        src135 <= 16'hd9fb;
        src136 <= 16'haa24;
        src137 <= 16'hdc60;
        src138 <= 16'h3b30;
        src139 <= 16'h8b45;
        src140 <= 16'h9934;
        src141 <= 16'h9598;
        src142 <= 16'hc848;
        src143 <= 16'hfe37;
        src144 <= 16'hb775;
        src145 <= 16'h81c8;
        src146 <= 16'h3abb;
        src147 <= 16'he293;
        src148 <= 16'h80b5;
        src149 <= 16'he7db;
        src150 <= 16'h1b93;
        src151 <= 16'h160b;
        src152 <= 16'hb515;
        src153 <= 16'hee5c;
        src154 <= 16'h725f;
        src155 <= 16'haa7d;
        src156 <= 16'h7cc3;
        src157 <= 16'ha789;
        src158 <= 16'h73ac;
        src159 <= 16'hd40a;
        src160 <= 16'haa0f;
        src161 <= 16'hf7d;
        src162 <= 16'hd3c1;
        src163 <= 16'h18f9;
        src164 <= 16'hc88a;
        src165 <= 16'h4150;
        src166 <= 16'haf78;
        src167 <= 16'h4169;
        src168 <= 16'h64b1;
        src169 <= 16'h59b5;
        src170 <= 16'hb0c4;
        src171 <= 16'hed3f;
        src172 <= 16'hfa77;
        src173 <= 16'hd987;
        src174 <= 16'h5e6c;
        src175 <= 16'hdb73;
        src176 <= 16'h194b;
        src177 <= 16'h17bf;
        src178 <= 16'h3c03;
        src179 <= 16'h6758;
        src180 <= 16'hee34;
        src181 <= 16'h6c83;
        src182 <= 16'h6327;
        src183 <= 16'hc537;
        src184 <= 16'hadf1;
        exp <= 24'h583b03;
        #1
        src0 <= 16'h3d23;
        src1 <= 16'he306;
        src2 <= 16'hff8c;
        src3 <= 16'h1509;
        src4 <= 16'h3e97;
        src5 <= 16'ha2e8;
        src6 <= 16'hbad3;
        src7 <= 16'h21b4;
        src8 <= 16'hadcc;
        src9 <= 16'h937;
        src10 <= 16'hcc1b;
        src11 <= 16'ha3a;
        src12 <= 16'h6715;
        src13 <= 16'ha7c8;
        src14 <= 16'h103e;
        src15 <= 16'h8af9;
        src16 <= 16'hfbe8;
        src17 <= 16'hb855;
        src18 <= 16'h4e8b;
        src19 <= 16'hb1aa;
        src20 <= 16'hb5f6;
        src21 <= 16'he7db;
        src22 <= 16'h5227;
        src23 <= 16'h12bf;
        src24 <= 16'h747a;
        src25 <= 16'h5131;
        src26 <= 16'h6296;
        src27 <= 16'h586c;
        src28 <= 16'h2b6d;
        src29 <= 16'h747f;
        src30 <= 16'hed09;
        src31 <= 16'h360;
        src32 <= 16'hbbce;
        src33 <= 16'h5e5;
        src34 <= 16'h1427;
        src35 <= 16'h1538;
        src36 <= 16'h52aa;
        src37 <= 16'h5c92;
        src38 <= 16'h2cb9;
        src39 <= 16'he746;
        src40 <= 16'hc4f4;
        src41 <= 16'h81a1;
        src42 <= 16'h1b40;
        src43 <= 16'h386f;
        src44 <= 16'hfec;
        src45 <= 16'hacfd;
        src46 <= 16'h7112;
        src47 <= 16'hff21;
        src48 <= 16'h8691;
        src49 <= 16'hb873;
        src50 <= 16'h3963;
        src51 <= 16'ha6ce;
        src52 <= 16'h3325;
        src53 <= 16'h5821;
        src54 <= 16'hf8b6;
        src55 <= 16'h257;
        src56 <= 16'h4863;
        src57 <= 16'h171f;
        src58 <= 16'hfcdd;
        src59 <= 16'h6ae2;
        src60 <= 16'h3cad;
        src61 <= 16'h7f92;
        src62 <= 16'hb510;
        src63 <= 16'h86c1;
        src64 <= 16'h60eb;
        src65 <= 16'ha6e1;
        src66 <= 16'hb9cd;
        src67 <= 16'hec64;
        src68 <= 16'hd9e0;
        src69 <= 16'h8c71;
        src70 <= 16'h88d1;
        src71 <= 16'h7022;
        src72 <= 16'h1ec2;
        src73 <= 16'h72c4;
        src74 <= 16'h8b10;
        src75 <= 16'hda70;
        src76 <= 16'hb427;
        src77 <= 16'h5ac4;
        src78 <= 16'h4aba;
        src79 <= 16'hab2c;
        src80 <= 16'hd37d;
        src81 <= 16'he955;
        src82 <= 16'h893a;
        src83 <= 16'h167f;
        src84 <= 16'hce7;
        src85 <= 16'h8d7d;
        src86 <= 16'he9fe;
        src87 <= 16'hb811;
        src88 <= 16'h6690;
        src89 <= 16'h55e9;
        src90 <= 16'h2530;
        src91 <= 16'h6391;
        src92 <= 16'h7adb;
        src93 <= 16'h76ec;
        src94 <= 16'h5513;
        src95 <= 16'hf3fb;
        src96 <= 16'hfa1;
        src97 <= 16'h815a;
        src98 <= 16'hb28d;
        src99 <= 16'hdff7;
        src100 <= 16'h9549;
        src101 <= 16'hcf0a;
        src102 <= 16'hc549;
        src103 <= 16'h9aa1;
        src104 <= 16'hdfcd;
        src105 <= 16'h54ab;
        src106 <= 16'hb1e6;
        src107 <= 16'hdb8e;
        src108 <= 16'h1c3b;
        src109 <= 16'h1f03;
        src110 <= 16'h78e2;
        src111 <= 16'hec2e;
        src112 <= 16'h11c0;
        src113 <= 16'h1a5a;
        src114 <= 16'he179;
        src115 <= 16'hbeb9;
        src116 <= 16'ha97a;
        src117 <= 16'he234;
        src118 <= 16'hd617;
        src119 <= 16'h51a9;
        src120 <= 16'hcece;
        src121 <= 16'h2f89;
        src122 <= 16'ha123;
        src123 <= 16'h78a4;
        src124 <= 16'h10f7;
        src125 <= 16'h35ea;
        src126 <= 16'haca4;
        src127 <= 16'h7b05;
        src128 <= 16'h3291;
        src129 <= 16'h77ef;
        src130 <= 16'h16d2;
        src131 <= 16'h1ce3;
        src132 <= 16'hd826;
        src133 <= 16'hf5a0;
        src134 <= 16'h1275;
        src135 <= 16'h724a;
        src136 <= 16'hd7df;
        src137 <= 16'h3347;
        src138 <= 16'hf0fd;
        src139 <= 16'h2909;
        src140 <= 16'ha27f;
        src141 <= 16'h2b3a;
        src142 <= 16'h6dfd;
        src143 <= 16'hd2df;
        src144 <= 16'hadfb;
        src145 <= 16'h6a0f;
        src146 <= 16'h82bb;
        src147 <= 16'hba81;
        src148 <= 16'hd070;
        src149 <= 16'hc7a;
        src150 <= 16'h6b5b;
        src151 <= 16'hbadc;
        src152 <= 16'h567d;
        src153 <= 16'h289e;
        src154 <= 16'heb85;
        src155 <= 16'h5333;
        src156 <= 16'h3ea9;
        src157 <= 16'he573;
        src158 <= 16'h7068;
        src159 <= 16'h1f7c;
        src160 <= 16'h3b96;
        src161 <= 16'h2756;
        src162 <= 16'h9079;
        src163 <= 16'h7f7d;
        src164 <= 16'h9353;
        src165 <= 16'h97e4;
        src166 <= 16'hfe2a;
        src167 <= 16'h2bad;
        src168 <= 16'haf33;
        src169 <= 16'hd728;
        src170 <= 16'h9c1d;
        src171 <= 16'hf799;
        src172 <= 16'hbc34;
        src173 <= 16'h5f3b;
        src174 <= 16'h78dc;
        src175 <= 16'hd98d;
        src176 <= 16'hf6ad;
        src177 <= 16'h1120;
        src178 <= 16'h458b;
        src179 <= 16'h65a7;
        src180 <= 16'hfe21;
        src181 <= 16'h7106;
        src182 <= 16'hc014;
        src183 <= 16'hc99c;
        src184 <= 16'ha059;
        exp <= 24'h5d0a1b;
        #1
        src0 <= 16'h8884;
        src1 <= 16'hb98a;
        src2 <= 16'h6e9b;
        src3 <= 16'hd12e;
        src4 <= 16'h56be;
        src5 <= 16'hc4b4;
        src6 <= 16'he382;
        src7 <= 16'h84b8;
        src8 <= 16'h8b37;
        src9 <= 16'he5fd;
        src10 <= 16'h2e23;
        src11 <= 16'h3ce1;
        src12 <= 16'hb624;
        src13 <= 16'hd045;
        src14 <= 16'haa3;
        src15 <= 16'hdc7d;
        src16 <= 16'hc0aa;
        src17 <= 16'hf50e;
        src18 <= 16'h84d6;
        src19 <= 16'hea7a;
        src20 <= 16'h3ffe;
        src21 <= 16'ha788;
        src22 <= 16'h49d7;
        src23 <= 16'hfacd;
        src24 <= 16'haa89;
        src25 <= 16'hbd2b;
        src26 <= 16'h5090;
        src27 <= 16'h108a;
        src28 <= 16'hc1b1;
        src29 <= 16'h9f23;
        src30 <= 16'h2f99;
        src31 <= 16'h9871;
        src32 <= 16'h1337;
        src33 <= 16'hc8f2;
        src34 <= 16'he0b7;
        src35 <= 16'h40eb;
        src36 <= 16'h4d15;
        src37 <= 16'hf4e9;
        src38 <= 16'h109;
        src39 <= 16'h7b2e;
        src40 <= 16'h3226;
        src41 <= 16'ha6ae;
        src42 <= 16'he5e1;
        src43 <= 16'hef22;
        src44 <= 16'ha746;
        src45 <= 16'h8c82;
        src46 <= 16'h6e55;
        src47 <= 16'h43ab;
        src48 <= 16'hd4f9;
        src49 <= 16'ha882;
        src50 <= 16'he25f;
        src51 <= 16'hc99c;
        src52 <= 16'h8;
        src53 <= 16'h742c;
        src54 <= 16'he150;
        src55 <= 16'h20d;
        src56 <= 16'h4627;
        src57 <= 16'h749d;
        src58 <= 16'haaca;
        src59 <= 16'hce1f;
        src60 <= 16'hfcf4;
        src61 <= 16'h4546;
        src62 <= 16'h152e;
        src63 <= 16'h205d;
        src64 <= 16'h5bd7;
        src65 <= 16'h2f57;
        src66 <= 16'hc1e9;
        src67 <= 16'h20dd;
        src68 <= 16'h4bb6;
        src69 <= 16'ha191;
        src70 <= 16'hae2d;
        src71 <= 16'hed40;
        src72 <= 16'hc322;
        src73 <= 16'h8929;
        src74 <= 16'h541f;
        src75 <= 16'h44be;
        src76 <= 16'hcc4d;
        src77 <= 16'h3b32;
        src78 <= 16'ha8f1;
        src79 <= 16'h7719;
        src80 <= 16'hba1b;
        src81 <= 16'h6d23;
        src82 <= 16'ha4cb;
        src83 <= 16'h5e74;
        src84 <= 16'hc699;
        src85 <= 16'h42a4;
        src86 <= 16'h2126;
        src87 <= 16'he685;
        src88 <= 16'h8af8;
        src89 <= 16'h3ecf;
        src90 <= 16'hdb9b;
        src91 <= 16'h54ac;
        src92 <= 16'h4b66;
        src93 <= 16'h6800;
        src94 <= 16'h66cb;
        src95 <= 16'hf8ed;
        src96 <= 16'h31d5;
        src97 <= 16'hb915;
        src98 <= 16'h9d6;
        src99 <= 16'h241f;
        src100 <= 16'h6c8e;
        src101 <= 16'hd446;
        src102 <= 16'h496e;
        src103 <= 16'h347d;
        src104 <= 16'h811c;
        src105 <= 16'h63d;
        src106 <= 16'he09b;
        src107 <= 16'h49f9;
        src108 <= 16'hb438;
        src109 <= 16'h8b11;
        src110 <= 16'hb61e;
        src111 <= 16'he3f;
        src112 <= 16'h98ca;
        src113 <= 16'h1437;
        src114 <= 16'h58fc;
        src115 <= 16'h4c56;
        src116 <= 16'h738f;
        src117 <= 16'h8b59;
        src118 <= 16'hc17b;
        src119 <= 16'he64b;
        src120 <= 16'hc2f;
        src121 <= 16'hec5c;
        src122 <= 16'hd77b;
        src123 <= 16'h176f;
        src124 <= 16'h4f0;
        src125 <= 16'h9f16;
        src126 <= 16'h9e4c;
        src127 <= 16'hcdfc;
        src128 <= 16'h2f94;
        src129 <= 16'h5d6d;
        src130 <= 16'h47aa;
        src131 <= 16'he1a5;
        src132 <= 16'hbf30;
        src133 <= 16'h57ff;
        src134 <= 16'hca34;
        src135 <= 16'h4f53;
        src136 <= 16'h3a27;
        src137 <= 16'h1167;
        src138 <= 16'h397f;
        src139 <= 16'h62fc;
        src140 <= 16'h96c4;
        src141 <= 16'hb391;
        src142 <= 16'h7026;
        src143 <= 16'h5d70;
        src144 <= 16'h4dec;
        src145 <= 16'hb731;
        src146 <= 16'hc486;
        src147 <= 16'h35b2;
        src148 <= 16'h4b6f;
        src149 <= 16'h8c6f;
        src150 <= 16'hba05;
        src151 <= 16'h887c;
        src152 <= 16'hb60f;
        src153 <= 16'h1d57;
        src154 <= 16'h9aa2;
        src155 <= 16'h1478;
        src156 <= 16'he4fa;
        src157 <= 16'h5eef;
        src158 <= 16'h2abd;
        src159 <= 16'hb78d;
        src160 <= 16'h646e;
        src161 <= 16'hcdb7;
        src162 <= 16'h3200;
        src163 <= 16'h620d;
        src164 <= 16'h9d7d;
        src165 <= 16'h9fd2;
        src166 <= 16'hf6d0;
        src167 <= 16'hbf2a;
        src168 <= 16'h9ae9;
        src169 <= 16'h5c56;
        src170 <= 16'he096;
        src171 <= 16'hb1e0;
        src172 <= 16'h6127;
        src173 <= 16'hccb5;
        src174 <= 16'he21;
        src175 <= 16'hc0f6;
        src176 <= 16'hd484;
        src177 <= 16'hf1ff;
        src178 <= 16'hbcb0;
        src179 <= 16'ha835;
        src180 <= 16'hfd81;
        src181 <= 16'h2aa9;
        src182 <= 16'hd1d0;
        src183 <= 16'hd9f6;
        src184 <= 16'h7022;
        exp <= 24'h603117;
        #1
        src0 <= 16'hbbbe;
        src1 <= 16'he08d;
        src2 <= 16'h579;
        src3 <= 16'h88e;
        src4 <= 16'h4e15;
        src5 <= 16'h4d35;
        src6 <= 16'h35d2;
        src7 <= 16'h8574;
        src8 <= 16'h1fd7;
        src9 <= 16'hea18;
        src10 <= 16'ha8b5;
        src11 <= 16'hfce8;
        src12 <= 16'hf5e4;
        src13 <= 16'hf120;
        src14 <= 16'h24fe;
        src15 <= 16'hf425;
        src16 <= 16'h2aea;
        src17 <= 16'hb0dc;
        src18 <= 16'hca9e;
        src19 <= 16'h543a;
        src20 <= 16'he7f;
        src21 <= 16'h80bd;
        src22 <= 16'h980c;
        src23 <= 16'h79ce;
        src24 <= 16'h6e99;
        src25 <= 16'hbe7c;
        src26 <= 16'hcc81;
        src27 <= 16'h1a1a;
        src28 <= 16'h7f70;
        src29 <= 16'haffb;
        src30 <= 16'h7e35;
        src31 <= 16'hfafe;
        src32 <= 16'h30c0;
        src33 <= 16'h8e10;
        src34 <= 16'h674b;
        src35 <= 16'hcea1;
        src36 <= 16'h8619;
        src37 <= 16'hc1d3;
        src38 <= 16'h7680;
        src39 <= 16'hbbdd;
        src40 <= 16'hf4ac;
        src41 <= 16'h68e0;
        src42 <= 16'h64d;
        src43 <= 16'h62a8;
        src44 <= 16'h9145;
        src45 <= 16'h4edb;
        src46 <= 16'hfe3c;
        src47 <= 16'h670f;
        src48 <= 16'hfcc;
        src49 <= 16'hfd2f;
        src50 <= 16'he2de;
        src51 <= 16'h3f38;
        src52 <= 16'h893b;
        src53 <= 16'h2271;
        src54 <= 16'h59ba;
        src55 <= 16'h57dd;
        src56 <= 16'hd9a;
        src57 <= 16'h32f8;
        src58 <= 16'h83af;
        src59 <= 16'hf282;
        src60 <= 16'hbf88;
        src61 <= 16'h8352;
        src62 <= 16'h5e4b;
        src63 <= 16'hec12;
        src64 <= 16'hecbf;
        src65 <= 16'hafd0;
        src66 <= 16'h50ab;
        src67 <= 16'hbb7d;
        src68 <= 16'he272;
        src69 <= 16'h5f35;
        src70 <= 16'h9a27;
        src71 <= 16'had62;
        src72 <= 16'h1e27;
        src73 <= 16'ha5e9;
        src74 <= 16'h75b7;
        src75 <= 16'hdc92;
        src76 <= 16'h7760;
        src77 <= 16'h4014;
        src78 <= 16'h7b2b;
        src79 <= 16'hddbe;
        src80 <= 16'h122f;
        src81 <= 16'h2dc9;
        src82 <= 16'h195c;
        src83 <= 16'habc2;
        src84 <= 16'h441c;
        src85 <= 16'h898b;
        src86 <= 16'h90d3;
        src87 <= 16'h27a0;
        src88 <= 16'h5ba6;
        src89 <= 16'hcd1f;
        src90 <= 16'h7518;
        src91 <= 16'he0f3;
        src92 <= 16'he72e;
        src93 <= 16'h4923;
        src94 <= 16'he1d3;
        src95 <= 16'h5725;
        src96 <= 16'hb19e;
        src97 <= 16'h5778;
        src98 <= 16'h7e5f;
        src99 <= 16'h3917;
        src100 <= 16'hfc04;
        src101 <= 16'h1216;
        src102 <= 16'h5dfb;
        src103 <= 16'hcdd;
        src104 <= 16'hec16;
        src105 <= 16'hf08d;
        src106 <= 16'hcf85;
        src107 <= 16'h8c6a;
        src108 <= 16'ha716;
        src109 <= 16'hfddc;
        src110 <= 16'h1d25;
        src111 <= 16'ha4cd;
        src112 <= 16'hefb9;
        src113 <= 16'hb7da;
        src114 <= 16'ha4fc;
        src115 <= 16'h42c1;
        src116 <= 16'he3d8;
        src117 <= 16'h878d;
        src118 <= 16'h9707;
        src119 <= 16'h4bca;
        src120 <= 16'h9d53;
        src121 <= 16'h1678;
        src122 <= 16'h461e;
        src123 <= 16'h14fc;
        src124 <= 16'h6a27;
        src125 <= 16'hcfea;
        src126 <= 16'h4af9;
        src127 <= 16'hdfb3;
        src128 <= 16'h3e10;
        src129 <= 16'hd6e7;
        src130 <= 16'hed11;
        src131 <= 16'hcf6e;
        src132 <= 16'h7734;
        src133 <= 16'h532e;
        src134 <= 16'hbc0d;
        src135 <= 16'hfafa;
        src136 <= 16'hc8fc;
        src137 <= 16'h250a;
        src138 <= 16'hdff7;
        src139 <= 16'hc5d5;
        src140 <= 16'h90fd;
        src141 <= 16'h7e7a;
        src142 <= 16'h2ddf;
        src143 <= 16'h790a;
        src144 <= 16'hcc55;
        src145 <= 16'hc4e0;
        src146 <= 16'h60b0;
        src147 <= 16'hcbd7;
        src148 <= 16'h6d3;
        src149 <= 16'h617a;
        src150 <= 16'he162;
        src151 <= 16'hd8c8;
        src152 <= 16'h9dc3;
        src153 <= 16'h7b53;
        src154 <= 16'h8ba9;
        src155 <= 16'h2b7e;
        src156 <= 16'h4212;
        src157 <= 16'h15e9;
        src158 <= 16'h374b;
        src159 <= 16'hf64d;
        src160 <= 16'h380f;
        src161 <= 16'hcde3;
        src162 <= 16'hbecd;
        src163 <= 16'hba92;
        src164 <= 16'h7f70;
        src165 <= 16'h43c5;
        src166 <= 16'h3863;
        src167 <= 16'h6de1;
        src168 <= 16'he0d;
        src169 <= 16'heece;
        src170 <= 16'h1002;
        src171 <= 16'h6441;
        src172 <= 16'hf02a;
        src173 <= 16'h7623;
        src174 <= 16'h7e6d;
        src175 <= 16'h22c1;
        src176 <= 16'h9b17;
        src177 <= 16'h2cb7;
        src178 <= 16'h88d9;
        src179 <= 16'hdf22;
        src180 <= 16'h48e6;
        src181 <= 16'h57a;
        src182 <= 16'h5107;
        src183 <= 16'hd3f;
        src184 <= 16'h1d50;
        exp <= 24'h5f780e;
        #1
        src0 <= 16'h4314;
        src1 <= 16'h78fc;
        src2 <= 16'h289e;
        src3 <= 16'h6422;
        src4 <= 16'h95d;
        src5 <= 16'h2535;
        src6 <= 16'h66f4;
        src7 <= 16'hbf36;
        src8 <= 16'h585b;
        src9 <= 16'ha09c;
        src10 <= 16'hc149;
        src11 <= 16'hfbcf;
        src12 <= 16'h200b;
        src13 <= 16'h87c6;
        src14 <= 16'h805a;
        src15 <= 16'h329;
        src16 <= 16'h327f;
        src17 <= 16'h2ac9;
        src18 <= 16'h7d20;
        src19 <= 16'hce49;
        src20 <= 16'h608e;
        src21 <= 16'h374d;
        src22 <= 16'h7585;
        src23 <= 16'h49ef;
        src24 <= 16'h8b4f;
        src25 <= 16'hfd96;
        src26 <= 16'he802;
        src27 <= 16'h3f40;
        src28 <= 16'h86b2;
        src29 <= 16'h506c;
        src30 <= 16'h7959;
        src31 <= 16'h72c4;
        src32 <= 16'hf47;
        src33 <= 16'ha62c;
        src34 <= 16'h974c;
        src35 <= 16'hdbff;
        src36 <= 16'h582;
        src37 <= 16'h4875;
        src38 <= 16'h877c;
        src39 <= 16'h4887;
        src40 <= 16'h3f3;
        src41 <= 16'h2ec1;
        src42 <= 16'hafc1;
        src43 <= 16'h88df;
        src44 <= 16'h9b87;
        src45 <= 16'h8e29;
        src46 <= 16'h430a;
        src47 <= 16'h9715;
        src48 <= 16'h6afc;
        src49 <= 16'ha629;
        src50 <= 16'h8b10;
        src51 <= 16'had84;
        src52 <= 16'h2e7;
        src53 <= 16'h7873;
        src54 <= 16'h7897;
        src55 <= 16'h7d90;
        src56 <= 16'h4a9b;
        src57 <= 16'h66e1;
        src58 <= 16'h711;
        src59 <= 16'h9450;
        src60 <= 16'h5617;
        src61 <= 16'hcb51;
        src62 <= 16'he4e6;
        src63 <= 16'hd7d1;
        src64 <= 16'hada8;
        src65 <= 16'h2c1f;
        src66 <= 16'he6e0;
        src67 <= 16'hc450;
        src68 <= 16'h4cef;
        src69 <= 16'h522d;
        src70 <= 16'h62f;
        src71 <= 16'hdcbc;
        src72 <= 16'hf81c;
        src73 <= 16'h8c6a;
        src74 <= 16'h25fc;
        src75 <= 16'h30c;
        src76 <= 16'hbd72;
        src77 <= 16'h85f9;
        src78 <= 16'h25fe;
        src79 <= 16'h8356;
        src80 <= 16'h6139;
        src81 <= 16'h1033;
        src82 <= 16'h253b;
        src83 <= 16'h1927;
        src84 <= 16'he636;
        src85 <= 16'h94cf;
        src86 <= 16'h6fe7;
        src87 <= 16'hfdec;
        src88 <= 16'hf6cd;
        src89 <= 16'ha108;
        src90 <= 16'h75ab;
        src91 <= 16'h3a4e;
        src92 <= 16'hd02e;
        src93 <= 16'he550;
        src94 <= 16'hd3bf;
        src95 <= 16'h2f53;
        src96 <= 16'h6fb0;
        src97 <= 16'ha6ca;
        src98 <= 16'h837d;
        src99 <= 16'h34c1;
        src100 <= 16'hd675;
        src101 <= 16'h6d6a;
        src102 <= 16'h6935;
        src103 <= 16'h663d;
        src104 <= 16'he4c9;
        src105 <= 16'heff2;
        src106 <= 16'hffaf;
        src107 <= 16'h51ac;
        src108 <= 16'hb727;
        src109 <= 16'hca02;
        src110 <= 16'h4cbf;
        src111 <= 16'h54b5;
        src112 <= 16'h328e;
        src113 <= 16'h53a8;
        src114 <= 16'h858;
        src115 <= 16'h3384;
        src116 <= 16'hd140;
        src117 <= 16'hfc7d;
        src118 <= 16'h3938;
        src119 <= 16'h9f4;
        src120 <= 16'h7bcc;
        src121 <= 16'hc926;
        src122 <= 16'h53c9;
        src123 <= 16'hdc2e;
        src124 <= 16'hb799;
        src125 <= 16'hf11a;
        src126 <= 16'hb96a;
        src127 <= 16'h46a4;
        src128 <= 16'h5bff;
        src129 <= 16'h1812;
        src130 <= 16'h9169;
        src131 <= 16'hf988;
        src132 <= 16'h63c1;
        src133 <= 16'he4b4;
        src134 <= 16'h921c;
        src135 <= 16'h545;
        src136 <= 16'h4d29;
        src137 <= 16'h1b73;
        src138 <= 16'h56f1;
        src139 <= 16'hdd5f;
        src140 <= 16'h3b33;
        src141 <= 16'h9512;
        src142 <= 16'hbf18;
        src143 <= 16'h4d17;
        src144 <= 16'h33c;
        src145 <= 16'h6e5c;
        src146 <= 16'he5d9;
        src147 <= 16'h4af7;
        src148 <= 16'h5532;
        src149 <= 16'hf42d;
        src150 <= 16'hc230;
        src151 <= 16'ha4ea;
        src152 <= 16'hc32d;
        src153 <= 16'h8566;
        src154 <= 16'h1cc4;
        src155 <= 16'h7fa1;
        src156 <= 16'hee06;
        src157 <= 16'h404a;
        src158 <= 16'hf2c0;
        src159 <= 16'h64d5;
        src160 <= 16'h9080;
        src161 <= 16'h4097;
        src162 <= 16'hb69c;
        src163 <= 16'hae58;
        src164 <= 16'hd402;
        src165 <= 16'hacf1;
        src166 <= 16'hfbf2;
        src167 <= 16'hc160;
        src168 <= 16'h5741;
        src169 <= 16'h39fd;
        src170 <= 16'hb36d;
        src171 <= 16'hc912;
        src172 <= 16'h7843;
        src173 <= 16'h412a;
        src174 <= 16'h36b4;
        src175 <= 16'h668b;
        src176 <= 16'h828d;
        src177 <= 16'h8e07;
        src178 <= 16'h1018;
        src179 <= 16'h25ef;
        src180 <= 16'hed32;
        src181 <= 16'hefba;
        src182 <= 16'h3bb3;
        src183 <= 16'h6f9;
        src184 <= 16'h65ff;
        exp <= 24'h5a9ef3;
        #1
        src0 <= 16'hf45b;
        src1 <= 16'h56ca;
        src2 <= 16'h1d89;
        src3 <= 16'he38b;
        src4 <= 16'hae10;
        src5 <= 16'hebe6;
        src6 <= 16'hd06d;
        src7 <= 16'h18cf;
        src8 <= 16'h405b;
        src9 <= 16'h43eb;
        src10 <= 16'h5e5c;
        src11 <= 16'hc714;
        src12 <= 16'he441;
        src13 <= 16'haa98;
        src14 <= 16'h8b29;
        src15 <= 16'h89e0;
        src16 <= 16'h10ef;
        src17 <= 16'h56fb;
        src18 <= 16'hacb0;
        src19 <= 16'hceb1;
        src20 <= 16'he5fb;
        src21 <= 16'hece7;
        src22 <= 16'ha0da;
        src23 <= 16'hf7a4;
        src24 <= 16'h98ca;
        src25 <= 16'haf0d;
        src26 <= 16'haa5;
        src27 <= 16'h93a5;
        src28 <= 16'h6a1b;
        src29 <= 16'h8eb1;
        src30 <= 16'hd69b;
        src31 <= 16'h2718;
        src32 <= 16'h666c;
        src33 <= 16'h9457;
        src34 <= 16'hdd07;
        src35 <= 16'h2d84;
        src36 <= 16'h924d;
        src37 <= 16'h1b26;
        src38 <= 16'h57ce;
        src39 <= 16'he220;
        src40 <= 16'hc3fc;
        src41 <= 16'h82dd;
        src42 <= 16'hf38e;
        src43 <= 16'hf3c3;
        src44 <= 16'h83b8;
        src45 <= 16'hc112;
        src46 <= 16'h2513;
        src47 <= 16'h59a4;
        src48 <= 16'h9509;
        src49 <= 16'hd1f3;
        src50 <= 16'h1d03;
        src51 <= 16'h9d7f;
        src52 <= 16'h83f8;
        src53 <= 16'he9f8;
        src54 <= 16'he7f7;
        src55 <= 16'h2f3a;
        src56 <= 16'h542b;
        src57 <= 16'h4834;
        src58 <= 16'ha27c;
        src59 <= 16'h6b8e;
        src60 <= 16'h81d3;
        src61 <= 16'hdf00;
        src62 <= 16'hf1c0;
        src63 <= 16'h5ca9;
        src64 <= 16'h8013;
        src65 <= 16'h31c2;
        src66 <= 16'h9668;
        src67 <= 16'hffd8;
        src68 <= 16'h8cc8;
        src69 <= 16'hcf6e;
        src70 <= 16'hda8f;
        src71 <= 16'heff3;
        src72 <= 16'he213;
        src73 <= 16'he725;
        src74 <= 16'hb7f5;
        src75 <= 16'h247f;
        src76 <= 16'haaac;
        src77 <= 16'he061;
        src78 <= 16'h52fc;
        src79 <= 16'h8889;
        src80 <= 16'h97e3;
        src81 <= 16'h5957;
        src82 <= 16'h8e78;
        src83 <= 16'h715d;
        src84 <= 16'h50a7;
        src85 <= 16'h11da;
        src86 <= 16'h9afc;
        src87 <= 16'h2461;
        src88 <= 16'h1e31;
        src89 <= 16'h238d;
        src90 <= 16'h90c2;
        src91 <= 16'h4092;
        src92 <= 16'h543e;
        src93 <= 16'h3475;
        src94 <= 16'h7fef;
        src95 <= 16'h3212;
        src96 <= 16'hf702;
        src97 <= 16'h6c31;
        src98 <= 16'h231e;
        src99 <= 16'ha26a;
        src100 <= 16'h585b;
        src101 <= 16'h1215;
        src102 <= 16'hb70;
        src103 <= 16'h57e0;
        src104 <= 16'hecc5;
        src105 <= 16'h1dfa;
        src106 <= 16'hb44d;
        src107 <= 16'h8768;
        src108 <= 16'h15c7;
        src109 <= 16'hc671;
        src110 <= 16'hc4b8;
        src111 <= 16'hb943;
        src112 <= 16'h3542;
        src113 <= 16'h4bfa;
        src114 <= 16'h81b5;
        src115 <= 16'h86a0;
        src116 <= 16'hfc7c;
        src117 <= 16'hf8b9;
        src118 <= 16'h5921;
        src119 <= 16'h34de;
        src120 <= 16'h79a6;
        src121 <= 16'he614;
        src122 <= 16'h587c;
        src123 <= 16'hbd16;
        src124 <= 16'ha71f;
        src125 <= 16'h51f0;
        src126 <= 16'h74b;
        src127 <= 16'hed3b;
        src128 <= 16'he640;
        src129 <= 16'h9a6;
        src130 <= 16'h5689;
        src131 <= 16'h977a;
        src132 <= 16'h5d47;
        src133 <= 16'h6e1e;
        src134 <= 16'hfce7;
        src135 <= 16'h445b;
        src136 <= 16'h72d1;
        src137 <= 16'h92ae;
        src138 <= 16'h7499;
        src139 <= 16'h3203;
        src140 <= 16'h9742;
        src141 <= 16'he31a;
        src142 <= 16'h548e;
        src143 <= 16'h3565;
        src144 <= 16'hc4bf;
        src145 <= 16'h36ff;
        src146 <= 16'hb17;
        src147 <= 16'hca8e;
        src148 <= 16'h4d2b;
        src149 <= 16'h4088;
        src150 <= 16'hd81f;
        src151 <= 16'h30e0;
        src152 <= 16'hf797;
        src153 <= 16'h3e95;
        src154 <= 16'hbe32;
        src155 <= 16'h522e;
        src156 <= 16'h6642;
        src157 <= 16'he7fe;
        src158 <= 16'h3cc2;
        src159 <= 16'h6a35;
        src160 <= 16'hb97f;
        src161 <= 16'h2e98;
        src162 <= 16'h8202;
        src163 <= 16'hc734;
        src164 <= 16'hc791;
        src165 <= 16'he592;
        src166 <= 16'h44f9;
        src167 <= 16'h8f04;
        src168 <= 16'hdeaf;
        src169 <= 16'h8550;
        src170 <= 16'ha102;
        src171 <= 16'h1f40;
        src172 <= 16'h39a6;
        src173 <= 16'h5677;
        src174 <= 16'ha6b6;
        src175 <= 16'ha881;
        src176 <= 16'hb1fa;
        src177 <= 16'hf1d6;
        src178 <= 16'heb7;
        src179 <= 16'hfdda;
        src180 <= 16'ha365;
        src181 <= 16'hedcd;
        src182 <= 16'hd9a7;
        src183 <= 16'he292;
        src184 <= 16'h7b6d;
        exp <= 24'h62777f;
        #1
        src0 <= 16'ha770;
        src1 <= 16'h6091;
        src2 <= 16'h301b;
        src3 <= 16'hcd2b;
        src4 <= 16'h11b3;
        src5 <= 16'hbee9;
        src6 <= 16'h8896;
        src7 <= 16'hbb82;
        src8 <= 16'h7df7;
        src9 <= 16'h8c71;
        src10 <= 16'hd4ab;
        src11 <= 16'hd557;
        src12 <= 16'hab24;
        src13 <= 16'h9ce4;
        src14 <= 16'h917;
        src15 <= 16'h3e63;
        src16 <= 16'h7cd5;
        src17 <= 16'h93e3;
        src18 <= 16'h1858;
        src19 <= 16'hcf2a;
        src20 <= 16'h519c;
        src21 <= 16'h4223;
        src22 <= 16'he77e;
        src23 <= 16'h3c21;
        src24 <= 16'h3e0c;
        src25 <= 16'hcbc7;
        src26 <= 16'h44a5;
        src27 <= 16'hde7a;
        src28 <= 16'he592;
        src29 <= 16'h7493;
        src30 <= 16'h56ad;
        src31 <= 16'h5702;
        src32 <= 16'h84a3;
        src33 <= 16'haf27;
        src34 <= 16'h5d89;
        src35 <= 16'hf0d0;
        src36 <= 16'he18a;
        src37 <= 16'ha29;
        src38 <= 16'h94f3;
        src39 <= 16'h86f4;
        src40 <= 16'hcda2;
        src41 <= 16'h798f;
        src42 <= 16'h5365;
        src43 <= 16'h5c29;
        src44 <= 16'h4bbb;
        src45 <= 16'hc6db;
        src46 <= 16'h465b;
        src47 <= 16'hdfa9;
        src48 <= 16'hbae6;
        src49 <= 16'hd368;
        src50 <= 16'h72d8;
        src51 <= 16'h6a8;
        src52 <= 16'h7949;
        src53 <= 16'h659;
        src54 <= 16'h162e;
        src55 <= 16'h1134;
        src56 <= 16'he73;
        src57 <= 16'hc2d9;
        src58 <= 16'h8be3;
        src59 <= 16'h2201;
        src60 <= 16'h38b6;
        src61 <= 16'hbbbc;
        src62 <= 16'h2e1c;
        src63 <= 16'h53d3;
        src64 <= 16'h6b48;
        src65 <= 16'he1da;
        src66 <= 16'hfcf3;
        src67 <= 16'hd4b5;
        src68 <= 16'hd414;
        src69 <= 16'h18f3;
        src70 <= 16'h7c75;
        src71 <= 16'h4c9b;
        src72 <= 16'h8353;
        src73 <= 16'h9ac8;
        src74 <= 16'hecdf;
        src75 <= 16'hd189;
        src76 <= 16'he712;
        src77 <= 16'h940c;
        src78 <= 16'h4c59;
        src79 <= 16'h7e47;
        src80 <= 16'hd0c0;
        src81 <= 16'h42b5;
        src82 <= 16'hc0e0;
        src83 <= 16'h968f;
        src84 <= 16'h878c;
        src85 <= 16'h4b05;
        src86 <= 16'h1c01;
        src87 <= 16'hf282;
        src88 <= 16'h9b2b;
        src89 <= 16'ha903;
        src90 <= 16'he61c;
        src91 <= 16'h6a45;
        src92 <= 16'h3e72;
        src93 <= 16'h6e08;
        src94 <= 16'hb7a7;
        src95 <= 16'h307a;
        src96 <= 16'h8561;
        src97 <= 16'h2961;
        src98 <= 16'h49b4;
        src99 <= 16'hd9b4;
        src100 <= 16'had22;
        src101 <= 16'hde24;
        src102 <= 16'h110a;
        src103 <= 16'he51b;
        src104 <= 16'h203e;
        src105 <= 16'h6acb;
        src106 <= 16'h8776;
        src107 <= 16'h3ca9;
        src108 <= 16'he8f6;
        src109 <= 16'hfb08;
        src110 <= 16'h8dcb;
        src111 <= 16'hcf7f;
        src112 <= 16'hdfcf;
        src113 <= 16'h3896;
        src114 <= 16'h8249;
        src115 <= 16'hfc6b;
        src116 <= 16'he9a4;
        src117 <= 16'hc34;
        src118 <= 16'h60e6;
        src119 <= 16'hec8f;
        src120 <= 16'h3ea0;
        src121 <= 16'hfe10;
        src122 <= 16'hb7ff;
        src123 <= 16'h2e61;
        src124 <= 16'h87d9;
        src125 <= 16'h7eb5;
        src126 <= 16'h4fe7;
        src127 <= 16'hc575;
        src128 <= 16'h82e;
        src129 <= 16'hc058;
        src130 <= 16'h23e8;
        src131 <= 16'hecfb;
        src132 <= 16'h7ff7;
        src133 <= 16'hadf0;
        src134 <= 16'h4324;
        src135 <= 16'h3f54;
        src136 <= 16'hb36f;
        src137 <= 16'h6163;
        src138 <= 16'hafe7;
        src139 <= 16'hb79e;
        src140 <= 16'hb8c6;
        src141 <= 16'h6ab7;
        src142 <= 16'hde4f;
        src143 <= 16'hc015;
        src144 <= 16'h7bbe;
        src145 <= 16'h3aa4;
        src146 <= 16'hc662;
        src147 <= 16'h8d0b;
        src148 <= 16'h287f;
        src149 <= 16'hae26;
        src150 <= 16'hb1c5;
        src151 <= 16'hbd38;
        src152 <= 16'hfb3e;
        src153 <= 16'h2af7;
        src154 <= 16'h5228;
        src155 <= 16'h173f;
        src156 <= 16'hfeda;
        src157 <= 16'heedf;
        src158 <= 16'hd603;
        src159 <= 16'ha86f;
        src160 <= 16'h5871;
        src161 <= 16'h10dc;
        src162 <= 16'h91e1;
        src163 <= 16'h2e07;
        src164 <= 16'h7832;
        src165 <= 16'h8705;
        src166 <= 16'hde8c;
        src167 <= 16'h8fb9;
        src168 <= 16'h73bc;
        src169 <= 16'hb5fd;
        src170 <= 16'hd2d;
        src171 <= 16'hfb9b;
        src172 <= 16'h22c2;
        src173 <= 16'hd63b;
        src174 <= 16'hc736;
        src175 <= 16'h5941;
        src176 <= 16'hb805;
        src177 <= 16'h6ad9;
        src178 <= 16'h422b;
        src179 <= 16'h27a8;
        src180 <= 16'hdbe4;
        src181 <= 16'h6877;
        src182 <= 16'h51cc;
        src183 <= 16'h92cc;
        src184 <= 16'h4d5b;
        exp <= 24'h610244;
        #1
        src0 <= 16'he3fd;
        src1 <= 16'hea0f;
        src2 <= 16'hf486;
        src3 <= 16'hd9b8;
        src4 <= 16'h5fea;
        src5 <= 16'h5b10;
        src6 <= 16'h3a24;
        src7 <= 16'had32;
        src8 <= 16'h9179;
        src9 <= 16'h9f8d;
        src10 <= 16'he0d9;
        src11 <= 16'ha195;
        src12 <= 16'h3474;
        src13 <= 16'h1223;
        src14 <= 16'heaa;
        src15 <= 16'haa2a;
        src16 <= 16'he590;
        src17 <= 16'h6c8e;
        src18 <= 16'h72d1;
        src19 <= 16'h478f;
        src20 <= 16'h5d6e;
        src21 <= 16'hbaeb;
        src22 <= 16'h2360;
        src23 <= 16'h9d9e;
        src24 <= 16'hdfe5;
        src25 <= 16'ha3b1;
        src26 <= 16'h3153;
        src27 <= 16'h61fd;
        src28 <= 16'h3447;
        src29 <= 16'h4a50;
        src30 <= 16'h9cd4;
        src31 <= 16'h2d49;
        src32 <= 16'h26ec;
        src33 <= 16'he217;
        src34 <= 16'h4b06;
        src35 <= 16'ha81a;
        src36 <= 16'he5d1;
        src37 <= 16'hd450;
        src38 <= 16'h7023;
        src39 <= 16'h8db6;
        src40 <= 16'hc710;
        src41 <= 16'h8d64;
        src42 <= 16'h71e2;
        src43 <= 16'h7dbc;
        src44 <= 16'hc697;
        src45 <= 16'h91ca;
        src46 <= 16'hdb74;
        src47 <= 16'h4811;
        src48 <= 16'hf72d;
        src49 <= 16'h906a;
        src50 <= 16'h2d59;
        src51 <= 16'h4dd3;
        src52 <= 16'hf349;
        src53 <= 16'h29f8;
        src54 <= 16'h6550;
        src55 <= 16'h2afe;
        src56 <= 16'hea62;
        src57 <= 16'h642c;
        src58 <= 16'h311a;
        src59 <= 16'hb342;
        src60 <= 16'he574;
        src61 <= 16'hba41;
        src62 <= 16'h1f71;
        src63 <= 16'h6733;
        src64 <= 16'h81b6;
        src65 <= 16'h4035;
        src66 <= 16'hdf9;
        src67 <= 16'hd22;
        src68 <= 16'he56;
        src69 <= 16'h4393;
        src70 <= 16'h35d9;
        src71 <= 16'hcbb4;
        src72 <= 16'hdcae;
        src73 <= 16'h274;
        src74 <= 16'h4772;
        src75 <= 16'h90f2;
        src76 <= 16'h3472;
        src77 <= 16'h2aa7;
        src78 <= 16'h411b;
        src79 <= 16'hf33a;
        src80 <= 16'hd37;
        src81 <= 16'h53b2;
        src82 <= 16'hd888;
        src83 <= 16'h93ce;
        src84 <= 16'hfe94;
        src85 <= 16'h9adb;
        src86 <= 16'h80ab;
        src87 <= 16'h7a5c;
        src88 <= 16'h982b;
        src89 <= 16'hcf87;
        src90 <= 16'h5b5c;
        src91 <= 16'h5ce1;
        src92 <= 16'h17ae;
        src93 <= 16'h43e1;
        src94 <= 16'h82fa;
        src95 <= 16'h9462;
        src96 <= 16'hae87;
        src97 <= 16'h1470;
        src98 <= 16'hb85d;
        src99 <= 16'h8d5b;
        src100 <= 16'h51ac;
        src101 <= 16'h5b37;
        src102 <= 16'h4338;
        src103 <= 16'h91e7;
        src104 <= 16'hce85;
        src105 <= 16'hb171;
        src106 <= 16'h1228;
        src107 <= 16'h913;
        src108 <= 16'hb374;
        src109 <= 16'h2a40;
        src110 <= 16'h4de4;
        src111 <= 16'hecbd;
        src112 <= 16'h7226;
        src113 <= 16'h2fb0;
        src114 <= 16'h5ec;
        src115 <= 16'h9b15;
        src116 <= 16'h1282;
        src117 <= 16'h3227;
        src118 <= 16'he29f;
        src119 <= 16'h6740;
        src120 <= 16'h2ceb;
        src121 <= 16'h5760;
        src122 <= 16'he21f;
        src123 <= 16'ha46f;
        src124 <= 16'h8636;
        src125 <= 16'h2471;
        src126 <= 16'h7715;
        src127 <= 16'hc5c4;
        src128 <= 16'h5208;
        src129 <= 16'h5280;
        src130 <= 16'h4e3c;
        src131 <= 16'hbf4a;
        src132 <= 16'h5743;
        src133 <= 16'he48a;
        src134 <= 16'hd833;
        src135 <= 16'h2ae6;
        src136 <= 16'ha166;
        src137 <= 16'ha96;
        src138 <= 16'h5fcd;
        src139 <= 16'h3d25;
        src140 <= 16'hb430;
        src141 <= 16'hc79d;
        src142 <= 16'ha782;
        src143 <= 16'h8d3e;
        src144 <= 16'h61e5;
        src145 <= 16'h528d;
        src146 <= 16'had0b;
        src147 <= 16'h9a4e;
        src148 <= 16'h96d2;
        src149 <= 16'hab0a;
        src150 <= 16'hbc64;
        src151 <= 16'h51e3;
        src152 <= 16'hf1d8;
        src153 <= 16'hd179;
        src154 <= 16'hdf38;
        src155 <= 16'hd6be;
        src156 <= 16'h1a00;
        src157 <= 16'hf39;
        src158 <= 16'hf9fd;
        src159 <= 16'h942c;
        src160 <= 16'h464c;
        src161 <= 16'h8e6c;
        src162 <= 16'hc445;
        src163 <= 16'hdadc;
        src164 <= 16'ha369;
        src165 <= 16'h4c18;
        src166 <= 16'hf44a;
        src167 <= 16'hf0c0;
        src168 <= 16'h32e8;
        src169 <= 16'hb9d8;
        src170 <= 16'h3162;
        src171 <= 16'hc960;
        src172 <= 16'h37af;
        src173 <= 16'h26a;
        src174 <= 16'ha5b2;
        src175 <= 16'h5717;
        src176 <= 16'he7f4;
        src177 <= 16'h1f1;
        src178 <= 16'h6c12;
        src179 <= 16'h6fa6;
        src180 <= 16'hd12b;
        src181 <= 16'h7668;
        src182 <= 16'h8249;
        src183 <= 16'h1e93;
        src184 <= 16'h1e8e;
        exp <= 24'h5ac0e8;
        #1
        src0 <= 16'h7e2b;
        src1 <= 16'h774e;
        src2 <= 16'hf236;
        src3 <= 16'h18bf;
        src4 <= 16'hc011;
        src5 <= 16'hc88f;
        src6 <= 16'h13a0;
        src7 <= 16'h222e;
        src8 <= 16'h428a;
        src9 <= 16'h1058;
        src10 <= 16'h6b32;
        src11 <= 16'h491e;
        src12 <= 16'h5e72;
        src13 <= 16'ha58b;
        src14 <= 16'haf0d;
        src15 <= 16'hb77b;
        src16 <= 16'h661f;
        src17 <= 16'ha361;
        src18 <= 16'h16;
        src19 <= 16'h2b98;
        src20 <= 16'h648b;
        src21 <= 16'h9abb;
        src22 <= 16'h27e3;
        src23 <= 16'h9bc7;
        src24 <= 16'hffec;
        src25 <= 16'h4d7;
        src26 <= 16'h6e11;
        src27 <= 16'hf14b;
        src28 <= 16'h90cc;
        src29 <= 16'h92b8;
        src30 <= 16'h6db3;
        src31 <= 16'h34c0;
        src32 <= 16'h65ef;
        src33 <= 16'hbc4a;
        src34 <= 16'h46db;
        src35 <= 16'h4dd2;
        src36 <= 16'h8ce8;
        src37 <= 16'h814c;
        src38 <= 16'h70c1;
        src39 <= 16'hb8b1;
        src40 <= 16'hd7c8;
        src41 <= 16'h46da;
        src42 <= 16'hc14c;
        src43 <= 16'h58f;
        src44 <= 16'hc43d;
        src45 <= 16'hc85d;
        src46 <= 16'h68da;
        src47 <= 16'hf6db;
        src48 <= 16'ha313;
        src49 <= 16'h6c7d;
        src50 <= 16'h4d72;
        src51 <= 16'h816e;
        src52 <= 16'h881c;
        src53 <= 16'h3720;
        src54 <= 16'h7b62;
        src55 <= 16'h4471;
        src56 <= 16'hee06;
        src57 <= 16'h9f77;
        src58 <= 16'hcd96;
        src59 <= 16'hc372;
        src60 <= 16'h96ce;
        src61 <= 16'hf057;
        src62 <= 16'h7b7f;
        src63 <= 16'h89bf;
        src64 <= 16'hce56;
        src65 <= 16'h1a63;
        src66 <= 16'h1a71;
        src67 <= 16'h84e3;
        src68 <= 16'h6dec;
        src69 <= 16'h55e1;
        src70 <= 16'h58a8;
        src71 <= 16'hfac2;
        src72 <= 16'h5b20;
        src73 <= 16'hdf69;
        src74 <= 16'hc82f;
        src75 <= 16'h3909;
        src76 <= 16'h14eb;
        src77 <= 16'h3eee;
        src78 <= 16'h4779;
        src79 <= 16'h6535;
        src80 <= 16'h3883;
        src81 <= 16'hc225;
        src82 <= 16'h28ee;
        src83 <= 16'haa3e;
        src84 <= 16'hd1c4;
        src85 <= 16'h57a3;
        src86 <= 16'h38ef;
        src87 <= 16'h821c;
        src88 <= 16'h2067;
        src89 <= 16'hbe6d;
        src90 <= 16'h3056;
        src91 <= 16'h9b3a;
        src92 <= 16'hd0a;
        src93 <= 16'h998e;
        src94 <= 16'h8b43;
        src95 <= 16'h813;
        src96 <= 16'h4f95;
        src97 <= 16'haca7;
        src98 <= 16'h1bb1;
        src99 <= 16'h3e0c;
        src100 <= 16'hf48a;
        src101 <= 16'hc5de;
        src102 <= 16'ha1f1;
        src103 <= 16'h48ec;
        src104 <= 16'hd392;
        src105 <= 16'ha872;
        src106 <= 16'h2f00;
        src107 <= 16'h682;
        src108 <= 16'h52e6;
        src109 <= 16'hc33e;
        src110 <= 16'h23d8;
        src111 <= 16'ha9de;
        src112 <= 16'hd48d;
        src113 <= 16'h3a7c;
        src114 <= 16'h19da;
        src115 <= 16'hc04b;
        src116 <= 16'h6844;
        src117 <= 16'h7ff3;
        src118 <= 16'h8029;
        src119 <= 16'hf006;
        src120 <= 16'h1174;
        src121 <= 16'hdee1;
        src122 <= 16'hf113;
        src123 <= 16'h5495;
        src124 <= 16'ha5c3;
        src125 <= 16'h4dd6;
        src126 <= 16'h6ba0;
        src127 <= 16'h8fb;
        src128 <= 16'hc797;
        src129 <= 16'hc062;
        src130 <= 16'h9e23;
        src131 <= 16'hbf50;
        src132 <= 16'h55b;
        src133 <= 16'hadb9;
        src134 <= 16'h3fbb;
        src135 <= 16'h7415;
        src136 <= 16'h917a;
        src137 <= 16'h6e28;
        src138 <= 16'h401f;
        src139 <= 16'h53ca;
        src140 <= 16'hea20;
        src141 <= 16'hd3b6;
        src142 <= 16'h5bf1;
        src143 <= 16'h351b;
        src144 <= 16'hd083;
        src145 <= 16'h18f;
        src146 <= 16'h3a87;
        src147 <= 16'h666e;
        src148 <= 16'h9396;
        src149 <= 16'hfd7;
        src150 <= 16'h5ecf;
        src151 <= 16'he3bc;
        src152 <= 16'hddc7;
        src153 <= 16'h6ccb;
        src154 <= 16'h3449;
        src155 <= 16'h5c72;
        src156 <= 16'h45a5;
        src157 <= 16'hf85a;
        src158 <= 16'hdaef;
        src159 <= 16'h9fdf;
        src160 <= 16'ha4f8;
        src161 <= 16'h7d3c;
        src162 <= 16'h83dd;
        src163 <= 16'h2e2d;
        src164 <= 16'hcdbc;
        src165 <= 16'h77f6;
        src166 <= 16'ha4ae;
        src167 <= 16'h118f;
        src168 <= 16'h6033;
        src169 <= 16'ha509;
        src170 <= 16'h48d4;
        src171 <= 16'hc293;
        src172 <= 16'hfee7;
        src173 <= 16'h9293;
        src174 <= 16'h53c6;
        src175 <= 16'he7f7;
        src176 <= 16'h62d2;
        src177 <= 16'hc146;
        src178 <= 16'h2bee;
        src179 <= 16'h1019;
        src180 <= 16'ha5e9;
        src181 <= 16'h1dd7;
        src182 <= 16'h7166;
        src183 <= 16'h45e6;
        src184 <= 16'h672;
        exp <= 24'h58a987;
        #1
        src0 <= 16'hc2ab;
        src1 <= 16'h5815;
        src2 <= 16'h2076;
        src3 <= 16'h1530;
        src4 <= 16'h6c0b;
        src5 <= 16'h6903;
        src6 <= 16'h4cfb;
        src7 <= 16'h3e6b;
        src8 <= 16'h2e64;
        src9 <= 16'heb72;
        src10 <= 16'he365;
        src11 <= 16'h3038;
        src12 <= 16'h45bb;
        src13 <= 16'h3e52;
        src14 <= 16'ha76d;
        src15 <= 16'h81f5;
        src16 <= 16'h8667;
        src17 <= 16'h39d5;
        src18 <= 16'hedf8;
        src19 <= 16'hf873;
        src20 <= 16'h9ee7;
        src21 <= 16'h13d7;
        src22 <= 16'h3e39;
        src23 <= 16'h21e2;
        src24 <= 16'h9544;
        src25 <= 16'h6025;
        src26 <= 16'h55bd;
        src27 <= 16'h93cb;
        src28 <= 16'h8d55;
        src29 <= 16'h81ab;
        src30 <= 16'h8ce4;
        src31 <= 16'h1dcf;
        src32 <= 16'h3676;
        src33 <= 16'hdebc;
        src34 <= 16'h9776;
        src35 <= 16'hafed;
        src36 <= 16'h1e1e;
        src37 <= 16'h84d2;
        src38 <= 16'he48c;
        src39 <= 16'h9fe1;
        src40 <= 16'ha4de;
        src41 <= 16'h69f6;
        src42 <= 16'h553f;
        src43 <= 16'h5ba2;
        src44 <= 16'h6e21;
        src45 <= 16'h71bc;
        src46 <= 16'h52fa;
        src47 <= 16'hd951;
        src48 <= 16'hb063;
        src49 <= 16'h1dd1;
        src50 <= 16'h3602;
        src51 <= 16'h6822;
        src52 <= 16'h8667;
        src53 <= 16'h2bbd;
        src54 <= 16'h9e76;
        src55 <= 16'hf042;
        src56 <= 16'h48f8;
        src57 <= 16'h713e;
        src58 <= 16'h3590;
        src59 <= 16'h6b90;
        src60 <= 16'h12fe;
        src61 <= 16'h30d9;
        src62 <= 16'h26ed;
        src63 <= 16'h7aeb;
        src64 <= 16'h2a8;
        src65 <= 16'h7109;
        src66 <= 16'h92c6;
        src67 <= 16'h22a4;
        src68 <= 16'hb82d;
        src69 <= 16'h9779;
        src70 <= 16'hbf35;
        src71 <= 16'h2b4a;
        src72 <= 16'hf293;
        src73 <= 16'h84c7;
        src74 <= 16'h6460;
        src75 <= 16'he908;
        src76 <= 16'h6ff7;
        src77 <= 16'h3dad;
        src78 <= 16'h5376;
        src79 <= 16'hc65c;
        src80 <= 16'h3088;
        src81 <= 16'hc6bd;
        src82 <= 16'hf1a9;
        src83 <= 16'h6f69;
        src84 <= 16'h1b45;
        src85 <= 16'hd2ea;
        src86 <= 16'h3f44;
        src87 <= 16'hc2d;
        src88 <= 16'h7455;
        src89 <= 16'he82f;
        src90 <= 16'hf45c;
        src91 <= 16'h5691;
        src92 <= 16'hc6ff;
        src93 <= 16'h679f;
        src94 <= 16'h5f27;
        src95 <= 16'h5a81;
        src96 <= 16'h55dd;
        src97 <= 16'h23b2;
        src98 <= 16'h677c;
        src99 <= 16'h804;
        src100 <= 16'h3078;
        src101 <= 16'hcf5d;
        src102 <= 16'h7bc1;
        src103 <= 16'hd85;
        src104 <= 16'hcef9;
        src105 <= 16'hf54d;
        src106 <= 16'h8534;
        src107 <= 16'h3fdc;
        src108 <= 16'h713c;
        src109 <= 16'h46f0;
        src110 <= 16'hfbc;
        src111 <= 16'hfb97;
        src112 <= 16'h5506;
        src113 <= 16'h1b52;
        src114 <= 16'h5cfe;
        src115 <= 16'h73bd;
        src116 <= 16'h9801;
        src117 <= 16'had5c;
        src118 <= 16'h7f1b;
        src119 <= 16'h4f50;
        src120 <= 16'h54a;
        src121 <= 16'he849;
        src122 <= 16'hb890;
        src123 <= 16'ha21e;
        src124 <= 16'hbf1d;
        src125 <= 16'hd884;
        src126 <= 16'hcc16;
        src127 <= 16'h85cb;
        src128 <= 16'h1b56;
        src129 <= 16'h107e;
        src130 <= 16'h6149;
        src131 <= 16'h5992;
        src132 <= 16'h8519;
        src133 <= 16'h5d63;
        src134 <= 16'hdfe4;
        src135 <= 16'h8987;
        src136 <= 16'h914e;
        src137 <= 16'h10aa;
        src138 <= 16'h7f6e;
        src139 <= 16'h7a4d;
        src140 <= 16'h8b87;
        src141 <= 16'h3088;
        src142 <= 16'h3c14;
        src143 <= 16'h4117;
        src144 <= 16'h9d7;
        src145 <= 16'h78fe;
        src146 <= 16'hdafe;
        src147 <= 16'h80a1;
        src148 <= 16'h8f9c;
        src149 <= 16'hc43c;
        src150 <= 16'hd36c;
        src151 <= 16'hb5b3;
        src152 <= 16'hb317;
        src153 <= 16'habf7;
        src154 <= 16'h1d08;
        src155 <= 16'h3387;
        src156 <= 16'he63d;
        src157 <= 16'hdea5;
        src158 <= 16'he5d6;
        src159 <= 16'he46;
        src160 <= 16'h2f63;
        src161 <= 16'haa4a;
        src162 <= 16'h4649;
        src163 <= 16'h89c1;
        src164 <= 16'hc948;
        src165 <= 16'hd862;
        src166 <= 16'hd75c;
        src167 <= 16'h4f1a;
        src168 <= 16'h553b;
        src169 <= 16'h942b;
        src170 <= 16'h761e;
        src171 <= 16'h6d9b;
        src172 <= 16'hfffe;
        src173 <= 16'h530d;
        src174 <= 16'hefb9;
        src175 <= 16'h5dfb;
        src176 <= 16'h1a30;
        src177 <= 16'h854;
        src178 <= 16'h6f3;
        src179 <= 16'h4391;
        src180 <= 16'hecc;
        src181 <= 16'h6c27;
        src182 <= 16'h1905;
        src183 <= 16'h33b5;
        src184 <= 16'he7e6;
        exp <= 24'h559a84;
        #1
        src0 <= 16'hc3ee;
        src1 <= 16'hab68;
        src2 <= 16'hcbcc;
        src3 <= 16'h66c9;
        src4 <= 16'h1347;
        src5 <= 16'h105;
        src6 <= 16'h6e1b;
        src7 <= 16'h1b1d;
        src8 <= 16'hbc89;
        src9 <= 16'h6c07;
        src10 <= 16'hd5b6;
        src11 <= 16'hf01;
        src12 <= 16'h83f7;
        src13 <= 16'h3dc8;
        src14 <= 16'h12b0;
        src15 <= 16'hb5c0;
        src16 <= 16'h3e1d;
        src17 <= 16'he3bd;
        src18 <= 16'h10fa;
        src19 <= 16'h951b;
        src20 <= 16'he03c;
        src21 <= 16'h4d88;
        src22 <= 16'h22e7;
        src23 <= 16'h47e4;
        src24 <= 16'h7367;
        src25 <= 16'heb42;
        src26 <= 16'hfb0;
        src27 <= 16'hd108;
        src28 <= 16'h2b75;
        src29 <= 16'h92f6;
        src30 <= 16'h4a9d;
        src31 <= 16'h40ab;
        src32 <= 16'hda20;
        src33 <= 16'ha320;
        src34 <= 16'h29e6;
        src35 <= 16'h2efa;
        src36 <= 16'hca46;
        src37 <= 16'h1ae3;
        src38 <= 16'hc203;
        src39 <= 16'hc5b2;
        src40 <= 16'h340f;
        src41 <= 16'hefa4;
        src42 <= 16'h70d6;
        src43 <= 16'he09e;
        src44 <= 16'h6270;
        src45 <= 16'hc20;
        src46 <= 16'ha682;
        src47 <= 16'h534d;
        src48 <= 16'h8cb8;
        src49 <= 16'hb228;
        src50 <= 16'h9276;
        src51 <= 16'h2104;
        src52 <= 16'he7b7;
        src53 <= 16'ha580;
        src54 <= 16'hc310;
        src55 <= 16'h3b28;
        src56 <= 16'h286b;
        src57 <= 16'h263a;
        src58 <= 16'h2f16;
        src59 <= 16'hc64d;
        src60 <= 16'h8e36;
        src61 <= 16'h8d57;
        src62 <= 16'h7948;
        src63 <= 16'heda4;
        src64 <= 16'hf430;
        src65 <= 16'hd57e;
        src66 <= 16'h90f6;
        src67 <= 16'hf609;
        src68 <= 16'hf4ca;
        src69 <= 16'h553c;
        src70 <= 16'h2b96;
        src71 <= 16'hbf65;
        src72 <= 16'h4bc3;
        src73 <= 16'h27c5;
        src74 <= 16'hc194;
        src75 <= 16'h4c97;
        src76 <= 16'hf200;
        src77 <= 16'h847;
        src78 <= 16'h249;
        src79 <= 16'h2894;
        src80 <= 16'hbeb;
        src81 <= 16'h5251;
        src82 <= 16'h7bd8;
        src83 <= 16'h49f3;
        src84 <= 16'hba52;
        src85 <= 16'h23be;
        src86 <= 16'h44b9;
        src87 <= 16'haabe;
        src88 <= 16'hb670;
        src89 <= 16'hf5aa;
        src90 <= 16'h829e;
        src91 <= 16'hae70;
        src92 <= 16'h78e1;
        src93 <= 16'h2ac9;
        src94 <= 16'h5fb3;
        src95 <= 16'h20b2;
        src96 <= 16'hb390;
        src97 <= 16'h6ab9;
        src98 <= 16'hd12f;
        src99 <= 16'h86f;
        src100 <= 16'h123f;
        src101 <= 16'h4319;
        src102 <= 16'h5c55;
        src103 <= 16'h65b8;
        src104 <= 16'h86bd;
        src105 <= 16'he3f2;
        src106 <= 16'he35c;
        src107 <= 16'h41ca;
        src108 <= 16'h261f;
        src109 <= 16'he93;
        src110 <= 16'h1a67;
        src111 <= 16'he22f;
        src112 <= 16'h9c35;
        src113 <= 16'hb73b;
        src114 <= 16'h5eab;
        src115 <= 16'he252;
        src116 <= 16'h1021;
        src117 <= 16'hd0a8;
        src118 <= 16'h66b3;
        src119 <= 16'h7728;
        src120 <= 16'hac59;
        src121 <= 16'hf3e5;
        src122 <= 16'hc903;
        src123 <= 16'hde89;
        src124 <= 16'he221;
        src125 <= 16'h60fe;
        src126 <= 16'hbf76;
        src127 <= 16'ha5b8;
        src128 <= 16'h968c;
        src129 <= 16'h616;
        src130 <= 16'h9cc3;
        src131 <= 16'h27f9;
        src132 <= 16'ha365;
        src133 <= 16'hdd49;
        src134 <= 16'hf2ca;
        src135 <= 16'hbf73;
        src136 <= 16'h84f4;
        src137 <= 16'h8d67;
        src138 <= 16'h8936;
        src139 <= 16'h86d0;
        src140 <= 16'hc2c0;
        src141 <= 16'he620;
        src142 <= 16'hddba;
        src143 <= 16'h2b41;
        src144 <= 16'hd4b5;
        src145 <= 16'h8570;
        src146 <= 16'he3fa;
        src147 <= 16'h3f27;
        src148 <= 16'hc1a2;
        src149 <= 16'h71d9;
        src150 <= 16'h3ddc;
        src151 <= 16'h1119;
        src152 <= 16'hdf67;
        src153 <= 16'hdcc4;
        src154 <= 16'hde3e;
        src155 <= 16'habc4;
        src156 <= 16'h2052;
        src157 <= 16'h2646;
        src158 <= 16'ha346;
        src159 <= 16'hd409;
        src160 <= 16'h9cc8;
        src161 <= 16'h5734;
        src162 <= 16'h91b0;
        src163 <= 16'h84e2;
        src164 <= 16'hfb6;
        src165 <= 16'hc2ab;
        src166 <= 16'h136c;
        src167 <= 16'hd28a;
        src168 <= 16'hbd72;
        src169 <= 16'h389d;
        src170 <= 16'hf812;
        src171 <= 16'h819a;
        src172 <= 16'haf1e;
        src173 <= 16'h1ecd;
        src174 <= 16'hbee5;
        src175 <= 16'h4c0e;
        src176 <= 16'h3260;
        src177 <= 16'h8549;
        src178 <= 16'h1ab3;
        src179 <= 16'h8ac0;
        src180 <= 16'h3fa1;
        src181 <= 16'hf23f;
        src182 <= 16'h686;
        src183 <= 16'h193c;
        src184 <= 16'h9acd;
        exp <= 24'h5c1978;
        #1
        src0 <= 16'hb67d;
        src1 <= 16'h792c;
        src2 <= 16'h9bb1;
        src3 <= 16'h68a;
        src4 <= 16'h25e3;
        src5 <= 16'h9bbd;
        src6 <= 16'haaf0;
        src7 <= 16'he16f;
        src8 <= 16'h64d4;
        src9 <= 16'hb30e;
        src10 <= 16'hb964;
        src11 <= 16'h9eed;
        src12 <= 16'he1c;
        src13 <= 16'h67be;
        src14 <= 16'ha02;
        src15 <= 16'h7238;
        src16 <= 16'hbe56;
        src17 <= 16'hf6aa;
        src18 <= 16'ha6dd;
        src19 <= 16'h78e1;
        src20 <= 16'h7c22;
        src21 <= 16'h7c84;
        src22 <= 16'h4c7b;
        src23 <= 16'h864e;
        src24 <= 16'he982;
        src25 <= 16'h4b7c;
        src26 <= 16'hda82;
        src27 <= 16'h97ed;
        src28 <= 16'ha88d;
        src29 <= 16'he84e;
        src30 <= 16'h2edd;
        src31 <= 16'h954d;
        src32 <= 16'h9a4e;
        src33 <= 16'h8c0f;
        src34 <= 16'h32f6;
        src35 <= 16'he87d;
        src36 <= 16'h3103;
        src37 <= 16'h5dc3;
        src38 <= 16'h9fae;
        src39 <= 16'ha0db;
        src40 <= 16'h8746;
        src41 <= 16'hb16c;
        src42 <= 16'ha63d;
        src43 <= 16'h6c8b;
        src44 <= 16'h883c;
        src45 <= 16'h7ac6;
        src46 <= 16'h9b45;
        src47 <= 16'hdf21;
        src48 <= 16'hdead;
        src49 <= 16'ha259;
        src50 <= 16'h8dd6;
        src51 <= 16'hf125;
        src52 <= 16'h1c90;
        src53 <= 16'ha6fb;
        src54 <= 16'h5f5a;
        src55 <= 16'hc137;
        src56 <= 16'h92d4;
        src57 <= 16'h3d9d;
        src58 <= 16'hb0eb;
        src59 <= 16'ha2bc;
        src60 <= 16'h5223;
        src61 <= 16'hdd79;
        src62 <= 16'he649;
        src63 <= 16'h39ad;
        src64 <= 16'hec3b;
        src65 <= 16'h774;
        src66 <= 16'h1580;
        src67 <= 16'h7b8e;
        src68 <= 16'ha869;
        src69 <= 16'h897;
        src70 <= 16'h20e6;
        src71 <= 16'hc92f;
        src72 <= 16'h6cab;
        src73 <= 16'hefff;
        src74 <= 16'h97ce;
        src75 <= 16'h3e99;
        src76 <= 16'h290d;
        src77 <= 16'hf5ff;
        src78 <= 16'hd810;
        src79 <= 16'h54ea;
        src80 <= 16'h59f4;
        src81 <= 16'ha443;
        src82 <= 16'hb370;
        src83 <= 16'hd1af;
        src84 <= 16'ha796;
        src85 <= 16'hdabf;
        src86 <= 16'hba7c;
        src87 <= 16'hefc9;
        src88 <= 16'h83aa;
        src89 <= 16'he2a7;
        src90 <= 16'hee1a;
        src91 <= 16'h7ef9;
        src92 <= 16'h9624;
        src93 <= 16'h8398;
        src94 <= 16'h74ce;
        src95 <= 16'hafa4;
        src96 <= 16'hd20a;
        src97 <= 16'h68e0;
        src98 <= 16'h347;
        src99 <= 16'hc0a7;
        src100 <= 16'h163a;
        src101 <= 16'h171c;
        src102 <= 16'hc222;
        src103 <= 16'hfa1e;
        src104 <= 16'hf585;
        src105 <= 16'h37e4;
        src106 <= 16'hde53;
        src107 <= 16'h1539;
        src108 <= 16'he57e;
        src109 <= 16'h57da;
        src110 <= 16'h64e;
        src111 <= 16'h2ab8;
        src112 <= 16'hbef5;
        src113 <= 16'h3827;
        src114 <= 16'h8c9d;
        src115 <= 16'h5402;
        src116 <= 16'h7f73;
        src117 <= 16'hd073;
        src118 <= 16'h1ca2;
        src119 <= 16'hbfe1;
        src120 <= 16'h71c1;
        src121 <= 16'h6be7;
        src122 <= 16'h357f;
        src123 <= 16'h9518;
        src124 <= 16'hc373;
        src125 <= 16'h60c3;
        src126 <= 16'h8a7;
        src127 <= 16'hcec0;
        src128 <= 16'h68df;
        src129 <= 16'h98f5;
        src130 <= 16'hd8d8;
        src131 <= 16'h5201;
        src132 <= 16'hee2e;
        src133 <= 16'hd27d;
        src134 <= 16'h37d7;
        src135 <= 16'ha734;
        src136 <= 16'hde21;
        src137 <= 16'h4fac;
        src138 <= 16'h778;
        src139 <= 16'h755d;
        src140 <= 16'hd7af;
        src141 <= 16'h3cd7;
        src142 <= 16'h1449;
        src143 <= 16'h4f03;
        src144 <= 16'h9e7;
        src145 <= 16'hbac1;
        src146 <= 16'h5ddf;
        src147 <= 16'hbac7;
        src148 <= 16'hcf17;
        src149 <= 16'hd46;
        src150 <= 16'h3c7f;
        src151 <= 16'hc645;
        src152 <= 16'h9d99;
        src153 <= 16'h54a2;
        src154 <= 16'hc6ed;
        src155 <= 16'h3461;
        src156 <= 16'ha14f;
        src157 <= 16'h3fce;
        src158 <= 16'hec8d;
        src159 <= 16'h490f;
        src160 <= 16'h156c;
        src161 <= 16'ha195;
        src162 <= 16'h3142;
        src163 <= 16'h74a0;
        src164 <= 16'h5adb;
        src165 <= 16'h8184;
        src166 <= 16'h50fb;
        src167 <= 16'ha0ab;
        src168 <= 16'hebb8;
        src169 <= 16'h51e9;
        src170 <= 16'h63ff;
        src171 <= 16'hd21b;
        src172 <= 16'he694;
        src173 <= 16'h809b;
        src174 <= 16'h3859;
        src175 <= 16'h315b;
        src176 <= 16'h77e;
        src177 <= 16'ha0f9;
        src178 <= 16'h5902;
        src179 <= 16'hb1ee;
        src180 <= 16'h6a15;
        src181 <= 16'ha8c1;
        src182 <= 16'hdeab;
        src183 <= 16'hcf85;
        src184 <= 16'hf802;
        exp <= 24'h615c3a;
        #1
        src0 <= 16'h89bf;
        src1 <= 16'haa06;
        src2 <= 16'h81a5;
        src3 <= 16'h6b75;
        src4 <= 16'h9105;
        src5 <= 16'h2784;
        src6 <= 16'hd8b9;
        src7 <= 16'h87a1;
        src8 <= 16'hbeb4;
        src9 <= 16'ha535;
        src10 <= 16'hde30;
        src11 <= 16'h8ba0;
        src12 <= 16'h836f;
        src13 <= 16'h5b66;
        src14 <= 16'h7a1c;
        src15 <= 16'h4caa;
        src16 <= 16'h4a61;
        src17 <= 16'hfaac;
        src18 <= 16'h3a5;
        src19 <= 16'h303;
        src20 <= 16'h7637;
        src21 <= 16'h52bf;
        src22 <= 16'hcf4f;
        src23 <= 16'h96c1;
        src24 <= 16'hffac;
        src25 <= 16'hf2ad;
        src26 <= 16'ha6d9;
        src27 <= 16'he1ed;
        src28 <= 16'hb1a3;
        src29 <= 16'h423;
        src30 <= 16'he578;
        src31 <= 16'h32b3;
        src32 <= 16'h4e5f;
        src33 <= 16'hcfbd;
        src34 <= 16'hf16b;
        src35 <= 16'h21a5;
        src36 <= 16'ha343;
        src37 <= 16'hbfe;
        src38 <= 16'h672f;
        src39 <= 16'hc3c0;
        src40 <= 16'h3c9a;
        src41 <= 16'h69ef;
        src42 <= 16'hdf8c;
        src43 <= 16'h2d05;
        src44 <= 16'h5b87;
        src45 <= 16'h8b7d;
        src46 <= 16'h8374;
        src47 <= 16'h43ed;
        src48 <= 16'h288a;
        src49 <= 16'h4c0c;
        src50 <= 16'hd423;
        src51 <= 16'h8b57;
        src52 <= 16'h2ad7;
        src53 <= 16'he6c4;
        src54 <= 16'hee13;
        src55 <= 16'hf1a0;
        src56 <= 16'h5ecb;
        src57 <= 16'hd21a;
        src58 <= 16'h8c65;
        src59 <= 16'h5f4f;
        src60 <= 16'h7884;
        src61 <= 16'h352d;
        src62 <= 16'hc30;
        src63 <= 16'h7617;
        src64 <= 16'hc074;
        src65 <= 16'hb61f;
        src66 <= 16'h87f4;
        src67 <= 16'h3f9d;
        src68 <= 16'h776a;
        src69 <= 16'hec4c;
        src70 <= 16'h1e8d;
        src71 <= 16'h2bcd;
        src72 <= 16'h1004;
        src73 <= 16'h83ef;
        src74 <= 16'h4cee;
        src75 <= 16'h42df;
        src76 <= 16'hc318;
        src77 <= 16'h2b51;
        src78 <= 16'h8add;
        src79 <= 16'h7402;
        src80 <= 16'ha3b;
        src81 <= 16'ha892;
        src82 <= 16'h23f0;
        src83 <= 16'h8971;
        src84 <= 16'hed68;
        src85 <= 16'hf647;
        src86 <= 16'h9369;
        src87 <= 16'hd0b;
        src88 <= 16'h8f6d;
        src89 <= 16'h3613;
        src90 <= 16'h1b1b;
        src91 <= 16'hd9b0;
        src92 <= 16'hd437;
        src93 <= 16'h7590;
        src94 <= 16'hd838;
        src95 <= 16'hb3d3;
        src96 <= 16'h13e8;
        src97 <= 16'h6412;
        src98 <= 16'h3d87;
        src99 <= 16'h73dc;
        src100 <= 16'h414b;
        src101 <= 16'ha04c;
        src102 <= 16'h5d41;
        src103 <= 16'h8141;
        src104 <= 16'hbbc8;
        src105 <= 16'h1a0;
        src106 <= 16'hed4b;
        src107 <= 16'h21ab;
        src108 <= 16'h1448;
        src109 <= 16'hca2a;
        src110 <= 16'h2659;
        src111 <= 16'haf9;
        src112 <= 16'h20b8;
        src113 <= 16'h253b;
        src114 <= 16'h5286;
        src115 <= 16'h3993;
        src116 <= 16'h12e3;
        src117 <= 16'h9798;
        src118 <= 16'he8f9;
        src119 <= 16'h3224;
        src120 <= 16'h8114;
        src121 <= 16'h7b0d;
        src122 <= 16'hf1c7;
        src123 <= 16'h9753;
        src124 <= 16'h1f89;
        src125 <= 16'h9e84;
        src126 <= 16'h5633;
        src127 <= 16'hfc1c;
        src128 <= 16'hf518;
        src129 <= 16'h9f68;
        src130 <= 16'h3de2;
        src131 <= 16'h9f1d;
        src132 <= 16'h8269;
        src133 <= 16'h8e48;
        src134 <= 16'hb938;
        src135 <= 16'hcd7a;
        src136 <= 16'h1247;
        src137 <= 16'h17bc;
        src138 <= 16'hdf37;
        src139 <= 16'h78d6;
        src140 <= 16'hc130;
        src141 <= 16'h3acb;
        src142 <= 16'hf439;
        src143 <= 16'h91fd;
        src144 <= 16'hb7da;
        src145 <= 16'h63a4;
        src146 <= 16'h12dc;
        src147 <= 16'h5212;
        src148 <= 16'h2444;
        src149 <= 16'had49;
        src150 <= 16'hfa6b;
        src151 <= 16'h9575;
        src152 <= 16'h8d78;
        src153 <= 16'h755e;
        src154 <= 16'h7766;
        src155 <= 16'h321e;
        src156 <= 16'hbe24;
        src157 <= 16'h1af0;
        src158 <= 16'hb9c6;
        src159 <= 16'h8077;
        src160 <= 16'hf9fa;
        src161 <= 16'h8b79;
        src162 <= 16'h5559;
        src163 <= 16'ha4ff;
        src164 <= 16'h31fd;
        src165 <= 16'hb43d;
        src166 <= 16'h9b16;
        src167 <= 16'ha92a;
        src168 <= 16'h8d31;
        src169 <= 16'h5d8a;
        src170 <= 16'hfab5;
        src171 <= 16'hbac2;
        src172 <= 16'h10d6;
        src173 <= 16'h971e;
        src174 <= 16'h4ef;
        src175 <= 16'hec51;
        src176 <= 16'h8198;
        src177 <= 16'hc48d;
        src178 <= 16'h4d3b;
        src179 <= 16'h92ad;
        src180 <= 16'hfee1;
        src181 <= 16'h4bca;
        src182 <= 16'h6056;
        src183 <= 16'hb61;
        src184 <= 16'h9882;
        exp <= 24'h5b5b6b;
        #1
        src0 <= 16'hc5c9;
        src1 <= 16'hf0ad;
        src2 <= 16'h5de;
        src3 <= 16'h8dec;
        src4 <= 16'h5af6;
        src5 <= 16'h2b8e;
        src6 <= 16'h4da6;
        src7 <= 16'h1cb7;
        src8 <= 16'h44a2;
        src9 <= 16'h334b;
        src10 <= 16'hf7af;
        src11 <= 16'h75ee;
        src12 <= 16'hed94;
        src13 <= 16'hb39a;
        src14 <= 16'h295f;
        src15 <= 16'h5e56;
        src16 <= 16'h84f8;
        src17 <= 16'hf8ae;
        src18 <= 16'hc26a;
        src19 <= 16'he58e;
        src20 <= 16'h7094;
        src21 <= 16'hc542;
        src22 <= 16'hea68;
        src23 <= 16'h5bc5;
        src24 <= 16'hfe6e;
        src25 <= 16'hbc44;
        src26 <= 16'hf9d3;
        src27 <= 16'h1d64;
        src28 <= 16'h2355;
        src29 <= 16'hf483;
        src30 <= 16'hfc81;
        src31 <= 16'h16d1;
        src32 <= 16'hf58c;
        src33 <= 16'h96c6;
        src34 <= 16'hae13;
        src35 <= 16'h31b1;
        src36 <= 16'hfa64;
        src37 <= 16'he598;
        src38 <= 16'hb29e;
        src39 <= 16'h4a22;
        src40 <= 16'ha825;
        src41 <= 16'hf387;
        src42 <= 16'ha318;
        src43 <= 16'h9039;
        src44 <= 16'h8b7e;
        src45 <= 16'h58fc;
        src46 <= 16'h7677;
        src47 <= 16'h4d;
        src48 <= 16'h9bac;
        src49 <= 16'hfb26;
        src50 <= 16'h7;
        src51 <= 16'hc994;
        src52 <= 16'h4de7;
        src53 <= 16'h1fb5;
        src54 <= 16'h3043;
        src55 <= 16'hcf4d;
        src56 <= 16'h8493;
        src57 <= 16'h3ae5;
        src58 <= 16'hf47f;
        src59 <= 16'h8a24;
        src60 <= 16'h267;
        src61 <= 16'h1ac7;
        src62 <= 16'h5eb4;
        src63 <= 16'h2780;
        src64 <= 16'h2067;
        src65 <= 16'hacd8;
        src66 <= 16'h8085;
        src67 <= 16'hb3ff;
        src68 <= 16'h57d0;
        src69 <= 16'h7ae9;
        src70 <= 16'h741;
        src71 <= 16'he91b;
        src72 <= 16'hde1f;
        src73 <= 16'hc4e7;
        src74 <= 16'h48a3;
        src75 <= 16'hf233;
        src76 <= 16'he6de;
        src77 <= 16'heb6f;
        src78 <= 16'h4a65;
        src79 <= 16'hb001;
        src80 <= 16'h6262;
        src81 <= 16'hf542;
        src82 <= 16'h2875;
        src83 <= 16'h1af9;
        src84 <= 16'h1c05;
        src85 <= 16'h8472;
        src86 <= 16'h957;
        src87 <= 16'hee25;
        src88 <= 16'hf3d3;
        src89 <= 16'h502d;
        src90 <= 16'h8bf5;
        src91 <= 16'h12f0;
        src92 <= 16'hd2b5;
        src93 <= 16'h7ef3;
        src94 <= 16'h698;
        src95 <= 16'hc143;
        src96 <= 16'h3bf7;
        src97 <= 16'h24bb;
        src98 <= 16'hc212;
        src99 <= 16'h3baa;
        src100 <= 16'h3a62;
        src101 <= 16'hbebd;
        src102 <= 16'h30de;
        src103 <= 16'hbdc7;
        src104 <= 16'h927b;
        src105 <= 16'hc686;
        src106 <= 16'h6d1d;
        src107 <= 16'h63a8;
        src108 <= 16'h3dca;
        src109 <= 16'hafa;
        src110 <= 16'h98d6;
        src111 <= 16'hc470;
        src112 <= 16'he721;
        src113 <= 16'h6074;
        src114 <= 16'hd9;
        src115 <= 16'h6500;
        src116 <= 16'h1d1b;
        src117 <= 16'h9219;
        src118 <= 16'h70ea;
        src119 <= 16'h58a9;
        src120 <= 16'h6af;
        src121 <= 16'h776f;
        src122 <= 16'h39f9;
        src123 <= 16'hc87d;
        src124 <= 16'hb284;
        src125 <= 16'he862;
        src126 <= 16'hf369;
        src127 <= 16'he5b3;
        src128 <= 16'h9439;
        src129 <= 16'hd559;
        src130 <= 16'h304f;
        src131 <= 16'ha26c;
        src132 <= 16'h9507;
        src133 <= 16'h675a;
        src134 <= 16'h4fac;
        src135 <= 16'h5362;
        src136 <= 16'h72b5;
        src137 <= 16'h6048;
        src138 <= 16'ha68b;
        src139 <= 16'h6cb4;
        src140 <= 16'hdf76;
        src141 <= 16'haf45;
        src142 <= 16'h95d5;
        src143 <= 16'hcd61;
        src144 <= 16'h1b73;
        src145 <= 16'had12;
        src146 <= 16'h8b31;
        src147 <= 16'h9678;
        src148 <= 16'h710d;
        src149 <= 16'h6a4;
        src150 <= 16'hc525;
        src151 <= 16'h63ca;
        src152 <= 16'h255f;
        src153 <= 16'hc072;
        src154 <= 16'h391a;
        src155 <= 16'h6059;
        src156 <= 16'h6fdd;
        src157 <= 16'hf608;
        src158 <= 16'h5e6a;
        src159 <= 16'heb45;
        src160 <= 16'hec25;
        src161 <= 16'h9a35;
        src162 <= 16'h10ae;
        src163 <= 16'h4f76;
        src164 <= 16'hf0a4;
        src165 <= 16'h78d7;
        src166 <= 16'h13ff;
        src167 <= 16'h308e;
        src168 <= 16'h24e8;
        src169 <= 16'h6590;
        src170 <= 16'hf8f8;
        src171 <= 16'hf871;
        src172 <= 16'h908f;
        src173 <= 16'h5962;
        src174 <= 16'h7307;
        src175 <= 16'h53f0;
        src176 <= 16'hd752;
        src177 <= 16'h6e8d;
        src178 <= 16'hd52b;
        src179 <= 16'hb63b;
        src180 <= 16'h4be5;
        src181 <= 16'hdccc;
        src182 <= 16'h3d88;
        src183 <= 16'hb06a;
        src184 <= 16'h19bb;
        exp <= 24'h5f0a87;
        #1
        src0 <= 16'he3dc;
        src1 <= 16'he26a;
        src2 <= 16'h747e;
        src3 <= 16'h56d0;
        src4 <= 16'hec4b;
        src5 <= 16'h81e6;
        src6 <= 16'h5479;
        src7 <= 16'h81a5;
        src8 <= 16'hcfc2;
        src9 <= 16'h887b;
        src10 <= 16'hc221;
        src11 <= 16'hb175;
        src12 <= 16'hc361;
        src13 <= 16'h5b13;
        src14 <= 16'h9a81;
        src15 <= 16'hce96;
        src16 <= 16'h2b57;
        src17 <= 16'hdb08;
        src18 <= 16'h558a;
        src19 <= 16'hb5bc;
        src20 <= 16'haac0;
        src21 <= 16'h29d6;
        src22 <= 16'h7fe0;
        src23 <= 16'h4b16;
        src24 <= 16'h5489;
        src25 <= 16'h9ab4;
        src26 <= 16'hf66a;
        src27 <= 16'hd979;
        src28 <= 16'hc645;
        src29 <= 16'hf893;
        src30 <= 16'h16da;
        src31 <= 16'h40bb;
        src32 <= 16'h7239;
        src33 <= 16'hc892;
        src34 <= 16'h2113;
        src35 <= 16'hb760;
        src36 <= 16'h1e66;
        src37 <= 16'hcabc;
        src38 <= 16'hdb58;
        src39 <= 16'h2597;
        src40 <= 16'h6cbe;
        src41 <= 16'hfe2d;
        src42 <= 16'h9c0a;
        src43 <= 16'hcd57;
        src44 <= 16'h2049;
        src45 <= 16'h40b;
        src46 <= 16'he177;
        src47 <= 16'h28db;
        src48 <= 16'hdf85;
        src49 <= 16'h5dd8;
        src50 <= 16'heed9;
        src51 <= 16'hc41b;
        src52 <= 16'hf7cd;
        src53 <= 16'hc5c0;
        src54 <= 16'hb318;
        src55 <= 16'hadae;
        src56 <= 16'h5905;
        src57 <= 16'hd53d;
        src58 <= 16'hb928;
        src59 <= 16'h72a0;
        src60 <= 16'haad8;
        src61 <= 16'h6458;
        src62 <= 16'hf74;
        src63 <= 16'hcc92;
        src64 <= 16'had51;
        src65 <= 16'haa92;
        src66 <= 16'hf910;
        src67 <= 16'hd4ff;
        src68 <= 16'hf942;
        src69 <= 16'h1fcf;
        src70 <= 16'h3185;
        src71 <= 16'hef;
        src72 <= 16'he28e;
        src73 <= 16'h21e0;
        src74 <= 16'h2559;
        src75 <= 16'hbac2;
        src76 <= 16'h43a4;
        src77 <= 16'h936b;
        src78 <= 16'hcac1;
        src79 <= 16'h187f;
        src80 <= 16'haa81;
        src81 <= 16'he6bb;
        src82 <= 16'h50b8;
        src83 <= 16'h6ecc;
        src84 <= 16'h33e5;
        src85 <= 16'hcd46;
        src86 <= 16'h1428;
        src87 <= 16'hf136;
        src88 <= 16'hb002;
        src89 <= 16'h9c8e;
        src90 <= 16'h2c11;
        src91 <= 16'hecd3;
        src92 <= 16'h99fa;
        src93 <= 16'h2974;
        src94 <= 16'hb5e6;
        src95 <= 16'h7335;
        src96 <= 16'h2700;
        src97 <= 16'h3cd8;
        src98 <= 16'h6d1a;
        src99 <= 16'hdc32;
        src100 <= 16'h8906;
        src101 <= 16'h8577;
        src102 <= 16'h38ae;
        src103 <= 16'h93a4;
        src104 <= 16'h1072;
        src105 <= 16'h3e28;
        src106 <= 16'hbc69;
        src107 <= 16'hcc82;
        src108 <= 16'hf517;
        src109 <= 16'hb87a;
        src110 <= 16'hee5;
        src111 <= 16'h984e;
        src112 <= 16'h745c;
        src113 <= 16'h64e;
        src114 <= 16'hf2c5;
        src115 <= 16'hd267;
        src116 <= 16'h9489;
        src117 <= 16'h62d1;
        src118 <= 16'h12c8;
        src119 <= 16'hf0ab;
        src120 <= 16'h2290;
        src121 <= 16'h6273;
        src122 <= 16'h2801;
        src123 <= 16'h3cb2;
        src124 <= 16'h49ce;
        src125 <= 16'h2988;
        src126 <= 16'hf2b6;
        src127 <= 16'he4bb;
        src128 <= 16'hf655;
        src129 <= 16'h4b31;
        src130 <= 16'h22d9;
        src131 <= 16'h58de;
        src132 <= 16'h55ea;
        src133 <= 16'h80cf;
        src134 <= 16'h5e46;
        src135 <= 16'h3cea;
        src136 <= 16'h7653;
        src137 <= 16'h35a6;
        src138 <= 16'he7fe;
        src139 <= 16'h7090;
        src140 <= 16'hd3c1;
        src141 <= 16'h7fa3;
        src142 <= 16'haf82;
        src143 <= 16'h16d6;
        src144 <= 16'h5a84;
        src145 <= 16'hee6c;
        src146 <= 16'h4a3f;
        src147 <= 16'h68f8;
        src148 <= 16'h6b09;
        src149 <= 16'he51;
        src150 <= 16'h9aa0;
        src151 <= 16'hbab0;
        src152 <= 16'ha79a;
        src153 <= 16'h8ac2;
        src154 <= 16'h84e0;
        src155 <= 16'ha758;
        src156 <= 16'h83e4;
        src157 <= 16'hb31e;
        src158 <= 16'hc6c0;
        src159 <= 16'h5975;
        src160 <= 16'hc0b;
        src161 <= 16'h2578;
        src162 <= 16'hcada;
        src163 <= 16'h98e7;
        src164 <= 16'h9a1a;
        src165 <= 16'hfcf2;
        src166 <= 16'he09d;
        src167 <= 16'h84ae;
        src168 <= 16'h485e;
        src169 <= 16'h69c1;
        src170 <= 16'h4b79;
        src171 <= 16'hc6bc;
        src172 <= 16'h3f43;
        src173 <= 16'h4f34;
        src174 <= 16'h95d3;
        src175 <= 16'h532f;
        src176 <= 16'h11d0;
        src177 <= 16'h6e60;
        src178 <= 16'h7c30;
        src179 <= 16'h25b4;
        src180 <= 16'h8df9;
        src181 <= 16'hb17f;
        src182 <= 16'hfdf;
        src183 <= 16'hf98b;
        src184 <= 16'h358c;
        exp <= 24'h601d04;
        #1
        src0 <= 16'h607e;
        src1 <= 16'h9ef7;
        src2 <= 16'h1cc6;
        src3 <= 16'h2674;
        src4 <= 16'h718b;
        src5 <= 16'hc9ab;
        src6 <= 16'hfc0d;
        src7 <= 16'h52c0;
        src8 <= 16'hc6f1;
        src9 <= 16'hb5d9;
        src10 <= 16'h4e62;
        src11 <= 16'he095;
        src12 <= 16'h5b6a;
        src13 <= 16'h6c03;
        src14 <= 16'hd550;
        src15 <= 16'hf821;
        src16 <= 16'h8135;
        src17 <= 16'h7c43;
        src18 <= 16'h40c;
        src19 <= 16'hd4d6;
        src20 <= 16'h9e0e;
        src21 <= 16'h5ab;
        src22 <= 16'hafe8;
        src23 <= 16'hac19;
        src24 <= 16'h5670;
        src25 <= 16'h78aa;
        src26 <= 16'he735;
        src27 <= 16'hb588;
        src28 <= 16'ha77;
        src29 <= 16'h1c93;
        src30 <= 16'h7c30;
        src31 <= 16'hab89;
        src32 <= 16'hd622;
        src33 <= 16'h469a;
        src34 <= 16'hb3d0;
        src35 <= 16'hada5;
        src36 <= 16'h1a02;
        src37 <= 16'h95bb;
        src38 <= 16'hd91;
        src39 <= 16'hbff9;
        src40 <= 16'h474b;
        src41 <= 16'h4565;
        src42 <= 16'h6320;
        src43 <= 16'h74cb;
        src44 <= 16'hd9c4;
        src45 <= 16'hcb99;
        src46 <= 16'hf9a7;
        src47 <= 16'h75d5;
        src48 <= 16'haa36;
        src49 <= 16'head2;
        src50 <= 16'h1e18;
        src51 <= 16'h8116;
        src52 <= 16'ha5c9;
        src53 <= 16'h166;
        src54 <= 16'h6f09;
        src55 <= 16'he8a6;
        src56 <= 16'ha45a;
        src57 <= 16'hd0cc;
        src58 <= 16'hd97;
        src59 <= 16'h927d;
        src60 <= 16'h21ec;
        src61 <= 16'he6db;
        src62 <= 16'hd741;
        src63 <= 16'h8453;
        src64 <= 16'h58d0;
        src65 <= 16'hba16;
        src66 <= 16'hd4fa;
        src67 <= 16'he3b0;
        src68 <= 16'h46eb;
        src69 <= 16'hfee3;
        src70 <= 16'h65e6;
        src71 <= 16'h3fb7;
        src72 <= 16'hce65;
        src73 <= 16'hb8c1;
        src74 <= 16'hd1fa;
        src75 <= 16'h602f;
        src76 <= 16'h2f8e;
        src77 <= 16'hd0f2;
        src78 <= 16'hadba;
        src79 <= 16'h5f05;
        src80 <= 16'h12a8;
        src81 <= 16'he67a;
        src82 <= 16'h9729;
        src83 <= 16'h388;
        src84 <= 16'h6379;
        src85 <= 16'had2e;
        src86 <= 16'hcfd2;
        src87 <= 16'h6e50;
        src88 <= 16'hd0ce;
        src89 <= 16'h2209;
        src90 <= 16'h7c;
        src91 <= 16'h8fb3;
        src92 <= 16'hb9d3;
        src93 <= 16'hd1d7;
        src94 <= 16'hdac6;
        src95 <= 16'hcfae;
        src96 <= 16'h2da3;
        src97 <= 16'hab6;
        src98 <= 16'h390c;
        src99 <= 16'h1911;
        src100 <= 16'h3612;
        src101 <= 16'hf880;
        src102 <= 16'h7781;
        src103 <= 16'hd3f5;
        src104 <= 16'hbcc3;
        src105 <= 16'hc6aa;
        src106 <= 16'h6af3;
        src107 <= 16'h4407;
        src108 <= 16'ha086;
        src109 <= 16'ha62e;
        src110 <= 16'hfb5c;
        src111 <= 16'h329e;
        src112 <= 16'h381f;
        src113 <= 16'h7412;
        src114 <= 16'h9467;
        src115 <= 16'h5b05;
        src116 <= 16'h2ae1;
        src117 <= 16'h82ed;
        src118 <= 16'hd81;
        src119 <= 16'he9f0;
        src120 <= 16'ha64c;
        src121 <= 16'h833b;
        src122 <= 16'ha7dd;
        src123 <= 16'haaab;
        src124 <= 16'h71d4;
        src125 <= 16'h544d;
        src126 <= 16'h37b7;
        src127 <= 16'h825d;
        src128 <= 16'h5c01;
        src129 <= 16'h3f66;
        src130 <= 16'ha5e2;
        src131 <= 16'hdec1;
        src132 <= 16'hf019;
        src133 <= 16'h9a4b;
        src134 <= 16'h8022;
        src135 <= 16'hf7ec;
        src136 <= 16'ha7c4;
        src137 <= 16'h4cc4;
        src138 <= 16'hcf5f;
        src139 <= 16'haa2f;
        src140 <= 16'hee76;
        src141 <= 16'h133a;
        src142 <= 16'hf6f2;
        src143 <= 16'h84f9;
        src144 <= 16'ha1b0;
        src145 <= 16'hdbd5;
        src146 <= 16'h29b6;
        src147 <= 16'h635f;
        src148 <= 16'hde1;
        src149 <= 16'h59f7;
        src150 <= 16'hd9d0;
        src151 <= 16'h7ccb;
        src152 <= 16'had4a;
        src153 <= 16'h739e;
        src154 <= 16'h9b43;
        src155 <= 16'hef2d;
        src156 <= 16'h4692;
        src157 <= 16'h977e;
        src158 <= 16'h8a23;
        src159 <= 16'h39d6;
        src160 <= 16'h6367;
        src161 <= 16'hb0be;
        src162 <= 16'h3b30;
        src163 <= 16'h24e5;
        src164 <= 16'hb206;
        src165 <= 16'h7f65;
        src166 <= 16'hffdf;
        src167 <= 16'h3c45;
        src168 <= 16'h78f5;
        src169 <= 16'headc;
        src170 <= 16'h16ef;
        src171 <= 16'hb786;
        src172 <= 16'hf8e6;
        src173 <= 16'h3887;
        src174 <= 16'h70e3;
        src175 <= 16'hd0b5;
        src176 <= 16'h37fe;
        src177 <= 16'h861d;
        src178 <= 16'h1e64;
        src179 <= 16'h34a0;
        src180 <= 16'h7941;
        src181 <= 16'h138;
        src182 <= 16'h4283;
        src183 <= 16'ha418;
        src184 <= 16'h51a2;
        exp <= 24'h603114;
        #1
        src0 <= 16'hb5db;
        src1 <= 16'h41ad;
        src2 <= 16'h3372;
        src3 <= 16'h2703;
        src4 <= 16'he187;
        src5 <= 16'h268;
        src6 <= 16'h4c6;
        src7 <= 16'h4d0e;
        src8 <= 16'hc172;
        src9 <= 16'hfd7b;
        src10 <= 16'hc86e;
        src11 <= 16'h2863;
        src12 <= 16'h86bb;
        src13 <= 16'h1360;
        src14 <= 16'h32ed;
        src15 <= 16'h8c41;
        src16 <= 16'h643d;
        src17 <= 16'h62df;
        src18 <= 16'h7de5;
        src19 <= 16'h17d3;
        src20 <= 16'hb047;
        src21 <= 16'hd1d;
        src22 <= 16'h697e;
        src23 <= 16'h8763;
        src24 <= 16'h5973;
        src25 <= 16'h3187;
        src26 <= 16'h9bf0;
        src27 <= 16'h8cc0;
        src28 <= 16'hb904;
        src29 <= 16'h4756;
        src30 <= 16'h4e7d;
        src31 <= 16'h6db6;
        src32 <= 16'h15b2;
        src33 <= 16'h83f;
        src34 <= 16'h5c8f;
        src35 <= 16'h49d8;
        src36 <= 16'h952d;
        src37 <= 16'h51d3;
        src38 <= 16'h3a99;
        src39 <= 16'h5b05;
        src40 <= 16'h90c2;
        src41 <= 16'hd1b;
        src42 <= 16'h9983;
        src43 <= 16'hf5ca;
        src44 <= 16'h7044;
        src45 <= 16'h633c;
        src46 <= 16'h5827;
        src47 <= 16'h2cb4;
        src48 <= 16'h5868;
        src49 <= 16'h5564;
        src50 <= 16'h6d44;
        src51 <= 16'h9d65;
        src52 <= 16'hdabe;
        src53 <= 16'hf5ea;
        src54 <= 16'h81d7;
        src55 <= 16'ha8b7;
        src56 <= 16'h413a;
        src57 <= 16'habc1;
        src58 <= 16'h2f80;
        src59 <= 16'hd978;
        src60 <= 16'h330c;
        src61 <= 16'h9c8d;
        src62 <= 16'h2dd7;
        src63 <= 16'hcaa5;
        src64 <= 16'h9357;
        src65 <= 16'h1b9;
        src66 <= 16'hba8c;
        src67 <= 16'hb87b;
        src68 <= 16'h3b01;
        src69 <= 16'h2e7e;
        src70 <= 16'hfa63;
        src71 <= 16'hb46c;
        src72 <= 16'hf86f;
        src73 <= 16'h67b7;
        src74 <= 16'hee13;
        src75 <= 16'h4faf;
        src76 <= 16'hf997;
        src77 <= 16'h45d6;
        src78 <= 16'hd113;
        src79 <= 16'h4d47;
        src80 <= 16'h1c73;
        src81 <= 16'hc702;
        src82 <= 16'h9e16;
        src83 <= 16'h236;
        src84 <= 16'hb1e0;
        src85 <= 16'h718a;
        src86 <= 16'hc898;
        src87 <= 16'h8797;
        src88 <= 16'h6043;
        src89 <= 16'hbc3a;
        src90 <= 16'h12a7;
        src91 <= 16'he152;
        src92 <= 16'ha2f3;
        src93 <= 16'h6f18;
        src94 <= 16'h9569;
        src95 <= 16'hcd98;
        src96 <= 16'habbd;
        src97 <= 16'hd3c8;
        src98 <= 16'hb3e6;
        src99 <= 16'hed5e;
        src100 <= 16'h572;
        src101 <= 16'hbe2b;
        src102 <= 16'h6901;
        src103 <= 16'h50fe;
        src104 <= 16'h49b0;
        src105 <= 16'h729f;
        src106 <= 16'h6a79;
        src107 <= 16'h36ef;
        src108 <= 16'hb833;
        src109 <= 16'he53e;
        src110 <= 16'hdbcf;
        src111 <= 16'h23c4;
        src112 <= 16'h540d;
        src113 <= 16'h9be;
        src114 <= 16'h2d08;
        src115 <= 16'hfa36;
        src116 <= 16'h99ec;
        src117 <= 16'hd21a;
        src118 <= 16'h407c;
        src119 <= 16'hfa26;
        src120 <= 16'h5585;
        src121 <= 16'hfd60;
        src122 <= 16'hf191;
        src123 <= 16'hcba9;
        src124 <= 16'h4664;
        src125 <= 16'he514;
        src126 <= 16'hbc48;
        src127 <= 16'h211d;
        src128 <= 16'hf42;
        src129 <= 16'hd964;
        src130 <= 16'h51bf;
        src131 <= 16'h9a72;
        src132 <= 16'hb08a;
        src133 <= 16'hd5b6;
        src134 <= 16'h8f51;
        src135 <= 16'h4d0c;
        src136 <= 16'h3247;
        src137 <= 16'hfac6;
        src138 <= 16'h5d5c;
        src139 <= 16'h57fd;
        src140 <= 16'h8f04;
        src141 <= 16'h6401;
        src142 <= 16'hf45e;
        src143 <= 16'he934;
        src144 <= 16'h8089;
        src145 <= 16'hf17a;
        src146 <= 16'hde99;
        src147 <= 16'ha5b;
        src148 <= 16'h183;
        src149 <= 16'h8ea1;
        src150 <= 16'hd22b;
        src151 <= 16'h768c;
        src152 <= 16'h5b1;
        src153 <= 16'h26a5;
        src154 <= 16'h4228;
        src155 <= 16'hd3ef;
        src156 <= 16'hbce4;
        src157 <= 16'hb15b;
        src158 <= 16'h46fe;
        src159 <= 16'hc5c4;
        src160 <= 16'h4f6a;
        src161 <= 16'h9b54;
        src162 <= 16'h5890;
        src163 <= 16'h4807;
        src164 <= 16'he266;
        src165 <= 16'h43cf;
        src166 <= 16'ha725;
        src167 <= 16'h334;
        src168 <= 16'hf969;
        src169 <= 16'h780f;
        src170 <= 16'h9a3b;
        src171 <= 16'h2de9;
        src172 <= 16'heba2;
        src173 <= 16'h58d6;
        src174 <= 16'h628;
        src175 <= 16'h2138;
        src176 <= 16'h452c;
        src177 <= 16'he2fe;
        src178 <= 16'he59a;
        src179 <= 16'h821d;
        src180 <= 16'h4898;
        src181 <= 16'h5892;
        src182 <= 16'hbda6;
        src183 <= 16'ha2ec;
        src184 <= 16'h17b;
        exp <= 24'h5b2b22;
        #1
        src0 <= 16'h7e48;
        src1 <= 16'hf5f3;
        src2 <= 16'h556a;
        src3 <= 16'h6093;
        src4 <= 16'h8bc8;
        src5 <= 16'hddec;
        src6 <= 16'ha5f8;
        src7 <= 16'hf41e;
        src8 <= 16'ha04d;
        src9 <= 16'h39d2;
        src10 <= 16'h365b;
        src11 <= 16'h10df;
        src12 <= 16'h419;
        src13 <= 16'h933;
        src14 <= 16'h8665;
        src15 <= 16'h7707;
        src16 <= 16'h5a;
        src17 <= 16'h96d;
        src18 <= 16'h4705;
        src19 <= 16'hcae2;
        src20 <= 16'hff68;
        src21 <= 16'hc608;
        src22 <= 16'hd29c;
        src23 <= 16'h9f59;
        src24 <= 16'hf3ec;
        src25 <= 16'h4ea4;
        src26 <= 16'h2415;
        src27 <= 16'hd63e;
        src28 <= 16'h5a71;
        src29 <= 16'h42d8;
        src30 <= 16'h8f4a;
        src31 <= 16'hf68d;
        src32 <= 16'hf37f;
        src33 <= 16'h103c;
        src34 <= 16'he8f1;
        src35 <= 16'h2897;
        src36 <= 16'h343e;
        src37 <= 16'hd38d;
        src38 <= 16'haad2;
        src39 <= 16'h9df8;
        src40 <= 16'hb5c;
        src41 <= 16'hf1c4;
        src42 <= 16'h7ef6;
        src43 <= 16'hf2a1;
        src44 <= 16'h91d;
        src45 <= 16'hde0;
        src46 <= 16'h46e4;
        src47 <= 16'hf7b9;
        src48 <= 16'h5031;
        src49 <= 16'h59f5;
        src50 <= 16'hd58c;
        src51 <= 16'h72f;
        src52 <= 16'hf087;
        src53 <= 16'hfffb;
        src54 <= 16'hda54;
        src55 <= 16'hd7ea;
        src56 <= 16'hb284;
        src57 <= 16'hb316;
        src58 <= 16'h3f3;
        src59 <= 16'h7b5b;
        src60 <= 16'hb954;
        src61 <= 16'h1a10;
        src62 <= 16'hfeeb;
        src63 <= 16'ha83a;
        src64 <= 16'h1e8a;
        src65 <= 16'h5ded;
        src66 <= 16'h6143;
        src67 <= 16'he446;
        src68 <= 16'h31b5;
        src69 <= 16'h3fb;
        src70 <= 16'h733a;
        src71 <= 16'h6d24;
        src72 <= 16'hdf8c;
        src73 <= 16'h7adf;
        src74 <= 16'h77a2;
        src75 <= 16'h3af3;
        src76 <= 16'hdfe0;
        src77 <= 16'h5f0f;
        src78 <= 16'h5023;
        src79 <= 16'h185;
        src80 <= 16'h6c24;
        src81 <= 16'h8cb0;
        src82 <= 16'h217b;
        src83 <= 16'hf8c;
        src84 <= 16'headc;
        src85 <= 16'hcd14;
        src86 <= 16'he75b;
        src87 <= 16'h6ef6;
        src88 <= 16'h9c48;
        src89 <= 16'h8e13;
        src90 <= 16'h7bfa;
        src91 <= 16'h1419;
        src92 <= 16'hc824;
        src93 <= 16'h7c09;
        src94 <= 16'h507e;
        src95 <= 16'he707;
        src96 <= 16'h3364;
        src97 <= 16'h8ab5;
        src98 <= 16'hdb7;
        src99 <= 16'h3d71;
        src100 <= 16'h2dfa;
        src101 <= 16'h94ef;
        src102 <= 16'hfa92;
        src103 <= 16'h2550;
        src104 <= 16'h264f;
        src105 <= 16'h3bed;
        src106 <= 16'hba18;
        src107 <= 16'hf955;
        src108 <= 16'h54f9;
        src109 <= 16'hc16;
        src110 <= 16'h1d20;
        src111 <= 16'h9785;
        src112 <= 16'h2a38;
        src113 <= 16'h7455;
        src114 <= 16'h18a2;
        src115 <= 16'h6fcc;
        src116 <= 16'h6f62;
        src117 <= 16'h121f;
        src118 <= 16'h968c;
        src119 <= 16'h3362;
        src120 <= 16'h9fd8;
        src121 <= 16'h8fa8;
        src122 <= 16'hff91;
        src123 <= 16'h8067;
        src124 <= 16'h1e75;
        src125 <= 16'h4671;
        src126 <= 16'h14c3;
        src127 <= 16'h42b0;
        src128 <= 16'h201d;
        src129 <= 16'h2803;
        src130 <= 16'h2ed3;
        src131 <= 16'h54de;
        src132 <= 16'h44a1;
        src133 <= 16'h65be;
        src134 <= 16'hceee;
        src135 <= 16'h55d4;
        src136 <= 16'h8f40;
        src137 <= 16'heaf0;
        src138 <= 16'h860c;
        src139 <= 16'hbbf2;
        src140 <= 16'hc4e0;
        src141 <= 16'ha1a0;
        src142 <= 16'hdd1b;
        src143 <= 16'h4c45;
        src144 <= 16'h782e;
        src145 <= 16'h377a;
        src146 <= 16'h8920;
        src147 <= 16'h98a;
        src148 <= 16'hff27;
        src149 <= 16'hb350;
        src150 <= 16'h1bdf;
        src151 <= 16'h183d;
        src152 <= 16'hc450;
        src153 <= 16'hbfe5;
        src154 <= 16'hfbd3;
        src155 <= 16'h942f;
        src156 <= 16'h79a;
        src157 <= 16'hcda0;
        src158 <= 16'h4684;
        src159 <= 16'h93f1;
        src160 <= 16'hd6dd;
        src161 <= 16'hc288;
        src162 <= 16'h558c;
        src163 <= 16'hbcf9;
        src164 <= 16'h8da;
        src165 <= 16'h89d4;
        src166 <= 16'h5a9e;
        src167 <= 16'h9010;
        src168 <= 16'h5c88;
        src169 <= 16'hb0c7;
        src170 <= 16'hdb5b;
        src171 <= 16'hcd9e;
        src172 <= 16'ha1dc;
        src173 <= 16'h65b9;
        src174 <= 16'h25f2;
        src175 <= 16'hc111;
        src176 <= 16'h7918;
        src177 <= 16'h5fab;
        src178 <= 16'hb8e6;
        src179 <= 16'ha260;
        src180 <= 16'h874e;
        src181 <= 16'hc951;
        src182 <= 16'h29b0;
        src183 <= 16'h302;
        src184 <= 16'h91d8;
        exp <= 24'h597f0c;
        #1
        src0 <= 16'h43c0;
        src1 <= 16'h97c3;
        src2 <= 16'h8ca1;
        src3 <= 16'h6cfe;
        src4 <= 16'h32a8;
        src5 <= 16'hf117;
        src6 <= 16'h36db;
        src7 <= 16'hd3c6;
        src8 <= 16'he26b;
        src9 <= 16'h3f54;
        src10 <= 16'h7358;
        src11 <= 16'hb998;
        src12 <= 16'h8116;
        src13 <= 16'haa00;
        src14 <= 16'hfec7;
        src15 <= 16'h86cf;
        src16 <= 16'h1555;
        src17 <= 16'h53a4;
        src18 <= 16'h2c7d;
        src19 <= 16'h6b90;
        src20 <= 16'heae7;
        src21 <= 16'h5602;
        src22 <= 16'h59be;
        src23 <= 16'h8e49;
        src24 <= 16'h8392;
        src25 <= 16'h353;
        src26 <= 16'hbe85;
        src27 <= 16'ha3b5;
        src28 <= 16'ha34f;
        src29 <= 16'h2a48;
        src30 <= 16'h85b9;
        src31 <= 16'h56fa;
        src32 <= 16'h2c;
        src33 <= 16'hba7;
        src34 <= 16'hab27;
        src35 <= 16'ha746;
        src36 <= 16'h2da7;
        src37 <= 16'h7dcc;
        src38 <= 16'h8120;
        src39 <= 16'h2bf6;
        src40 <= 16'h42ab;
        src41 <= 16'hc7ac;
        src42 <= 16'h66f5;
        src43 <= 16'h8ce3;
        src44 <= 16'h4320;
        src45 <= 16'hd370;
        src46 <= 16'h98f9;
        src47 <= 16'h7c6d;
        src48 <= 16'hd134;
        src49 <= 16'hc632;
        src50 <= 16'hf14c;
        src51 <= 16'hfde5;
        src52 <= 16'h2ce7;
        src53 <= 16'hb45;
        src54 <= 16'hf6b5;
        src55 <= 16'h7678;
        src56 <= 16'hddbb;
        src57 <= 16'hcaaa;
        src58 <= 16'hf31a;
        src59 <= 16'hb047;
        src60 <= 16'h137e;
        src61 <= 16'h2fcf;
        src62 <= 16'hb02e;
        src63 <= 16'hacb2;
        src64 <= 16'hceb9;
        src65 <= 16'h24c4;
        src66 <= 16'h4d9b;
        src67 <= 16'h6694;
        src68 <= 16'h1e8f;
        src69 <= 16'hc680;
        src70 <= 16'he18;
        src71 <= 16'hd800;
        src72 <= 16'h2f25;
        src73 <= 16'haf51;
        src74 <= 16'hbbe0;
        src75 <= 16'h8b80;
        src76 <= 16'hcd0d;
        src77 <= 16'h5e0e;
        src78 <= 16'he395;
        src79 <= 16'heccb;
        src80 <= 16'hfff4;
        src81 <= 16'hbaba;
        src82 <= 16'h5ff9;
        src83 <= 16'h42dc;
        src84 <= 16'hc97a;
        src85 <= 16'hed70;
        src86 <= 16'he949;
        src87 <= 16'h95da;
        src88 <= 16'h919;
        src89 <= 16'hcae;
        src90 <= 16'h1355;
        src91 <= 16'hdc1f;
        src92 <= 16'h93c7;
        src93 <= 16'h9116;
        src94 <= 16'h99aa;
        src95 <= 16'h873e;
        src96 <= 16'hed8a;
        src97 <= 16'ha55;
        src98 <= 16'hcf13;
        src99 <= 16'h25a;
        src100 <= 16'h67bf;
        src101 <= 16'h3692;
        src102 <= 16'h6b2b;
        src103 <= 16'h3659;
        src104 <= 16'hb149;
        src105 <= 16'heff8;
        src106 <= 16'h890a;
        src107 <= 16'h2e31;
        src108 <= 16'h79cb;
        src109 <= 16'he5dc;
        src110 <= 16'h5e98;
        src111 <= 16'h2f01;
        src112 <= 16'h3497;
        src113 <= 16'h2d66;
        src114 <= 16'h5a4a;
        src115 <= 16'h2438;
        src116 <= 16'he820;
        src117 <= 16'h210;
        src118 <= 16'h5892;
        src119 <= 16'h84fd;
        src120 <= 16'he7e;
        src121 <= 16'h39d3;
        src122 <= 16'hbb8e;
        src123 <= 16'hb71d;
        src124 <= 16'hfb36;
        src125 <= 16'hedf9;
        src126 <= 16'h5936;
        src127 <= 16'hd34a;
        src128 <= 16'ha463;
        src129 <= 16'hbc24;
        src130 <= 16'hb1cf;
        src131 <= 16'hb514;
        src132 <= 16'h7f55;
        src133 <= 16'h11c9;
        src134 <= 16'hd9d6;
        src135 <= 16'h7344;
        src136 <= 16'he453;
        src137 <= 16'hf755;
        src138 <= 16'h14cd;
        src139 <= 16'h46a6;
        src140 <= 16'h3384;
        src141 <= 16'ha6e2;
        src142 <= 16'hf52a;
        src143 <= 16'h9735;
        src144 <= 16'he722;
        src145 <= 16'h59a5;
        src146 <= 16'h5dbb;
        src147 <= 16'h53c4;
        src148 <= 16'ha8c0;
        src149 <= 16'h8210;
        src150 <= 16'h2710;
        src151 <= 16'he799;
        src152 <= 16'h5761;
        src153 <= 16'h78aa;
        src154 <= 16'h58bb;
        src155 <= 16'hb4de;
        src156 <= 16'h81f4;
        src157 <= 16'hde52;
        src158 <= 16'h2526;
        src159 <= 16'ha408;
        src160 <= 16'h22ec;
        src161 <= 16'hab22;
        src162 <= 16'hddb4;
        src163 <= 16'h5b75;
        src164 <= 16'h7541;
        src165 <= 16'h19d7;
        src166 <= 16'h851a;
        src167 <= 16'haf72;
        src168 <= 16'hf8f6;
        src169 <= 16'h2912;
        src170 <= 16'h815e;
        src171 <= 16'h7d97;
        src172 <= 16'hc503;
        src173 <= 16'h7491;
        src174 <= 16'h4a40;
        src175 <= 16'h1697;
        src176 <= 16'h199a;
        src177 <= 16'h3b4c;
        src178 <= 16'h5d15;
        src179 <= 16'h5cd3;
        src180 <= 16'had57;
        src181 <= 16'h4ff6;
        src182 <= 16'h92d9;
        src183 <= 16'h4488;
        src184 <= 16'h7e34;
        exp <= 24'h5d51d3;
        #1
        src0 <= 16'h1203;
        src1 <= 16'hd7bd;
        src2 <= 16'hcf5f;
        src3 <= 16'h4753;
        src4 <= 16'hf63d;
        src5 <= 16'haf6a;
        src6 <= 16'hf660;
        src7 <= 16'hed48;
        src8 <= 16'hf64e;
        src9 <= 16'hcb8a;
        src10 <= 16'h22a8;
        src11 <= 16'h4b93;
        src12 <= 16'h9ebd;
        src13 <= 16'hd1a3;
        src14 <= 16'h9c7f;
        src15 <= 16'hfc4;
        src16 <= 16'h828f;
        src17 <= 16'h887a;
        src18 <= 16'h704;
        src19 <= 16'ha627;
        src20 <= 16'h2799;
        src21 <= 16'h626e;
        src22 <= 16'h7f75;
        src23 <= 16'h1176;
        src24 <= 16'hbc5e;
        src25 <= 16'hc539;
        src26 <= 16'hb80b;
        src27 <= 16'hcc4a;
        src28 <= 16'h613d;
        src29 <= 16'hc152;
        src30 <= 16'h8284;
        src31 <= 16'h4ed4;
        src32 <= 16'h479a;
        src33 <= 16'h4c06;
        src34 <= 16'h6b25;
        src35 <= 16'hdb05;
        src36 <= 16'h2141;
        src37 <= 16'hceac;
        src38 <= 16'he5bd;
        src39 <= 16'hf85d;
        src40 <= 16'hed50;
        src41 <= 16'h84bf;
        src42 <= 16'h4da3;
        src43 <= 16'hc516;
        src44 <= 16'h5907;
        src45 <= 16'h32d7;
        src46 <= 16'h7c73;
        src47 <= 16'hf799;
        src48 <= 16'h32f5;
        src49 <= 16'h24ff;
        src50 <= 16'hba21;
        src51 <= 16'heb72;
        src52 <= 16'heb67;
        src53 <= 16'hd43a;
        src54 <= 16'h9eac;
        src55 <= 16'h2a4f;
        src56 <= 16'ha80a;
        src57 <= 16'h8e0;
        src58 <= 16'hb3c6;
        src59 <= 16'h585a;
        src60 <= 16'ha6e1;
        src61 <= 16'hff40;
        src62 <= 16'hf919;
        src63 <= 16'h599c;
        src64 <= 16'he375;
        src65 <= 16'h91a8;
        src66 <= 16'h5885;
        src67 <= 16'h2aaa;
        src68 <= 16'hac41;
        src69 <= 16'h783c;
        src70 <= 16'h613f;
        src71 <= 16'h77bf;
        src72 <= 16'h17c;
        src73 <= 16'he023;
        src74 <= 16'ha88a;
        src75 <= 16'h6dd6;
        src76 <= 16'hdd2d;
        src77 <= 16'hd955;
        src78 <= 16'h53d3;
        src79 <= 16'hf86;
        src80 <= 16'h1726;
        src81 <= 16'h434d;
        src82 <= 16'h60c4;
        src83 <= 16'h7b4f;
        src84 <= 16'h4e1c;
        src85 <= 16'h5b2d;
        src86 <= 16'h18f;
        src87 <= 16'hca;
        src88 <= 16'h84ad;
        src89 <= 16'he54d;
        src90 <= 16'h361f;
        src91 <= 16'hb79a;
        src92 <= 16'h1e30;
        src93 <= 16'h7335;
        src94 <= 16'ha994;
        src95 <= 16'h6eed;
        src96 <= 16'h46de;
        src97 <= 16'he501;
        src98 <= 16'ha8c1;
        src99 <= 16'h603;
        src100 <= 16'h4246;
        src101 <= 16'hf489;
        src102 <= 16'hcd9;
        src103 <= 16'hb776;
        src104 <= 16'h23ea;
        src105 <= 16'h5387;
        src106 <= 16'hd370;
        src107 <= 16'h481a;
        src108 <= 16'h7673;
        src109 <= 16'h1cec;
        src110 <= 16'h6db8;
        src111 <= 16'h5523;
        src112 <= 16'h1d0e;
        src113 <= 16'h8534;
        src114 <= 16'h1eab;
        src115 <= 16'h4b9d;
        src116 <= 16'he52f;
        src117 <= 16'h4ef8;
        src118 <= 16'hd335;
        src119 <= 16'h7fc9;
        src120 <= 16'h7b6f;
        src121 <= 16'h3180;
        src122 <= 16'h6172;
        src123 <= 16'h17ad;
        src124 <= 16'h2405;
        src125 <= 16'hf07e;
        src126 <= 16'h33c9;
        src127 <= 16'h85c2;
        src128 <= 16'h1b86;
        src129 <= 16'h245a;
        src130 <= 16'h5ed0;
        src131 <= 16'hb257;
        src132 <= 16'h2c40;
        src133 <= 16'h5be8;
        src134 <= 16'h47eb;
        src135 <= 16'h9a2a;
        src136 <= 16'h156e;
        src137 <= 16'hf5ec;
        src138 <= 16'h15ef;
        src139 <= 16'h3e1f;
        src140 <= 16'hd9c3;
        src141 <= 16'h14b3;
        src142 <= 16'h32fb;
        src143 <= 16'hc950;
        src144 <= 16'h94a5;
        src145 <= 16'h1088;
        src146 <= 16'h7c7d;
        src147 <= 16'h8b3f;
        src148 <= 16'h2094;
        src149 <= 16'hba17;
        src150 <= 16'h8ca8;
        src151 <= 16'hd71b;
        src152 <= 16'h1188;
        src153 <= 16'hc43f;
        src154 <= 16'h7797;
        src155 <= 16'hf50e;
        src156 <= 16'h1c97;
        src157 <= 16'h433;
        src158 <= 16'ha960;
        src159 <= 16'h8d85;
        src160 <= 16'h88d1;
        src161 <= 16'hf2fe;
        src162 <= 16'h342d;
        src163 <= 16'h6463;
        src164 <= 16'hc78f;
        src165 <= 16'h438;
        src166 <= 16'h6c6f;
        src167 <= 16'h6dcc;
        src168 <= 16'hf785;
        src169 <= 16'h5ccc;
        src170 <= 16'h5805;
        src171 <= 16'he533;
        src172 <= 16'h827e;
        src173 <= 16'h753b;
        src174 <= 16'h22f2;
        src175 <= 16'hc690;
        src176 <= 16'he8bd;
        src177 <= 16'h87f3;
        src178 <= 16'h768e;
        src179 <= 16'he0fd;
        src180 <= 16'h50d1;
        src181 <= 16'hd621;
        src182 <= 16'h5b19;
        src183 <= 16'h63f;
        src184 <= 16'h8f4d;
        exp <= 24'h59d5ef;
        #1
        src0 <= 16'h4d91;
        src1 <= 16'h1ac2;
        src2 <= 16'h7259;
        src3 <= 16'h27ea;
        src4 <= 16'hee65;
        src5 <= 16'h1baf;
        src6 <= 16'h561f;
        src7 <= 16'h7d30;
        src8 <= 16'he05f;
        src9 <= 16'h8fb1;
        src10 <= 16'h3658;
        src11 <= 16'h2ee7;
        src12 <= 16'hcbc3;
        src13 <= 16'hf0d2;
        src14 <= 16'ha277;
        src15 <= 16'h65e3;
        src16 <= 16'h8f0;
        src17 <= 16'h9e28;
        src18 <= 16'h5ce9;
        src19 <= 16'h4b36;
        src20 <= 16'h9111;
        src21 <= 16'h5c1c;
        src22 <= 16'hc9f9;
        src23 <= 16'hb978;
        src24 <= 16'h6ac7;
        src25 <= 16'h41d8;
        src26 <= 16'h51db;
        src27 <= 16'h2963;
        src28 <= 16'hd081;
        src29 <= 16'hccc1;
        src30 <= 16'hc79b;
        src31 <= 16'h3125;
        src32 <= 16'ha86e;
        src33 <= 16'h5cd3;
        src34 <= 16'he98b;
        src35 <= 16'h1c53;
        src36 <= 16'h576e;
        src37 <= 16'hba4a;
        src38 <= 16'h8db4;
        src39 <= 16'h3b70;
        src40 <= 16'h455d;
        src41 <= 16'hfcdc;
        src42 <= 16'h4294;
        src43 <= 16'hfc4e;
        src44 <= 16'ha677;
        src45 <= 16'h49f8;
        src46 <= 16'hf8f4;
        src47 <= 16'h1aa;
        src48 <= 16'hb640;
        src49 <= 16'h48a;
        src50 <= 16'ha4ae;
        src51 <= 16'hd0c7;
        src52 <= 16'hb56f;
        src53 <= 16'h857c;
        src54 <= 16'hb598;
        src55 <= 16'h644e;
        src56 <= 16'h210c;
        src57 <= 16'h880b;
        src58 <= 16'h6922;
        src59 <= 16'hf523;
        src60 <= 16'hee98;
        src61 <= 16'h27d5;
        src62 <= 16'h5f17;
        src63 <= 16'h3525;
        src64 <= 16'h1cfc;
        src65 <= 16'ha71c;
        src66 <= 16'h9db;
        src67 <= 16'hbff1;
        src68 <= 16'h61e5;
        src69 <= 16'h1ac3;
        src70 <= 16'h7331;
        src71 <= 16'h3481;
        src72 <= 16'he4ba;
        src73 <= 16'h16b5;
        src74 <= 16'hc1e3;
        src75 <= 16'h3f41;
        src76 <= 16'he410;
        src77 <= 16'h7c8;
        src78 <= 16'hc27a;
        src79 <= 16'h14a9;
        src80 <= 16'h34bb;
        src81 <= 16'h9d58;
        src82 <= 16'h63ad;
        src83 <= 16'h1fe;
        src84 <= 16'h6109;
        src85 <= 16'hba2;
        src86 <= 16'h5489;
        src87 <= 16'hf887;
        src88 <= 16'h5e7;
        src89 <= 16'h8fd6;
        src90 <= 16'he23b;
        src91 <= 16'hb4a9;
        src92 <= 16'h826e;
        src93 <= 16'h2dd9;
        src94 <= 16'h1a76;
        src95 <= 16'hfaf0;
        src96 <= 16'h3a95;
        src97 <= 16'h9170;
        src98 <= 16'h336f;
        src99 <= 16'h4967;
        src100 <= 16'he3e4;
        src101 <= 16'hfd76;
        src102 <= 16'h70ab;
        src103 <= 16'h2c3a;
        src104 <= 16'hc57a;
        src105 <= 16'h2591;
        src106 <= 16'ha6af;
        src107 <= 16'h3df1;
        src108 <= 16'h2e20;
        src109 <= 16'h8a90;
        src110 <= 16'hfb71;
        src111 <= 16'h659f;
        src112 <= 16'hc0d5;
        src113 <= 16'h21da;
        src114 <= 16'h50ac;
        src115 <= 16'h59ab;
        src116 <= 16'h1ea1;
        src117 <= 16'h2336;
        src118 <= 16'h23d0;
        src119 <= 16'hf2b;
        src120 <= 16'h18cc;
        src121 <= 16'he03d;
        src122 <= 16'hbf61;
        src123 <= 16'h127c;
        src124 <= 16'h92d7;
        src125 <= 16'hb224;
        src126 <= 16'hc7ab;
        src127 <= 16'hf7df;
        src128 <= 16'ha5b7;
        src129 <= 16'h62ed;
        src130 <= 16'h7002;
        src131 <= 16'h9f71;
        src132 <= 16'h1655;
        src133 <= 16'hace9;
        src134 <= 16'h18c;
        src135 <= 16'h492c;
        src136 <= 16'h76d;
        src137 <= 16'h208b;
        src138 <= 16'hc417;
        src139 <= 16'heeca;
        src140 <= 16'hbc8b;
        src141 <= 16'hac2c;
        src142 <= 16'hc7f6;
        src143 <= 16'h27b7;
        src144 <= 16'h8b94;
        src145 <= 16'ha648;
        src146 <= 16'hed81;
        src147 <= 16'hf9e4;
        src148 <= 16'h8106;
        src149 <= 16'hb0bc;
        src150 <= 16'he1e;
        src151 <= 16'h85cc;
        src152 <= 16'hba0a;
        src153 <= 16'h7d7e;
        src154 <= 16'hcfb8;
        src155 <= 16'h183;
        src156 <= 16'hf7f1;
        src157 <= 16'h7432;
        src158 <= 16'h45e;
        src159 <= 16'hcac6;
        src160 <= 16'hb1f0;
        src161 <= 16'h8c0;
        src162 <= 16'haf3a;
        src163 <= 16'hb861;
        src164 <= 16'hd427;
        src165 <= 16'h62b4;
        src166 <= 16'h7c57;
        src167 <= 16'h5ed1;
        src168 <= 16'h1135;
        src169 <= 16'h7e77;
        src170 <= 16'h4f2c;
        src171 <= 16'h26d9;
        src172 <= 16'hb0e0;
        src173 <= 16'haa6b;
        src174 <= 16'hfebe;
        src175 <= 16'hd267;
        src176 <= 16'hfa2e;
        src177 <= 16'h6874;
        src178 <= 16'h91a1;
        src179 <= 16'he354;
        src180 <= 16'hb2f7;
        src181 <= 16'hcbcf;
        src182 <= 16'h4da8;
        src183 <= 16'h559e;
        src184 <= 16'h59b;
        exp <= 24'h593a6c;
        #1
        src0 <= 16'hadd;
        src1 <= 16'he542;
        src2 <= 16'h3a08;
        src3 <= 16'he5c6;
        src4 <= 16'hc662;
        src5 <= 16'h401f;
        src6 <= 16'hfccb;
        src7 <= 16'h16ff;
        src8 <= 16'he20f;
        src9 <= 16'h3147;
        src10 <= 16'ha9c2;
        src11 <= 16'hc04f;
        src12 <= 16'hc11b;
        src13 <= 16'h44e1;
        src14 <= 16'h7e17;
        src15 <= 16'h45ab;
        src16 <= 16'he3ab;
        src17 <= 16'h118d;
        src18 <= 16'h94e;
        src19 <= 16'h9dea;
        src20 <= 16'ha627;
        src21 <= 16'h6bde;
        src22 <= 16'h7f1e;
        src23 <= 16'h95b;
        src24 <= 16'h71fa;
        src25 <= 16'h3582;
        src26 <= 16'hbe14;
        src27 <= 16'h5fd0;
        src28 <= 16'hc66a;
        src29 <= 16'h5d40;
        src30 <= 16'hea22;
        src31 <= 16'h5f0c;
        src32 <= 16'h3e49;
        src33 <= 16'hb04f;
        src34 <= 16'h2e50;
        src35 <= 16'hcddc;
        src36 <= 16'h9ecf;
        src37 <= 16'h710d;
        src38 <= 16'hcd6;
        src39 <= 16'h552e;
        src40 <= 16'ha115;
        src41 <= 16'h8215;
        src42 <= 16'h547f;
        src43 <= 16'h82b2;
        src44 <= 16'ha497;
        src45 <= 16'h17d1;
        src46 <= 16'h1534;
        src47 <= 16'h7f2a;
        src48 <= 16'h6728;
        src49 <= 16'h5e1d;
        src50 <= 16'h5473;
        src51 <= 16'ha43e;
        src52 <= 16'hb436;
        src53 <= 16'h6d50;
        src54 <= 16'h3f1e;
        src55 <= 16'hfcc7;
        src56 <= 16'hc599;
        src57 <= 16'h5db9;
        src58 <= 16'h686b;
        src59 <= 16'h1b42;
        src60 <= 16'hc49d;
        src61 <= 16'h71bf;
        src62 <= 16'h8709;
        src63 <= 16'he1db;
        src64 <= 16'h7391;
        src65 <= 16'h960f;
        src66 <= 16'h2e2a;
        src67 <= 16'h57f1;
        src68 <= 16'h227a;
        src69 <= 16'he6a9;
        src70 <= 16'h9460;
        src71 <= 16'hd7eb;
        src72 <= 16'h7eb6;
        src73 <= 16'ha58a;
        src74 <= 16'hdf8;
        src75 <= 16'h5580;
        src76 <= 16'hfeb6;
        src77 <= 16'h9fa4;
        src78 <= 16'hf72e;
        src79 <= 16'hf92c;
        src80 <= 16'h808f;
        src81 <= 16'hab67;
        src82 <= 16'h81dc;
        src83 <= 16'h2e11;
        src84 <= 16'hb0e6;
        src85 <= 16'h2446;
        src86 <= 16'h4837;
        src87 <= 16'hec43;
        src88 <= 16'ha460;
        src89 <= 16'hced;
        src90 <= 16'h9485;
        src91 <= 16'he574;
        src92 <= 16'h8fe4;
        src93 <= 16'hfb;
        src94 <= 16'hf7a7;
        src95 <= 16'h56c6;
        src96 <= 16'h3a07;
        src97 <= 16'hcc3c;
        src98 <= 16'h21ff;
        src99 <= 16'hb84c;
        src100 <= 16'hd89c;
        src101 <= 16'h709e;
        src102 <= 16'h816e;
        src103 <= 16'h75e7;
        src104 <= 16'h1c7b;
        src105 <= 16'hb7f3;
        src106 <= 16'hc0a3;
        src107 <= 16'h7cfe;
        src108 <= 16'h7454;
        src109 <= 16'h8ed2;
        src110 <= 16'he186;
        src111 <= 16'hfaef;
        src112 <= 16'hc6fa;
        src113 <= 16'hf43d;
        src114 <= 16'h4929;
        src115 <= 16'h806d;
        src116 <= 16'h8fd0;
        src117 <= 16'h160b;
        src118 <= 16'he7d0;
        src119 <= 16'h5dd8;
        src120 <= 16'hec0e;
        src121 <= 16'he8cf;
        src122 <= 16'h757e;
        src123 <= 16'h4713;
        src124 <= 16'h500e;
        src125 <= 16'h3c1;
        src126 <= 16'h907d;
        src127 <= 16'h29bc;
        src128 <= 16'hf115;
        src129 <= 16'hea78;
        src130 <= 16'hc73b;
        src131 <= 16'h1bfd;
        src132 <= 16'h1041;
        src133 <= 16'hf1b8;
        src134 <= 16'h4ff6;
        src135 <= 16'h5b0f;
        src136 <= 16'hce63;
        src137 <= 16'h4ca5;
        src138 <= 16'h58cd;
        src139 <= 16'hb34f;
        src140 <= 16'h5e24;
        src141 <= 16'hbcf;
        src142 <= 16'h484b;
        src143 <= 16'h9e3;
        src144 <= 16'h27cf;
        src145 <= 16'h334c;
        src146 <= 16'hc63b;
        src147 <= 16'h765b;
        src148 <= 16'hf663;
        src149 <= 16'h8ed1;
        src150 <= 16'hf13b;
        src151 <= 16'h1a6e;
        src152 <= 16'hca03;
        src153 <= 16'he0a1;
        src154 <= 16'h40cd;
        src155 <= 16'ha445;
        src156 <= 16'h7ad;
        src157 <= 16'h90fb;
        src158 <= 16'hbd53;
        src159 <= 16'hae67;
        src160 <= 16'hd94;
        src161 <= 16'h2ad4;
        src162 <= 16'hb3c5;
        src163 <= 16'h8fa4;
        src164 <= 16'h4da4;
        src165 <= 16'hfb00;
        src166 <= 16'h4876;
        src167 <= 16'hf5f3;
        src168 <= 16'hc48c;
        src169 <= 16'h3d30;
        src170 <= 16'h2db8;
        src171 <= 16'h5745;
        src172 <= 16'ha397;
        src173 <= 16'h8a98;
        src174 <= 16'h6e73;
        src175 <= 16'hb821;
        src176 <= 16'h79b3;
        src177 <= 16'ha4f3;
        src178 <= 16'h8db9;
        src179 <= 16'h8f6e;
        src180 <= 16'h502f;
        src181 <= 16'h5d1a;
        src182 <= 16'h7f32;
        src183 <= 16'h3b42;
        src184 <= 16'h36bd;
        exp <= 24'h5cd674;
        #1
        src0 <= 16'hd632;
        src1 <= 16'h8efe;
        src2 <= 16'ha4db;
        src3 <= 16'h5884;
        src4 <= 16'h5d22;
        src5 <= 16'h7cd8;
        src6 <= 16'hb656;
        src7 <= 16'h834e;
        src8 <= 16'h672e;
        src9 <= 16'he596;
        src10 <= 16'hd558;
        src11 <= 16'ha7d2;
        src12 <= 16'h58c7;
        src13 <= 16'h51c1;
        src14 <= 16'h2974;
        src15 <= 16'h8fc;
        src16 <= 16'h669d;
        src17 <= 16'habb9;
        src18 <= 16'h8333;
        src19 <= 16'hb5db;
        src20 <= 16'h51bb;
        src21 <= 16'hb3e9;
        src22 <= 16'h537c;
        src23 <= 16'hedcf;
        src24 <= 16'h335c;
        src25 <= 16'h3295;
        src26 <= 16'h76e7;
        src27 <= 16'haeb;
        src28 <= 16'hcc45;
        src29 <= 16'h56d2;
        src30 <= 16'h3f76;
        src31 <= 16'hc43;
        src32 <= 16'h7620;
        src33 <= 16'h9722;
        src34 <= 16'hb479;
        src35 <= 16'h5d6d;
        src36 <= 16'h56f9;
        src37 <= 16'h1731;
        src38 <= 16'h8e20;
        src39 <= 16'hee88;
        src40 <= 16'hc8a7;
        src41 <= 16'hee76;
        src42 <= 16'haaf5;
        src43 <= 16'ha9b8;
        src44 <= 16'h7e31;
        src45 <= 16'h7ee;
        src46 <= 16'h85c0;
        src47 <= 16'h2233;
        src48 <= 16'h8deb;
        src49 <= 16'hdea7;
        src50 <= 16'h8608;
        src51 <= 16'hbf46;
        src52 <= 16'hd0ff;
        src53 <= 16'hefe6;
        src54 <= 16'h80c9;
        src55 <= 16'hacf2;
        src56 <= 16'ha512;
        src57 <= 16'h459b;
        src58 <= 16'hb15;
        src59 <= 16'he222;
        src60 <= 16'h6866;
        src61 <= 16'h9e75;
        src62 <= 16'h274c;
        src63 <= 16'h115d;
        src64 <= 16'h2679;
        src65 <= 16'hec55;
        src66 <= 16'habf3;
        src67 <= 16'hc473;
        src68 <= 16'h8130;
        src69 <= 16'h1e47;
        src70 <= 16'h9e51;
        src71 <= 16'h40e3;
        src72 <= 16'hcd0e;
        src73 <= 16'hc05c;
        src74 <= 16'h48e9;
        src75 <= 16'h524e;
        src76 <= 16'he3e1;
        src77 <= 16'hf854;
        src78 <= 16'hd60b;
        src79 <= 16'hcc41;
        src80 <= 16'hdbf1;
        src81 <= 16'hb0f8;
        src82 <= 16'h8f89;
        src83 <= 16'he898;
        src84 <= 16'h4523;
        src85 <= 16'h74c9;
        src86 <= 16'h44b5;
        src87 <= 16'h308d;
        src88 <= 16'h2cb3;
        src89 <= 16'hc633;
        src90 <= 16'h6c5e;
        src91 <= 16'h2830;
        src92 <= 16'h7ae4;
        src93 <= 16'h1f86;
        src94 <= 16'hc277;
        src95 <= 16'h18ee;
        src96 <= 16'h45b5;
        src97 <= 16'h61ad;
        src98 <= 16'hc224;
        src99 <= 16'h8325;
        src100 <= 16'he011;
        src101 <= 16'hf2a8;
        src102 <= 16'h2f9;
        src103 <= 16'h3bab;
        src104 <= 16'hb15a;
        src105 <= 16'h2ac7;
        src106 <= 16'hcebc;
        src107 <= 16'ha88d;
        src108 <= 16'h6b00;
        src109 <= 16'h8c4;
        src110 <= 16'h1cb;
        src111 <= 16'hef2a;
        src112 <= 16'h9b3e;
        src113 <= 16'h8b1a;
        src114 <= 16'h54ed;
        src115 <= 16'h138e;
        src116 <= 16'h97f5;
        src117 <= 16'h7d28;
        src118 <= 16'h5215;
        src119 <= 16'hedb6;
        src120 <= 16'hb753;
        src121 <= 16'h6a96;
        src122 <= 16'hc240;
        src123 <= 16'hb50c;
        src124 <= 16'h9265;
        src125 <= 16'h2f25;
        src126 <= 16'h6d61;
        src127 <= 16'h7682;
        src128 <= 16'h8ca5;
        src129 <= 16'haa66;
        src130 <= 16'he29b;
        src131 <= 16'hd64d;
        src132 <= 16'h24fe;
        src133 <= 16'hba27;
        src134 <= 16'h14ff;
        src135 <= 16'h2ebf;
        src136 <= 16'h3d39;
        src137 <= 16'h8b6e;
        src138 <= 16'hf538;
        src139 <= 16'h1505;
        src140 <= 16'hc71e;
        src141 <= 16'had87;
        src142 <= 16'h74a1;
        src143 <= 16'h2899;
        src144 <= 16'hc87b;
        src145 <= 16'ha2b0;
        src146 <= 16'h9160;
        src147 <= 16'h3f2;
        src148 <= 16'ha28c;
        src149 <= 16'h1898;
        src150 <= 16'h2c5b;
        src151 <= 16'h1bfc;
        src152 <= 16'hb675;
        src153 <= 16'h519f;
        src154 <= 16'hc6f6;
        src155 <= 16'h443d;
        src156 <= 16'h5ac4;
        src157 <= 16'haf77;
        src158 <= 16'hdb2d;
        src159 <= 16'h5cfa;
        src160 <= 16'h10;
        src161 <= 16'h9ea2;
        src162 <= 16'hf1fa;
        src163 <= 16'hf3db;
        src164 <= 16'h9740;
        src165 <= 16'hf52;
        src166 <= 16'ha0ff;
        src167 <= 16'hf411;
        src168 <= 16'hc460;
        src169 <= 16'h202b;
        src170 <= 16'hef85;
        src171 <= 16'hcc9d;
        src172 <= 16'h7f8a;
        src173 <= 16'h2c93;
        src174 <= 16'h807b;
        src175 <= 16'hd78f;
        src176 <= 16'h9783;
        src177 <= 16'h29cf;
        src178 <= 16'h617c;
        src179 <= 16'hb891;
        src180 <= 16'h389;
        src181 <= 16'h7f72;
        src182 <= 16'h4957;
        src183 <= 16'h1fa5;
        src184 <= 16'h33b6;
        exp <= 24'h5c65fe;
        #1
        src0 <= 16'h85ff;
        src1 <= 16'hdf1;
        src2 <= 16'h8dd1;
        src3 <= 16'hf6f4;
        src4 <= 16'ha790;
        src5 <= 16'h946;
        src6 <= 16'h9099;
        src7 <= 16'haad;
        src8 <= 16'hb25e;
        src9 <= 16'h61d9;
        src10 <= 16'hc662;
        src11 <= 16'hd711;
        src12 <= 16'hb7dc;
        src13 <= 16'hfeec;
        src14 <= 16'hcf10;
        src15 <= 16'h4c8f;
        src16 <= 16'h735;
        src17 <= 16'h8bb6;
        src18 <= 16'h1d39;
        src19 <= 16'hb59;
        src20 <= 16'had7a;
        src21 <= 16'h285f;
        src22 <= 16'h83e2;
        src23 <= 16'h4db5;
        src24 <= 16'h88b8;
        src25 <= 16'h88bc;
        src26 <= 16'h734c;
        src27 <= 16'h7b75;
        src28 <= 16'h8141;
        src29 <= 16'h789a;
        src30 <= 16'hdd70;
        src31 <= 16'h19fe;
        src32 <= 16'h35b1;
        src33 <= 16'h35be;
        src34 <= 16'hfc07;
        src35 <= 16'h89aa;
        src36 <= 16'hae2;
        src37 <= 16'hd8c;
        src38 <= 16'h589f;
        src39 <= 16'hbfe5;
        src40 <= 16'hd36f;
        src41 <= 16'h5958;
        src42 <= 16'h90c5;
        src43 <= 16'h4c0a;
        src44 <= 16'h6cea;
        src45 <= 16'h9d54;
        src46 <= 16'h2983;
        src47 <= 16'h5c46;
        src48 <= 16'h1d54;
        src49 <= 16'h1582;
        src50 <= 16'he962;
        src51 <= 16'h5d5;
        src52 <= 16'h2176;
        src53 <= 16'h43ac;
        src54 <= 16'he7bc;
        src55 <= 16'h3dd6;
        src56 <= 16'hcc6d;
        src57 <= 16'h32fe;
        src58 <= 16'hba9e;
        src59 <= 16'he431;
        src60 <= 16'h3f30;
        src61 <= 16'hd39b;
        src62 <= 16'h7f2c;
        src63 <= 16'hb038;
        src64 <= 16'h8af8;
        src65 <= 16'h86e1;
        src66 <= 16'hd951;
        src67 <= 16'ha854;
        src68 <= 16'hc397;
        src69 <= 16'h746d;
        src70 <= 16'ha6a6;
        src71 <= 16'h7498;
        src72 <= 16'he3c0;
        src73 <= 16'hf702;
        src74 <= 16'h48c4;
        src75 <= 16'h4fe1;
        src76 <= 16'hda45;
        src77 <= 16'h9aec;
        src78 <= 16'h2987;
        src79 <= 16'he128;
        src80 <= 16'h989f;
        src81 <= 16'hbf95;
        src82 <= 16'h766;
        src83 <= 16'h16e0;
        src84 <= 16'hbdab;
        src85 <= 16'h517f;
        src86 <= 16'h1208;
        src87 <= 16'h7770;
        src88 <= 16'ha098;
        src89 <= 16'h4003;
        src90 <= 16'h71a5;
        src91 <= 16'hcffc;
        src92 <= 16'h2167;
        src93 <= 16'h2974;
        src94 <= 16'hb6df;
        src95 <= 16'h436b;
        src96 <= 16'hdb06;
        src97 <= 16'h1c3f;
        src98 <= 16'hbef3;
        src99 <= 16'h1afd;
        src100 <= 16'hf9de;
        src101 <= 16'ha3bf;
        src102 <= 16'hda7a;
        src103 <= 16'h2052;
        src104 <= 16'h5de;
        src105 <= 16'h6dae;
        src106 <= 16'h832e;
        src107 <= 16'h8e54;
        src108 <= 16'h2179;
        src109 <= 16'h5757;
        src110 <= 16'he16b;
        src111 <= 16'h8a16;
        src112 <= 16'heec0;
        src113 <= 16'ha70;
        src114 <= 16'h50a8;
        src115 <= 16'he1a5;
        src116 <= 16'hb7b1;
        src117 <= 16'h3b54;
        src118 <= 16'ha996;
        src119 <= 16'h645c;
        src120 <= 16'h3e9b;
        src121 <= 16'hc5;
        src122 <= 16'h4171;
        src123 <= 16'h3802;
        src124 <= 16'h622f;
        src125 <= 16'hdbc5;
        src126 <= 16'hd429;
        src127 <= 16'hdba8;
        src128 <= 16'h2f3a;
        src129 <= 16'h8080;
        src130 <= 16'h3a14;
        src131 <= 16'he5ae;
        src132 <= 16'h5fc6;
        src133 <= 16'hba75;
        src134 <= 16'h74;
        src135 <= 16'hf358;
        src136 <= 16'h1c7b;
        src137 <= 16'hbd1f;
        src138 <= 16'hba5c;
        src139 <= 16'hb38c;
        src140 <= 16'ha2b8;
        src141 <= 16'h835a;
        src142 <= 16'h9227;
        src143 <= 16'h812a;
        src144 <= 16'hcc51;
        src145 <= 16'ha128;
        src146 <= 16'h3e7f;
        src147 <= 16'hb3a7;
        src148 <= 16'h47d3;
        src149 <= 16'h204d;
        src150 <= 16'h7328;
        src151 <= 16'h6d42;
        src152 <= 16'ha5f6;
        src153 <= 16'ha310;
        src154 <= 16'h2c2f;
        src155 <= 16'hd6d2;
        src156 <= 16'h77df;
        src157 <= 16'h4ad0;
        src158 <= 16'h39d0;
        src159 <= 16'h5647;
        src160 <= 16'hbb10;
        src161 <= 16'h9aa1;
        src162 <= 16'h4cc9;
        src163 <= 16'h9a51;
        src164 <= 16'h4c9b;
        src165 <= 16'h15ad;
        src166 <= 16'ha02e;
        src167 <= 16'he9bc;
        src168 <= 16'hebbc;
        src169 <= 16'hc489;
        src170 <= 16'hfd2c;
        src171 <= 16'h4eab;
        src172 <= 16'hbff4;
        src173 <= 16'h3c7a;
        src174 <= 16'hacfa;
        src175 <= 16'hd27d;
        src176 <= 16'h6cf2;
        src177 <= 16'hf914;
        src178 <= 16'hc678;
        src179 <= 16'hff53;
        src180 <= 16'h60fa;
        src181 <= 16'h8793;
        src182 <= 16'h22d5;
        src183 <= 16'hdbe7;
        src184 <= 16'hf675;
        exp <= 24'h5ccc9e;
        #1
        src0 <= 16'hddfd;
        src1 <= 16'h51db;
        src2 <= 16'hef38;
        src3 <= 16'hb0e;
        src4 <= 16'haeaf;
        src5 <= 16'hc92d;
        src6 <= 16'hcc54;
        src7 <= 16'h4a77;
        src8 <= 16'h1e7f;
        src9 <= 16'h968;
        src10 <= 16'hc6a5;
        src11 <= 16'hb47;
        src12 <= 16'h65d8;
        src13 <= 16'h83cb;
        src14 <= 16'h31a;
        src15 <= 16'h4895;
        src16 <= 16'hcf0e;
        src17 <= 16'h9ed1;
        src18 <= 16'h6d28;
        src19 <= 16'h32e6;
        src20 <= 16'h8616;
        src21 <= 16'h1c13;
        src22 <= 16'heab8;
        src23 <= 16'h6670;
        src24 <= 16'h3a23;
        src25 <= 16'h6f37;
        src26 <= 16'hdfa5;
        src27 <= 16'h7582;
        src28 <= 16'h3615;
        src29 <= 16'hee4e;
        src30 <= 16'h280c;
        src31 <= 16'ha38b;
        src32 <= 16'h8fb;
        src33 <= 16'h23b9;
        src34 <= 16'hc75c;
        src35 <= 16'h1387;
        src36 <= 16'h66c4;
        src37 <= 16'h26de;
        src38 <= 16'hed0d;
        src39 <= 16'he297;
        src40 <= 16'hca0b;
        src41 <= 16'hb1a8;
        src42 <= 16'he172;
        src43 <= 16'hd735;
        src44 <= 16'h686c;
        src45 <= 16'h8bbb;
        src46 <= 16'haf5f;
        src47 <= 16'hf0d8;
        src48 <= 16'h4f74;
        src49 <= 16'h7547;
        src50 <= 16'h1ffb;
        src51 <= 16'h3edd;
        src52 <= 16'hb7c2;
        src53 <= 16'h99b1;
        src54 <= 16'h5d34;
        src55 <= 16'he08e;
        src56 <= 16'hfe29;
        src57 <= 16'hf0c0;
        src58 <= 16'ha350;
        src59 <= 16'h9e9c;
        src60 <= 16'h2279;
        src61 <= 16'had6f;
        src62 <= 16'h8718;
        src63 <= 16'h11f2;
        src64 <= 16'hce75;
        src65 <= 16'h5277;
        src66 <= 16'hcfb0;
        src67 <= 16'h328b;
        src68 <= 16'hb4c3;
        src69 <= 16'h956c;
        src70 <= 16'h976b;
        src71 <= 16'hfaf0;
        src72 <= 16'hcc6f;
        src73 <= 16'h3765;
        src74 <= 16'h380d;
        src75 <= 16'h56ff;
        src76 <= 16'ha23d;
        src77 <= 16'h8426;
        src78 <= 16'hbd85;
        src79 <= 16'hb4d2;
        src80 <= 16'h9e79;
        src81 <= 16'hc004;
        src82 <= 16'h37d0;
        src83 <= 16'h934b;
        src84 <= 16'h95b1;
        src85 <= 16'hc405;
        src86 <= 16'hebc5;
        src87 <= 16'habc0;
        src88 <= 16'haedd;
        src89 <= 16'h6374;
        src90 <= 16'h7ee1;
        src91 <= 16'h6b9b;
        src92 <= 16'hfa63;
        src93 <= 16'h673e;
        src94 <= 16'h1192;
        src95 <= 16'hacbd;
        src96 <= 16'hafbf;
        src97 <= 16'h42dd;
        src98 <= 16'h6e4a;
        src99 <= 16'h97c4;
        src100 <= 16'ha009;
        src101 <= 16'hf413;
        src102 <= 16'h8f6d;
        src103 <= 16'h7522;
        src104 <= 16'h185c;
        src105 <= 16'h4a84;
        src106 <= 16'hc59b;
        src107 <= 16'ha408;
        src108 <= 16'he2e6;
        src109 <= 16'h2df3;
        src110 <= 16'h2158;
        src111 <= 16'h3314;
        src112 <= 16'h87f5;
        src113 <= 16'h4c42;
        src114 <= 16'h8d4e;
        src115 <= 16'h7d94;
        src116 <= 16'h4f9f;
        src117 <= 16'hfb0c;
        src118 <= 16'hb839;
        src119 <= 16'h762f;
        src120 <= 16'hba0e;
        src121 <= 16'h1b99;
        src122 <= 16'hbfa2;
        src123 <= 16'he340;
        src124 <= 16'h8290;
        src125 <= 16'haf2;
        src126 <= 16'he349;
        src127 <= 16'hfc5;
        src128 <= 16'h8207;
        src129 <= 16'haeda;
        src130 <= 16'h2dd6;
        src131 <= 16'h48b8;
        src132 <= 16'h947c;
        src133 <= 16'hefdd;
        src134 <= 16'he0e6;
        src135 <= 16'h6bb;
        src136 <= 16'hbfbe;
        src137 <= 16'h7be3;
        src138 <= 16'h1e72;
        src139 <= 16'hab5d;
        src140 <= 16'hfc78;
        src141 <= 16'hcfee;
        src142 <= 16'h2cf6;
        src143 <= 16'hd146;
        src144 <= 16'h54fd;
        src145 <= 16'h4374;
        src146 <= 16'hfe0d;
        src147 <= 16'h8eb6;
        src148 <= 16'h91db;
        src149 <= 16'hf1d8;
        src150 <= 16'hce3;
        src151 <= 16'h581c;
        src152 <= 16'hfad;
        src153 <= 16'he24f;
        src154 <= 16'hbfcd;
        src155 <= 16'haa01;
        src156 <= 16'h93b7;
        src157 <= 16'h714d;
        src158 <= 16'h368;
        src159 <= 16'hf656;
        src160 <= 16'h4521;
        src161 <= 16'hd19a;
        src162 <= 16'h9bb2;
        src163 <= 16'h707f;
        src164 <= 16'hb231;
        src165 <= 16'hfe85;
        src166 <= 16'h2b86;
        src167 <= 16'h96d0;
        src168 <= 16'hd889;
        src169 <= 16'h387b;
        src170 <= 16'h532e;
        src171 <= 16'hb81b;
        src172 <= 16'h45e8;
        src173 <= 16'hd5b9;
        src174 <= 16'h15cb;
        src175 <= 16'hf805;
        src176 <= 16'h8bd1;
        src177 <= 16'h7ed5;
        src178 <= 16'h67b9;
        src179 <= 16'h5b85;
        src180 <= 16'h52f8;
        src181 <= 16'h139;
        src182 <= 16'h4328;
        src183 <= 16'hb705;
        src184 <= 16'h43ba;
        exp <= 24'h6050a3;
        #1
        src0 <= 16'hb79f;
        src1 <= 16'h66c0;
        src2 <= 16'h5868;
        src3 <= 16'he75d;
        src4 <= 16'h1963;
        src5 <= 16'h455a;
        src6 <= 16'h227e;
        src7 <= 16'hcb54;
        src8 <= 16'h3302;
        src9 <= 16'hf4d2;
        src10 <= 16'h5b12;
        src11 <= 16'h5f6a;
        src12 <= 16'h199d;
        src13 <= 16'hac26;
        src14 <= 16'h2269;
        src15 <= 16'hd73e;
        src16 <= 16'h90c8;
        src17 <= 16'hab68;
        src18 <= 16'h3279;
        src19 <= 16'h6cbf;
        src20 <= 16'h2e63;
        src21 <= 16'h4870;
        src22 <= 16'h4b24;
        src23 <= 16'hde1c;
        src24 <= 16'he864;
        src25 <= 16'ha647;
        src26 <= 16'hbc85;
        src27 <= 16'h69c0;
        src28 <= 16'h820b;
        src29 <= 16'h6dd2;
        src30 <= 16'hcf8b;
        src31 <= 16'h1cb0;
        src32 <= 16'h6804;
        src33 <= 16'h3025;
        src34 <= 16'hc9bd;
        src35 <= 16'h3a0;
        src36 <= 16'h4658;
        src37 <= 16'h19b1;
        src38 <= 16'h6e3a;
        src39 <= 16'h9abb;
        src40 <= 16'h563e;
        src41 <= 16'h4e7a;
        src42 <= 16'h189c;
        src43 <= 16'h9320;
        src44 <= 16'h74e5;
        src45 <= 16'h5760;
        src46 <= 16'hf5d4;
        src47 <= 16'h2441;
        src48 <= 16'h5753;
        src49 <= 16'h3a0c;
        src50 <= 16'h7182;
        src51 <= 16'h6d91;
        src52 <= 16'h1a2b;
        src53 <= 16'hf5cd;
        src54 <= 16'haf29;
        src55 <= 16'h7089;
        src56 <= 16'h7f8;
        src57 <= 16'hd4f;
        src58 <= 16'h749a;
        src59 <= 16'h4f8;
        src60 <= 16'hc4b2;
        src61 <= 16'h8eff;
        src62 <= 16'h7569;
        src63 <= 16'h6da5;
        src64 <= 16'h8252;
        src65 <= 16'hb625;
        src66 <= 16'h4627;
        src67 <= 16'hc384;
        src68 <= 16'h661c;
        src69 <= 16'h7502;
        src70 <= 16'had66;
        src71 <= 16'hb32c;
        src72 <= 16'hf65d;
        src73 <= 16'h312d;
        src74 <= 16'h5be7;
        src75 <= 16'hd914;
        src76 <= 16'hea22;
        src77 <= 16'h73cd;
        src78 <= 16'he950;
        src79 <= 16'h3565;
        src80 <= 16'ha617;
        src81 <= 16'hb9de;
        src82 <= 16'h67a4;
        src83 <= 16'hc19c;
        src84 <= 16'h10db;
        src85 <= 16'h7c03;
        src86 <= 16'ha6c3;
        src87 <= 16'h20e5;
        src88 <= 16'h1876;
        src89 <= 16'hcf0c;
        src90 <= 16'h847d;
        src91 <= 16'ha621;
        src92 <= 16'hfeb9;
        src93 <= 16'hfc0f;
        src94 <= 16'habe;
        src95 <= 16'h765e;
        src96 <= 16'hcada;
        src97 <= 16'heab5;
        src98 <= 16'h2253;
        src99 <= 16'hb82e;
        src100 <= 16'hf437;
        src101 <= 16'h79f8;
        src102 <= 16'h1a4a;
        src103 <= 16'h5949;
        src104 <= 16'h4542;
        src105 <= 16'h87ca;
        src106 <= 16'hd19d;
        src107 <= 16'h817;
        src108 <= 16'h56a3;
        src109 <= 16'hf5e5;
        src110 <= 16'hdc3f;
        src111 <= 16'h1378;
        src112 <= 16'h9039;
        src113 <= 16'h4c90;
        src114 <= 16'h4cd8;
        src115 <= 16'h5384;
        src116 <= 16'hecf1;
        src117 <= 16'h9289;
        src118 <= 16'h878b;
        src119 <= 16'he9f2;
        src120 <= 16'hc684;
        src121 <= 16'hf21a;
        src122 <= 16'h5981;
        src123 <= 16'hab9e;
        src124 <= 16'hfe2a;
        src125 <= 16'h3597;
        src126 <= 16'h1e0f;
        src127 <= 16'he670;
        src128 <= 16'hbe99;
        src129 <= 16'hbd21;
        src130 <= 16'h447d;
        src131 <= 16'h77ea;
        src132 <= 16'hf8bd;
        src133 <= 16'h55ef;
        src134 <= 16'h6d8e;
        src135 <= 16'hd42c;
        src136 <= 16'hb162;
        src137 <= 16'h4c2;
        src138 <= 16'ha03a;
        src139 <= 16'hb12e;
        src140 <= 16'h7504;
        src141 <= 16'h50f1;
        src142 <= 16'hcc6a;
        src143 <= 16'h9a91;
        src144 <= 16'h4a24;
        src145 <= 16'h8751;
        src146 <= 16'ha8ca;
        src147 <= 16'hcb64;
        src148 <= 16'hc548;
        src149 <= 16'h7356;
        src150 <= 16'h19fe;
        src151 <= 16'hb861;
        src152 <= 16'h3f28;
        src153 <= 16'h1872;
        src154 <= 16'hd985;
        src155 <= 16'hafd5;
        src156 <= 16'hc979;
        src157 <= 16'hff5c;
        src158 <= 16'h9aab;
        src159 <= 16'h199e;
        src160 <= 16'hca97;
        src161 <= 16'hb6d9;
        src162 <= 16'hd14e;
        src163 <= 16'h34d3;
        src164 <= 16'h23fb;
        src165 <= 16'ha4c;
        src166 <= 16'h9e27;
        src167 <= 16'h1331;
        src168 <= 16'he3d1;
        src169 <= 16'hbed9;
        src170 <= 16'hb5f8;
        src171 <= 16'h9e92;
        src172 <= 16'h9f89;
        src173 <= 16'hf33;
        src174 <= 16'h41f9;
        src175 <= 16'h391;
        src176 <= 16'h584b;
        src177 <= 16'he703;
        src178 <= 16'h3524;
        src179 <= 16'h7375;
        src180 <= 16'he868;
        src181 <= 16'h9f0;
        src182 <= 16'ha44f;
        src183 <= 16'ha96;
        src184 <= 16'hc6f8;
        exp <= 24'h5c8e15;
        #1
        src0 <= 16'h6bb6;
        src1 <= 16'h4cdb;
        src2 <= 16'h688b;
        src3 <= 16'h9615;
        src4 <= 16'h8545;
        src5 <= 16'h5501;
        src6 <= 16'hb5a1;
        src7 <= 16'h5f09;
        src8 <= 16'h6f8;
        src9 <= 16'hcf4a;
        src10 <= 16'h83b;
        src11 <= 16'hbfef;
        src12 <= 16'h9b6c;
        src13 <= 16'h7e63;
        src14 <= 16'h164f;
        src15 <= 16'h1732;
        src16 <= 16'h8fef;
        src17 <= 16'h9269;
        src18 <= 16'h215b;
        src19 <= 16'hd403;
        src20 <= 16'hb7e1;
        src21 <= 16'h5c16;
        src22 <= 16'h4f18;
        src23 <= 16'h18fc;
        src24 <= 16'h7c8e;
        src25 <= 16'hd0b3;
        src26 <= 16'h945f;
        src27 <= 16'h1c8;
        src28 <= 16'h473a;
        src29 <= 16'h3d;
        src30 <= 16'hd3a3;
        src31 <= 16'h7ed9;
        src32 <= 16'h8d1d;
        src33 <= 16'hc1c9;
        src34 <= 16'hf5;
        src35 <= 16'hd4a6;
        src36 <= 16'h155e;
        src37 <= 16'h7be9;
        src38 <= 16'h5f96;
        src39 <= 16'h7fb7;
        src40 <= 16'hb917;
        src41 <= 16'hb040;
        src42 <= 16'h866b;
        src43 <= 16'hef75;
        src44 <= 16'h75b7;
        src45 <= 16'h6301;
        src46 <= 16'h4aba;
        src47 <= 16'hc0a;
        src48 <= 16'h585a;
        src49 <= 16'h89bd;
        src50 <= 16'h457;
        src51 <= 16'h5a2;
        src52 <= 16'h3131;
        src53 <= 16'h8cde;
        src54 <= 16'hb094;
        src55 <= 16'h60bc;
        src56 <= 16'hd95;
        src57 <= 16'hbe22;
        src58 <= 16'h9b71;
        src59 <= 16'hc3b2;
        src60 <= 16'hd058;
        src61 <= 16'h7b5e;
        src62 <= 16'h8973;
        src63 <= 16'h60fc;
        src64 <= 16'h8375;
        src65 <= 16'h50c6;
        src66 <= 16'hf363;
        src67 <= 16'h70b5;
        src68 <= 16'h249e;
        src69 <= 16'h9643;
        src70 <= 16'hfa2a;
        src71 <= 16'h239c;
        src72 <= 16'h45d2;
        src73 <= 16'h62e8;
        src74 <= 16'hfb82;
        src75 <= 16'h4f10;
        src76 <= 16'h598;
        src77 <= 16'h5c04;
        src78 <= 16'h5a7c;
        src79 <= 16'h33a1;
        src80 <= 16'hccf6;
        src81 <= 16'h7338;
        src82 <= 16'h3e48;
        src83 <= 16'h95e0;
        src84 <= 16'h38af;
        src85 <= 16'hfdb7;
        src86 <= 16'h2b3e;
        src87 <= 16'hd56d;
        src88 <= 16'he962;
        src89 <= 16'h47f9;
        src90 <= 16'h20ee;
        src91 <= 16'h41e0;
        src92 <= 16'h3167;
        src93 <= 16'he86b;
        src94 <= 16'h82c3;
        src95 <= 16'hf814;
        src96 <= 16'h5e10;
        src97 <= 16'ha2f0;
        src98 <= 16'h7fc7;
        src99 <= 16'h5237;
        src100 <= 16'hb7bd;
        src101 <= 16'h3915;
        src102 <= 16'hc88a;
        src103 <= 16'he8c9;
        src104 <= 16'h4d9d;
        src105 <= 16'h6324;
        src106 <= 16'h463c;
        src107 <= 16'h3821;
        src108 <= 16'he3e1;
        src109 <= 16'h1333;
        src110 <= 16'h4408;
        src111 <= 16'ha33c;
        src112 <= 16'h258;
        src113 <= 16'he3e4;
        src114 <= 16'ha0d8;
        src115 <= 16'he064;
        src116 <= 16'h300b;
        src117 <= 16'haa73;
        src118 <= 16'h1e36;
        src119 <= 16'h9497;
        src120 <= 16'haba0;
        src121 <= 16'h6976;
        src122 <= 16'h64ca;
        src123 <= 16'h7d74;
        src124 <= 16'hfba8;
        src125 <= 16'h180d;
        src126 <= 16'hfcf5;
        src127 <= 16'hcd54;
        src128 <= 16'he1b3;
        src129 <= 16'h9b17;
        src130 <= 16'h7235;
        src131 <= 16'h6f8b;
        src132 <= 16'h691a;
        src133 <= 16'h26c0;
        src134 <= 16'hd1ee;
        src135 <= 16'hc66a;
        src136 <= 16'h7941;
        src137 <= 16'hc9dd;
        src138 <= 16'h1480;
        src139 <= 16'h6fd4;
        src140 <= 16'h1f96;
        src141 <= 16'hc0;
        src142 <= 16'h6d3b;
        src143 <= 16'h17bd;
        src144 <= 16'ha2be;
        src145 <= 16'h91c6;
        src146 <= 16'h2341;
        src147 <= 16'hb5eb;
        src148 <= 16'h34af;
        src149 <= 16'h3304;
        src150 <= 16'h348d;
        src151 <= 16'h2e6b;
        src152 <= 16'h52ee;
        src153 <= 16'hc0ab;
        src154 <= 16'h4178;
        src155 <= 16'h7ffd;
        src156 <= 16'ha217;
        src157 <= 16'h8613;
        src158 <= 16'h6dd9;
        src159 <= 16'hef96;
        src160 <= 16'h28dc;
        src161 <= 16'h1968;
        src162 <= 16'h6277;
        src163 <= 16'h1a95;
        src164 <= 16'h4a58;
        src165 <= 16'hbbf4;
        src166 <= 16'h50c0;
        src167 <= 16'hff4c;
        src168 <= 16'hab8f;
        src169 <= 16'h3ef1;
        src170 <= 16'he51b;
        src171 <= 16'hf115;
        src172 <= 16'h7b2c;
        src173 <= 16'h3c7;
        src174 <= 16'h3e28;
        src175 <= 16'h8fb8;
        src176 <= 16'h98fb;
        src177 <= 16'h3492;
        src178 <= 16'h7ba7;
        src179 <= 16'h589;
        src180 <= 16'ha77a;
        src181 <= 16'h80f5;
        src182 <= 16'h27a0;
        src183 <= 16'h51f4;
        src184 <= 16'h43f2;
        exp <= 24'h549070;
        #1
        src0 <= 16'h26ce;
        src1 <= 16'h80a;
        src2 <= 16'h6b48;
        src3 <= 16'hf526;
        src4 <= 16'h3cc2;
        src5 <= 16'h5f10;
        src6 <= 16'h456;
        src7 <= 16'hd744;
        src8 <= 16'h3fa9;
        src9 <= 16'h2fef;
        src10 <= 16'h6d4a;
        src11 <= 16'h80eb;
        src12 <= 16'h4bb4;
        src13 <= 16'hb20a;
        src14 <= 16'h79c8;
        src15 <= 16'h943e;
        src16 <= 16'h8810;
        src17 <= 16'hb3a0;
        src18 <= 16'hb8c5;
        src19 <= 16'hc9cd;
        src20 <= 16'h700d;
        src21 <= 16'hef2c;
        src22 <= 16'h1959;
        src23 <= 16'hacca;
        src24 <= 16'h8746;
        src25 <= 16'h9af4;
        src26 <= 16'h608e;
        src27 <= 16'h7e4e;
        src28 <= 16'h87ea;
        src29 <= 16'ha195;
        src30 <= 16'h5334;
        src31 <= 16'h4f78;
        src32 <= 16'he688;
        src33 <= 16'h61c8;
        src34 <= 16'hb335;
        src35 <= 16'h4964;
        src36 <= 16'h2328;
        src37 <= 16'hde60;
        src38 <= 16'hc82b;
        src39 <= 16'h9ce5;
        src40 <= 16'hd0de;
        src41 <= 16'hbbd4;
        src42 <= 16'he1b2;
        src43 <= 16'h45c1;
        src44 <= 16'h4750;
        src45 <= 16'hda28;
        src46 <= 16'hb6f0;
        src47 <= 16'h6042;
        src48 <= 16'h6a68;
        src49 <= 16'h4991;
        src50 <= 16'h5c36;
        src51 <= 16'h432d;
        src52 <= 16'h6e0b;
        src53 <= 16'h966e;
        src54 <= 16'h3a97;
        src55 <= 16'h7a35;
        src56 <= 16'h34b4;
        src57 <= 16'h5bd5;
        src58 <= 16'hbf07;
        src59 <= 16'hc2ce;
        src60 <= 16'ha743;
        src61 <= 16'h4333;
        src62 <= 16'h5256;
        src63 <= 16'ha99a;
        src64 <= 16'hef1b;
        src65 <= 16'he826;
        src66 <= 16'h69;
        src67 <= 16'h5437;
        src68 <= 16'hbaa0;
        src69 <= 16'hdf44;
        src70 <= 16'hcf10;
        src71 <= 16'h3883;
        src72 <= 16'h94e7;
        src73 <= 16'h465c;
        src74 <= 16'ha752;
        src75 <= 16'he3c6;
        src76 <= 16'h100;
        src77 <= 16'h387b;
        src78 <= 16'h3919;
        src79 <= 16'hc2b4;
        src80 <= 16'h9120;
        src81 <= 16'he400;
        src82 <= 16'hce25;
        src83 <= 16'h57d7;
        src84 <= 16'ha49e;
        src85 <= 16'hd567;
        src86 <= 16'h5ba0;
        src87 <= 16'h3408;
        src88 <= 16'h6a73;
        src89 <= 16'h6a9b;
        src90 <= 16'h4eba;
        src91 <= 16'h9d73;
        src92 <= 16'hddf3;
        src93 <= 16'hca04;
        src94 <= 16'hc88a;
        src95 <= 16'h8082;
        src96 <= 16'hbcc1;
        src97 <= 16'h73fd;
        src98 <= 16'hab28;
        src99 <= 16'h2fae;
        src100 <= 16'ha9f9;
        src101 <= 16'h251b;
        src102 <= 16'h526e;
        src103 <= 16'he5c5;
        src104 <= 16'h3b41;
        src105 <= 16'ha54b;
        src106 <= 16'he640;
        src107 <= 16'he1d3;
        src108 <= 16'he89c;
        src109 <= 16'hbcf0;
        src110 <= 16'hd9d7;
        src111 <= 16'hc26d;
        src112 <= 16'hdf24;
        src113 <= 16'hfc77;
        src114 <= 16'hac63;
        src115 <= 16'h2335;
        src116 <= 16'h56f4;
        src117 <= 16'h10d7;
        src118 <= 16'h8ca2;
        src119 <= 16'h2cb;
        src120 <= 16'h5622;
        src121 <= 16'h5ff0;
        src122 <= 16'h98a9;
        src123 <= 16'h8c46;
        src124 <= 16'hf7df;
        src125 <= 16'h2211;
        src126 <= 16'h85f9;
        src127 <= 16'h1135;
        src128 <= 16'hd208;
        src129 <= 16'h68ab;
        src130 <= 16'h6242;
        src131 <= 16'hd7d3;
        src132 <= 16'h4862;
        src133 <= 16'h24c8;
        src134 <= 16'h77c8;
        src135 <= 16'hb999;
        src136 <= 16'h498f;
        src137 <= 16'h3469;
        src138 <= 16'h7221;
        src139 <= 16'hc1b0;
        src140 <= 16'h91c8;
        src141 <= 16'hf613;
        src142 <= 16'h895f;
        src143 <= 16'h3ccf;
        src144 <= 16'h6a4b;
        src145 <= 16'h59a6;
        src146 <= 16'h3935;
        src147 <= 16'h574b;
        src148 <= 16'h16d2;
        src149 <= 16'h1731;
        src150 <= 16'h2767;
        src151 <= 16'h143d;
        src152 <= 16'hcc0;
        src153 <= 16'hb203;
        src154 <= 16'hf312;
        src155 <= 16'h1920;
        src156 <= 16'hf3b0;
        src157 <= 16'h4071;
        src158 <= 16'h7fa1;
        src159 <= 16'h86a3;
        src160 <= 16'hb18c;
        src161 <= 16'h1d08;
        src162 <= 16'h5afd;
        src163 <= 16'h2690;
        src164 <= 16'h9d52;
        src165 <= 16'h193d;
        src166 <= 16'h942b;
        src167 <= 16'hfaa7;
        src168 <= 16'hd164;
        src169 <= 16'h79c9;
        src170 <= 16'h161d;
        src171 <= 16'h4707;
        src172 <= 16'hc6e7;
        src173 <= 16'h2fe0;
        src174 <= 16'he78a;
        src175 <= 16'h7160;
        src176 <= 16'ha91e;
        src177 <= 16'hd201;
        src178 <= 16'h3a30;
        src179 <= 16'hd6ab;
        src180 <= 16'h2d5d;
        src181 <= 16'h4159;
        src182 <= 16'h7ddc;
        src183 <= 16'h73d6;
        src184 <= 16'hc222;
        exp <= 24'h5cbd4c;
        #1
        src0 <= 16'hfa48;
        src1 <= 16'hde98;
        src2 <= 16'hf5e;
        src3 <= 16'h8e30;
        src4 <= 16'h2646;
        src5 <= 16'h8621;
        src6 <= 16'h5bc9;
        src7 <= 16'ha4db;
        src8 <= 16'h7b7;
        src9 <= 16'h35a8;
        src10 <= 16'h9c8e;
        src11 <= 16'h78ca;
        src12 <= 16'h3ce0;
        src13 <= 16'h6408;
        src14 <= 16'h4853;
        src15 <= 16'hf305;
        src16 <= 16'hacd;
        src17 <= 16'hf7be;
        src18 <= 16'hec16;
        src19 <= 16'hc234;
        src20 <= 16'h7ad6;
        src21 <= 16'hb469;
        src22 <= 16'h7bac;
        src23 <= 16'h9966;
        src24 <= 16'hf2f1;
        src25 <= 16'he684;
        src26 <= 16'he4f9;
        src27 <= 16'h40ed;
        src28 <= 16'h5d4b;
        src29 <= 16'hd7e7;
        src30 <= 16'hb962;
        src31 <= 16'h669c;
        src32 <= 16'h9667;
        src33 <= 16'h5058;
        src34 <= 16'hc3fa;
        src35 <= 16'hd92f;
        src36 <= 16'h140;
        src37 <= 16'h4b74;
        src38 <= 16'h39d5;
        src39 <= 16'hda39;
        src40 <= 16'h78db;
        src41 <= 16'h9d4d;
        src42 <= 16'h9251;
        src43 <= 16'h51e5;
        src44 <= 16'ha333;
        src45 <= 16'h5acf;
        src46 <= 16'h9598;
        src47 <= 16'hc953;
        src48 <= 16'hd88b;
        src49 <= 16'h573a;
        src50 <= 16'h1ba0;
        src51 <= 16'h84cd;
        src52 <= 16'h4562;
        src53 <= 16'h13c1;
        src54 <= 16'h6346;
        src55 <= 16'hda7;
        src56 <= 16'h6576;
        src57 <= 16'hc2ee;
        src58 <= 16'h69ba;
        src59 <= 16'hb774;
        src60 <= 16'h6763;
        src61 <= 16'h165f;
        src62 <= 16'h33cf;
        src63 <= 16'hd85;
        src64 <= 16'ha538;
        src65 <= 16'h9119;
        src66 <= 16'ha6f8;
        src67 <= 16'h83e4;
        src68 <= 16'h6195;
        src69 <= 16'he992;
        src70 <= 16'h47cf;
        src71 <= 16'h6397;
        src72 <= 16'h4c90;
        src73 <= 16'hb8e2;
        src74 <= 16'h8ade;
        src75 <= 16'hd5e0;
        src76 <= 16'he172;
        src77 <= 16'h2985;
        src78 <= 16'hd870;
        src79 <= 16'h6b84;
        src80 <= 16'hecba;
        src81 <= 16'ha0ce;
        src82 <= 16'h4c39;
        src83 <= 16'he59f;
        src84 <= 16'h48d6;
        src85 <= 16'h5694;
        src86 <= 16'he9eb;
        src87 <= 16'hcf4c;
        src88 <= 16'h44e4;
        src89 <= 16'ha2a4;
        src90 <= 16'hb4dc;
        src91 <= 16'h71f7;
        src92 <= 16'he26e;
        src93 <= 16'h2daf;
        src94 <= 16'haf2c;
        src95 <= 16'hfaa6;
        src96 <= 16'ha752;
        src97 <= 16'h4bf9;
        src98 <= 16'h1a17;
        src99 <= 16'h4b3;
        src100 <= 16'ha29c;
        src101 <= 16'hb8a0;
        src102 <= 16'he117;
        src103 <= 16'h2bf7;
        src104 <= 16'h1c2c;
        src105 <= 16'hac8f;
        src106 <= 16'h7275;
        src107 <= 16'hdd70;
        src108 <= 16'h5ea9;
        src109 <= 16'hd84c;
        src110 <= 16'h40d3;
        src111 <= 16'hba1a;
        src112 <= 16'h918b;
        src113 <= 16'hd213;
        src114 <= 16'h2258;
        src115 <= 16'h5536;
        src116 <= 16'hd734;
        src117 <= 16'h398f;
        src118 <= 16'h537c;
        src119 <= 16'ha095;
        src120 <= 16'h27f;
        src121 <= 16'hb213;
        src122 <= 16'hf733;
        src123 <= 16'hde75;
        src124 <= 16'h8d4c;
        src125 <= 16'ha8bf;
        src126 <= 16'h6e6d;
        src127 <= 16'hb408;
        src128 <= 16'h37f3;
        src129 <= 16'h1d86;
        src130 <= 16'hb72d;
        src131 <= 16'he21f;
        src132 <= 16'h91eb;
        src133 <= 16'hbf1a;
        src134 <= 16'h1ee5;
        src135 <= 16'hca42;
        src136 <= 16'h46d;
        src137 <= 16'hd85;
        src138 <= 16'h87cc;
        src139 <= 16'h1302;
        src140 <= 16'hf717;
        src141 <= 16'hce93;
        src142 <= 16'ha083;
        src143 <= 16'hdff9;
        src144 <= 16'heca7;
        src145 <= 16'h38e8;
        src146 <= 16'h5aa6;
        src147 <= 16'he8b4;
        src148 <= 16'hdda4;
        src149 <= 16'h6c60;
        src150 <= 16'h1773;
        src151 <= 16'he5fb;
        src152 <= 16'h1df7;
        src153 <= 16'h3461;
        src154 <= 16'h747a;
        src155 <= 16'h3ae6;
        src156 <= 16'hee0b;
        src157 <= 16'hfc96;
        src158 <= 16'he1ce;
        src159 <= 16'hb2cf;
        src160 <= 16'hba76;
        src161 <= 16'h9eaf;
        src162 <= 16'h50a7;
        src163 <= 16'h8604;
        src164 <= 16'h7edd;
        src165 <= 16'hcfea;
        src166 <= 16'h28e2;
        src167 <= 16'hfd46;
        src168 <= 16'h401;
        src169 <= 16'h9128;
        src170 <= 16'h52bf;
        src171 <= 16'hb57f;
        src172 <= 16'hf4e8;
        src173 <= 16'h4572;
        src174 <= 16'h6b83;
        src175 <= 16'h9631;
        src176 <= 16'h850;
        src177 <= 16'hb46a;
        src178 <= 16'h2a60;
        src179 <= 16'h399f;
        src180 <= 16'h98c6;
        src181 <= 16'habd2;
        src182 <= 16'h371;
        src183 <= 16'h3852;
        src184 <= 16'h4133;
        exp <= 24'h5f9d5e;
        #1
        src0 <= 16'h63d1;
        src1 <= 16'h4ff;
        src2 <= 16'h45cc;
        src3 <= 16'h7831;
        src4 <= 16'h42f0;
        src5 <= 16'h69e6;
        src6 <= 16'hc3ff;
        src7 <= 16'h5f62;
        src8 <= 16'hd377;
        src9 <= 16'h88b8;
        src10 <= 16'h7ec;
        src11 <= 16'h4fe3;
        src12 <= 16'h4c48;
        src13 <= 16'h44f6;
        src14 <= 16'h2519;
        src15 <= 16'h56c0;
        src16 <= 16'hd9cd;
        src17 <= 16'hf947;
        src18 <= 16'hd9c1;
        src19 <= 16'hfdf4;
        src20 <= 16'ha17f;
        src21 <= 16'h51ce;
        src22 <= 16'hca9b;
        src23 <= 16'hbf26;
        src24 <= 16'hd6d0;
        src25 <= 16'h129;
        src26 <= 16'hf0cb;
        src27 <= 16'hdb60;
        src28 <= 16'hc361;
        src29 <= 16'h5ad3;
        src30 <= 16'h5142;
        src31 <= 16'h2aae;
        src32 <= 16'h8f48;
        src33 <= 16'hba41;
        src34 <= 16'h95d9;
        src35 <= 16'ha462;
        src36 <= 16'h847f;
        src37 <= 16'h4787;
        src38 <= 16'h3779;
        src39 <= 16'h862;
        src40 <= 16'h7d03;
        src41 <= 16'h946f;
        src42 <= 16'h27bb;
        src43 <= 16'h7934;
        src44 <= 16'hc264;
        src45 <= 16'he9d5;
        src46 <= 16'h57fe;
        src47 <= 16'h2f55;
        src48 <= 16'hab7b;
        src49 <= 16'he465;
        src50 <= 16'h42cc;
        src51 <= 16'h1ddb;
        src52 <= 16'ha8b9;
        src53 <= 16'ha438;
        src54 <= 16'h358;
        src55 <= 16'he4d4;
        src56 <= 16'h2e8;
        src57 <= 16'hf62e;
        src58 <= 16'h7b94;
        src59 <= 16'h8bda;
        src60 <= 16'h8ea9;
        src61 <= 16'hd90f;
        src62 <= 16'he8dd;
        src63 <= 16'h13c3;
        src64 <= 16'hf5b6;
        src65 <= 16'h29a7;
        src66 <= 16'h693c;
        src67 <= 16'h4678;
        src68 <= 16'hccb3;
        src69 <= 16'h7dc7;
        src70 <= 16'h2b68;
        src71 <= 16'hc1d1;
        src72 <= 16'hbb11;
        src73 <= 16'h526c;
        src74 <= 16'h933;
        src75 <= 16'h4a42;
        src76 <= 16'h6a88;
        src77 <= 16'hef0a;
        src78 <= 16'hb0b4;
        src79 <= 16'h96cd;
        src80 <= 16'hbd46;
        src81 <= 16'h4be;
        src82 <= 16'hf5d5;
        src83 <= 16'h58cf;
        src84 <= 16'h676;
        src85 <= 16'h36f0;
        src86 <= 16'hea62;
        src87 <= 16'h1e07;
        src88 <= 16'h5168;
        src89 <= 16'hb3dd;
        src90 <= 16'h44b2;
        src91 <= 16'h3a51;
        src92 <= 16'h70dc;
        src93 <= 16'hd933;
        src94 <= 16'ha77d;
        src95 <= 16'h410f;
        src96 <= 16'hbeb2;
        src97 <= 16'h85a0;
        src98 <= 16'h30b4;
        src99 <= 16'h500a;
        src100 <= 16'hcf2d;
        src101 <= 16'h3d64;
        src102 <= 16'h675;
        src103 <= 16'he37;
        src104 <= 16'hd2da;
        src105 <= 16'hea31;
        src106 <= 16'h35fc;
        src107 <= 16'h53e;
        src108 <= 16'hb523;
        src109 <= 16'hc2c8;
        src110 <= 16'h702d;
        src111 <= 16'hc630;
        src112 <= 16'hb0d;
        src113 <= 16'he62b;
        src114 <= 16'h4eaf;
        src115 <= 16'h310c;
        src116 <= 16'h16d0;
        src117 <= 16'hdc75;
        src118 <= 16'h2c7f;
        src119 <= 16'h1800;
        src120 <= 16'h9c4a;
        src121 <= 16'hb939;
        src122 <= 16'hca7f;
        src123 <= 16'hacc1;
        src124 <= 16'hafa6;
        src125 <= 16'h5ce4;
        src126 <= 16'h564a;
        src127 <= 16'h77aa;
        src128 <= 16'hdb72;
        src129 <= 16'hfcd4;
        src130 <= 16'h53f4;
        src131 <= 16'h4be2;
        src132 <= 16'had03;
        src133 <= 16'hea99;
        src134 <= 16'hd10b;
        src135 <= 16'h6129;
        src136 <= 16'hd3d2;
        src137 <= 16'hbb3b;
        src138 <= 16'ha84c;
        src139 <= 16'h6e09;
        src140 <= 16'hccb2;
        src141 <= 16'ha15d;
        src142 <= 16'hb744;
        src143 <= 16'hbac3;
        src144 <= 16'ha32b;
        src145 <= 16'h6e63;
        src146 <= 16'h671a;
        src147 <= 16'he0eb;
        src148 <= 16'h3ef;
        src149 <= 16'h9e3d;
        src150 <= 16'hbe37;
        src151 <= 16'h9a96;
        src152 <= 16'h43b2;
        src153 <= 16'h7fed;
        src154 <= 16'h4ff0;
        src155 <= 16'hceab;
        src156 <= 16'h8f82;
        src157 <= 16'h4e53;
        src158 <= 16'h4629;
        src159 <= 16'h6d45;
        src160 <= 16'h4b31;
        src161 <= 16'h33b4;
        src162 <= 16'hd25b;
        src163 <= 16'hfcc2;
        src164 <= 16'hcfa4;
        src165 <= 16'h2b03;
        src166 <= 16'h30da;
        src167 <= 16'heee2;
        src168 <= 16'ha7;
        src169 <= 16'h95e3;
        src170 <= 16'h705f;
        src171 <= 16'hd164;
        src172 <= 16'h572f;
        src173 <= 16'h89c7;
        src174 <= 16'h198;
        src175 <= 16'h2f68;
        src176 <= 16'h8ffc;
        src177 <= 16'he218;
        src178 <= 16'h8f20;
        src179 <= 16'h7940;
        src180 <= 16'h7e1a;
        src181 <= 16'h8efe;
        src182 <= 16'h9df4;
        src183 <= 16'h512d;
        src184 <= 16'hcf80;
        exp <= 24'h5d3981;
        #1
        src0 <= 16'heef6;
        src1 <= 16'hc119;
        src2 <= 16'h7e8d;
        src3 <= 16'h6dac;
        src4 <= 16'h2087;
        src5 <= 16'hbcad;
        src6 <= 16'h19ad;
        src7 <= 16'h5142;
        src8 <= 16'h8487;
        src9 <= 16'hac79;
        src10 <= 16'h1d3c;
        src11 <= 16'hfa84;
        src12 <= 16'h3310;
        src13 <= 16'h3e2b;
        src14 <= 16'hb2f2;
        src15 <= 16'hf3da;
        src16 <= 16'h9dd2;
        src17 <= 16'hfe2;
        src18 <= 16'hd864;
        src19 <= 16'hdf2d;
        src20 <= 16'ha5d6;
        src21 <= 16'h105a;
        src22 <= 16'hc0e7;
        src23 <= 16'h69ad;
        src24 <= 16'h386a;
        src25 <= 16'h5715;
        src26 <= 16'h4a04;
        src27 <= 16'ha0b3;
        src28 <= 16'hcf3c;
        src29 <= 16'hc2ce;
        src30 <= 16'h1d73;
        src31 <= 16'h31ed;
        src32 <= 16'h9adb;
        src33 <= 16'h510;
        src34 <= 16'h8434;
        src35 <= 16'h8b94;
        src36 <= 16'hfc8d;
        src37 <= 16'h8e9a;
        src38 <= 16'h3dd6;
        src39 <= 16'h17d;
        src40 <= 16'he55c;
        src41 <= 16'h692c;
        src42 <= 16'he28c;
        src43 <= 16'h1a94;
        src44 <= 16'hd57e;
        src45 <= 16'h8641;
        src46 <= 16'he799;
        src47 <= 16'h9811;
        src48 <= 16'h38e4;
        src49 <= 16'h3d02;
        src50 <= 16'h2572;
        src51 <= 16'h10ae;
        src52 <= 16'h495c;
        src53 <= 16'hdb46;
        src54 <= 16'h4a6f;
        src55 <= 16'ha891;
        src56 <= 16'hc705;
        src57 <= 16'hbdc9;
        src58 <= 16'h846;
        src59 <= 16'hc764;
        src60 <= 16'h1854;
        src61 <= 16'h4145;
        src62 <= 16'h4678;
        src63 <= 16'hb539;
        src64 <= 16'h36c5;
        src65 <= 16'h66c8;
        src66 <= 16'h5cab;
        src67 <= 16'hf537;
        src68 <= 16'he2bc;
        src69 <= 16'h6d54;
        src70 <= 16'h811e;
        src71 <= 16'h30e4;
        src72 <= 16'hef4d;
        src73 <= 16'h816;
        src74 <= 16'hd291;
        src75 <= 16'h9aab;
        src76 <= 16'hb1af;
        src77 <= 16'h8596;
        src78 <= 16'ha6f5;
        src79 <= 16'hc440;
        src80 <= 16'h661f;
        src81 <= 16'hbe04;
        src82 <= 16'hab34;
        src83 <= 16'hdd07;
        src84 <= 16'h44f3;
        src85 <= 16'h92ec;
        src86 <= 16'h74fb;
        src87 <= 16'ha04e;
        src88 <= 16'he5d1;
        src89 <= 16'hfdc8;
        src90 <= 16'hdf76;
        src91 <= 16'h4119;
        src92 <= 16'h99ff;
        src93 <= 16'ha986;
        src94 <= 16'hc047;
        src95 <= 16'hb3f4;
        src96 <= 16'hd287;
        src97 <= 16'h2c26;
        src98 <= 16'h3364;
        src99 <= 16'he1fb;
        src100 <= 16'h9fed;
        src101 <= 16'h5a7c;
        src102 <= 16'h5eba;
        src103 <= 16'hfd48;
        src104 <= 16'h2ade;
        src105 <= 16'h7533;
        src106 <= 16'h6375;
        src107 <= 16'h21f7;
        src108 <= 16'h6465;
        src109 <= 16'h284e;
        src110 <= 16'h7e58;
        src111 <= 16'h2f09;
        src112 <= 16'h478a;
        src113 <= 16'h5a96;
        src114 <= 16'h71f4;
        src115 <= 16'hc48b;
        src116 <= 16'h6cae;
        src117 <= 16'h5479;
        src118 <= 16'h3fd1;
        src119 <= 16'h3b27;
        src120 <= 16'h5b32;
        src121 <= 16'hb27b;
        src122 <= 16'h5d3a;
        src123 <= 16'hdce3;
        src124 <= 16'he4b9;
        src125 <= 16'h5801;
        src126 <= 16'hb2ed;
        src127 <= 16'h4158;
        src128 <= 16'h3cdb;
        src129 <= 16'h61fb;
        src130 <= 16'h61df;
        src131 <= 16'hd6f9;
        src132 <= 16'hc10e;
        src133 <= 16'h417f;
        src134 <= 16'hccdb;
        src135 <= 16'hdcf5;
        src136 <= 16'h4aeb;
        src137 <= 16'h348;
        src138 <= 16'hf3ba;
        src139 <= 16'h5a45;
        src140 <= 16'h89cf;
        src141 <= 16'hb14c;
        src142 <= 16'h2aaa;
        src143 <= 16'h1030;
        src144 <= 16'hbc27;
        src145 <= 16'h549b;
        src146 <= 16'hbb71;
        src147 <= 16'h28be;
        src148 <= 16'hfaa6;
        src149 <= 16'h353f;
        src150 <= 16'h9d0e;
        src151 <= 16'h1b90;
        src152 <= 16'h7bb4;
        src153 <= 16'h20f5;
        src154 <= 16'hb484;
        src155 <= 16'hd9fc;
        src156 <= 16'h5db;
        src157 <= 16'h98fc;
        src158 <= 16'hfe61;
        src159 <= 16'hd7b5;
        src160 <= 16'h9bd1;
        src161 <= 16'hb2e9;
        src162 <= 16'h76dd;
        src163 <= 16'haca9;
        src164 <= 16'h637;
        src165 <= 16'h573d;
        src166 <= 16'h6b1c;
        src167 <= 16'h42c;
        src168 <= 16'ha1b6;
        src169 <= 16'h3496;
        src170 <= 16'h1607;
        src171 <= 16'he0f9;
        src172 <= 16'hb5ee;
        src173 <= 16'h9c5c;
        src174 <= 16'he916;
        src175 <= 16'h6271;
        src176 <= 16'hc12e;
        src177 <= 16'hf483;
        src178 <= 16'h166a;
        src179 <= 16'h1dbb;
        src180 <= 16'h9e9a;
        src181 <= 16'h1b8f;
        src182 <= 16'h9eea;
        src183 <= 16'h4c35;
        src184 <= 16'h53b2;
        exp <= 24'h5c3bbf;
        #1
        src0 <= 16'h3dad;
        src1 <= 16'h628a;
        src2 <= 16'h6dde;
        src3 <= 16'h6e49;
        src4 <= 16'hf2ee;
        src5 <= 16'h2939;
        src6 <= 16'hc03a;
        src7 <= 16'h1061;
        src8 <= 16'h34db;
        src9 <= 16'hd51a;
        src10 <= 16'hf23c;
        src11 <= 16'h33b;
        src12 <= 16'hbc2a;
        src13 <= 16'h5043;
        src14 <= 16'hd2ce;
        src15 <= 16'h518d;
        src16 <= 16'h77cf;
        src17 <= 16'h74a4;
        src18 <= 16'h9673;
        src19 <= 16'hf9fe;
        src20 <= 16'hc201;
        src21 <= 16'h55b7;
        src22 <= 16'hdc0a;
        src23 <= 16'h7d1e;
        src24 <= 16'h3e52;
        src25 <= 16'hd1db;
        src26 <= 16'hca4a;
        src27 <= 16'hb97f;
        src28 <= 16'h89cb;
        src29 <= 16'h3d77;
        src30 <= 16'h122e;
        src31 <= 16'h3b07;
        src32 <= 16'h5a20;
        src33 <= 16'hd93a;
        src34 <= 16'he724;
        src35 <= 16'h8b5a;
        src36 <= 16'h23e;
        src37 <= 16'hf6a4;
        src38 <= 16'hf0f9;
        src39 <= 16'h31ea;
        src40 <= 16'hbda9;
        src41 <= 16'h94bc;
        src42 <= 16'h15fe;
        src43 <= 16'h2289;
        src44 <= 16'h5408;
        src45 <= 16'he3d3;
        src46 <= 16'hf3be;
        src47 <= 16'h1de0;
        src48 <= 16'h342a;
        src49 <= 16'h2733;
        src50 <= 16'h234c;
        src51 <= 16'ha1bc;
        src52 <= 16'h4bbb;
        src53 <= 16'h6ebd;
        src54 <= 16'hf946;
        src55 <= 16'h2db5;
        src56 <= 16'hffb3;
        src57 <= 16'h269c;
        src58 <= 16'haa21;
        src59 <= 16'h706d;
        src60 <= 16'h4628;
        src61 <= 16'h4fab;
        src62 <= 16'h2b3;
        src63 <= 16'h8a11;
        src64 <= 16'h76a2;
        src65 <= 16'h5136;
        src66 <= 16'h564a;
        src67 <= 16'h2fb9;
        src68 <= 16'h5330;
        src69 <= 16'h9af9;
        src70 <= 16'h6465;
        src71 <= 16'h14ea;
        src72 <= 16'hc373;
        src73 <= 16'h50f;
        src74 <= 16'he54;
        src75 <= 16'hfd17;
        src76 <= 16'h63ec;
        src77 <= 16'h6a00;
        src78 <= 16'hd105;
        src79 <= 16'h97ff;
        src80 <= 16'h920d;
        src81 <= 16'hd922;
        src82 <= 16'h54c3;
        src83 <= 16'h149a;
        src84 <= 16'h34e4;
        src85 <= 16'h377a;
        src86 <= 16'h341f;
        src87 <= 16'h81;
        src88 <= 16'h5d7;
        src89 <= 16'hcdb6;
        src90 <= 16'hd2b5;
        src91 <= 16'h44d0;
        src92 <= 16'ha270;
        src93 <= 16'h53fc;
        src94 <= 16'h7d3d;
        src95 <= 16'h200;
        src96 <= 16'h909d;
        src97 <= 16'hc9c3;
        src98 <= 16'h1af5;
        src99 <= 16'h296c;
        src100 <= 16'h8d17;
        src101 <= 16'h7116;
        src102 <= 16'h19bf;
        src103 <= 16'h8243;
        src104 <= 16'hc221;
        src105 <= 16'hcc52;
        src106 <= 16'hf85c;
        src107 <= 16'h648;
        src108 <= 16'hdb86;
        src109 <= 16'hd7b3;
        src110 <= 16'hf57a;
        src111 <= 16'hbfa1;
        src112 <= 16'h1047;
        src113 <= 16'h2d4;
        src114 <= 16'h1add;
        src115 <= 16'h100b;
        src116 <= 16'h8847;
        src117 <= 16'h21d3;
        src118 <= 16'hf0ec;
        src119 <= 16'hce2;
        src120 <= 16'h929d;
        src121 <= 16'hf4b9;
        src122 <= 16'hf2b2;
        src123 <= 16'h423;
        src124 <= 16'h8499;
        src125 <= 16'h314e;
        src126 <= 16'h470c;
        src127 <= 16'hd75;
        src128 <= 16'he278;
        src129 <= 16'hdeb3;
        src130 <= 16'h8df8;
        src131 <= 16'h824e;
        src132 <= 16'h3abf;
        src133 <= 16'h1b23;
        src134 <= 16'h8506;
        src135 <= 16'h4bf5;
        src136 <= 16'he035;
        src137 <= 16'h21b2;
        src138 <= 16'h227c;
        src139 <= 16'h15fa;
        src140 <= 16'hf72;
        src141 <= 16'hefb0;
        src142 <= 16'h4d02;
        src143 <= 16'h723e;
        src144 <= 16'hb516;
        src145 <= 16'h3803;
        src146 <= 16'h181c;
        src147 <= 16'hf4f4;
        src148 <= 16'h3d4e;
        src149 <= 16'hf71d;
        src150 <= 16'h4867;
        src151 <= 16'h1922;
        src152 <= 16'h2dbe;
        src153 <= 16'h893a;
        src154 <= 16'h1ad0;
        src155 <= 16'h2c53;
        src156 <= 16'h6fd0;
        src157 <= 16'h2bf4;
        src158 <= 16'h741f;
        src159 <= 16'h7025;
        src160 <= 16'h2120;
        src161 <= 16'h9666;
        src162 <= 16'ha153;
        src163 <= 16'hd96;
        src164 <= 16'hb3a9;
        src165 <= 16'h26c6;
        src166 <= 16'he72d;
        src167 <= 16'hee70;
        src168 <= 16'h3b0f;
        src169 <= 16'h970e;
        src170 <= 16'h583f;
        src171 <= 16'h9d37;
        src172 <= 16'h2bdf;
        src173 <= 16'h37d9;
        src174 <= 16'h55a1;
        src175 <= 16'h5e38;
        src176 <= 16'h81c;
        src177 <= 16'h74f4;
        src178 <= 16'h8508;
        src179 <= 16'hc18b;
        src180 <= 16'h282b;
        src181 <= 16'hb104;
        src182 <= 16'h7fdc;
        src183 <= 16'h28d7;
        src184 <= 16'h7ac3;
        exp <= 24'h521355;
        #1
        src0 <= 16'hb043;
        src1 <= 16'h153e;
        src2 <= 16'he3f2;
        src3 <= 16'h24cc;
        src4 <= 16'hfd72;
        src5 <= 16'h467c;
        src6 <= 16'h537a;
        src7 <= 16'h8bc;
        src8 <= 16'hf4b4;
        src9 <= 16'h9730;
        src10 <= 16'h6b64;
        src11 <= 16'h8024;
        src12 <= 16'h6cb;
        src13 <= 16'h7410;
        src14 <= 16'hebe5;
        src15 <= 16'hbfc4;
        src16 <= 16'hfb2;
        src17 <= 16'h9d28;
        src18 <= 16'h5265;
        src19 <= 16'hc025;
        src20 <= 16'h484c;
        src21 <= 16'h187b;
        src22 <= 16'h7189;
        src23 <= 16'h92d6;
        src24 <= 16'hd082;
        src25 <= 16'h434b;
        src26 <= 16'hfacd;
        src27 <= 16'hb1cf;
        src28 <= 16'hd0f4;
        src29 <= 16'he391;
        src30 <= 16'hf555;
        src31 <= 16'h993e;
        src32 <= 16'hd523;
        src33 <= 16'hef48;
        src34 <= 16'h55f7;
        src35 <= 16'h7f62;
        src36 <= 16'h134;
        src37 <= 16'h82b;
        src38 <= 16'h1435;
        src39 <= 16'h9a4f;
        src40 <= 16'hcc1;
        src41 <= 16'hbe20;
        src42 <= 16'h30b7;
        src43 <= 16'h29cc;
        src44 <= 16'h944b;
        src45 <= 16'h942;
        src46 <= 16'ha44c;
        src47 <= 16'h1020;
        src48 <= 16'hb1d;
        src49 <= 16'hdeff;
        src50 <= 16'h445b;
        src51 <= 16'h5559;
        src52 <= 16'h73c3;
        src53 <= 16'h11a4;
        src54 <= 16'hcd6e;
        src55 <= 16'h419c;
        src56 <= 16'h7bc0;
        src57 <= 16'h3ec3;
        src58 <= 16'h2f04;
        src59 <= 16'h2186;
        src60 <= 16'h6639;
        src61 <= 16'h2800;
        src62 <= 16'h4ce;
        src63 <= 16'hd8c5;
        src64 <= 16'h5d6f;
        src65 <= 16'hcda9;
        src66 <= 16'h106;
        src67 <= 16'hdabf;
        src68 <= 16'h4439;
        src69 <= 16'ha26b;
        src70 <= 16'hc565;
        src71 <= 16'hd393;
        src72 <= 16'hd552;
        src73 <= 16'hdf18;
        src74 <= 16'he0da;
        src75 <= 16'hd170;
        src76 <= 16'h894d;
        src77 <= 16'had98;
        src78 <= 16'hc6a8;
        src79 <= 16'h58a1;
        src80 <= 16'h4d3f;
        src81 <= 16'hbbd9;
        src82 <= 16'h519f;
        src83 <= 16'h8d56;
        src84 <= 16'hd478;
        src85 <= 16'hcf95;
        src86 <= 16'h8e34;
        src87 <= 16'hf937;
        src88 <= 16'h11b0;
        src89 <= 16'hf2a1;
        src90 <= 16'h62b1;
        src91 <= 16'hc2a6;
        src92 <= 16'hf3d6;
        src93 <= 16'h42ca;
        src94 <= 16'h48e;
        src95 <= 16'haf55;
        src96 <= 16'hb71;
        src97 <= 16'h9dad;
        src98 <= 16'hd875;
        src99 <= 16'haabe;
        src100 <= 16'h6161;
        src101 <= 16'h7568;
        src102 <= 16'h3e90;
        src103 <= 16'h57f4;
        src104 <= 16'h7fb9;
        src105 <= 16'h71d2;
        src106 <= 16'h76f6;
        src107 <= 16'h4bc2;
        src108 <= 16'h949d;
        src109 <= 16'hd6e6;
        src110 <= 16'h635e;
        src111 <= 16'h7e57;
        src112 <= 16'h5f25;
        src113 <= 16'hecdf;
        src114 <= 16'h24e3;
        src115 <= 16'h6e41;
        src116 <= 16'hf8dc;
        src117 <= 16'h6608;
        src118 <= 16'ha5af;
        src119 <= 16'hd73c;
        src120 <= 16'h79a4;
        src121 <= 16'h3c4d;
        src122 <= 16'h7aa5;
        src123 <= 16'hb6a7;
        src124 <= 16'h137d;
        src125 <= 16'h99f9;
        src126 <= 16'hee3c;
        src127 <= 16'h5b55;
        src128 <= 16'h45eb;
        src129 <= 16'hf51b;
        src130 <= 16'hc729;
        src131 <= 16'he38c;
        src132 <= 16'h296;
        src133 <= 16'h67a4;
        src134 <= 16'h3bc7;
        src135 <= 16'he0ec;
        src136 <= 16'ha229;
        src137 <= 16'hba03;
        src138 <= 16'h5c82;
        src139 <= 16'hf904;
        src140 <= 16'hed28;
        src141 <= 16'h4b0c;
        src142 <= 16'hfc0d;
        src143 <= 16'h76d7;
        src144 <= 16'h457f;
        src145 <= 16'hfe1e;
        src146 <= 16'hdcb2;
        src147 <= 16'hc63b;
        src148 <= 16'hc072;
        src149 <= 16'hd8dd;
        src150 <= 16'heaef;
        src151 <= 16'h1869;
        src152 <= 16'hf96c;
        src153 <= 16'hc4b;
        src154 <= 16'hc696;
        src155 <= 16'h4043;
        src156 <= 16'h278a;
        src157 <= 16'hbdfc;
        src158 <= 16'h3e54;
        src159 <= 16'h9e4c;
        src160 <= 16'h3ac2;
        src161 <= 16'h5d25;
        src162 <= 16'h16de;
        src163 <= 16'h2e39;
        src164 <= 16'h61d6;
        src165 <= 16'ha7a1;
        src166 <= 16'hf680;
        src167 <= 16'h40ee;
        src168 <= 16'h6722;
        src169 <= 16'hd2c7;
        src170 <= 16'h5c1;
        src171 <= 16'hbe86;
        src172 <= 16'h10b8;
        src173 <= 16'h74c4;
        src174 <= 16'heb9f;
        src175 <= 16'h12ab;
        src176 <= 16'h9180;
        src177 <= 16'h9f0d;
        src178 <= 16'h958b;
        src179 <= 16'hbdda;
        src180 <= 16'h6ebc;
        src181 <= 16'hafcf;
        src182 <= 16'h1f65;
        src183 <= 16'hd732;
        src184 <= 16'h61e4;
        exp <= 24'h5ee205;
        #1
        src0 <= 16'h359d;
        src1 <= 16'h36cf;
        src2 <= 16'h4adc;
        src3 <= 16'h5798;
        src4 <= 16'heb7a;
        src5 <= 16'h28e0;
        src6 <= 16'h9bfd;
        src7 <= 16'h9bbd;
        src8 <= 16'ha5fd;
        src9 <= 16'he9f7;
        src10 <= 16'h5e31;
        src11 <= 16'h8722;
        src12 <= 16'h3b95;
        src13 <= 16'ha6d1;
        src14 <= 16'h8961;
        src15 <= 16'had17;
        src16 <= 16'he948;
        src17 <= 16'h920a;
        src18 <= 16'h61a2;
        src19 <= 16'he61f;
        src20 <= 16'he43b;
        src21 <= 16'h141e;
        src22 <= 16'hc285;
        src23 <= 16'h361f;
        src24 <= 16'hfb9d;
        src25 <= 16'h3a63;
        src26 <= 16'hbcad;
        src27 <= 16'h4e4;
        src28 <= 16'hf0ab;
        src29 <= 16'h9846;
        src30 <= 16'h64d4;
        src31 <= 16'h8d5e;
        src32 <= 16'h4f88;
        src33 <= 16'hb40d;
        src34 <= 16'h5dfd;
        src35 <= 16'hea83;
        src36 <= 16'h87df;
        src37 <= 16'hf26b;
        src38 <= 16'h6642;
        src39 <= 16'h950d;
        src40 <= 16'hc2d;
        src41 <= 16'h24ee;
        src42 <= 16'hda16;
        src43 <= 16'h48ae;
        src44 <= 16'h4c8b;
        src45 <= 16'h9efe;
        src46 <= 16'h98d8;
        src47 <= 16'ha233;
        src48 <= 16'he16b;
        src49 <= 16'hb88c;
        src50 <= 16'ha333;
        src51 <= 16'h6951;
        src52 <= 16'hc7f3;
        src53 <= 16'h8082;
        src54 <= 16'h416d;
        src55 <= 16'hae79;
        src56 <= 16'h5d06;
        src57 <= 16'h980b;
        src58 <= 16'h7ea6;
        src59 <= 16'h55f7;
        src60 <= 16'h9ac2;
        src61 <= 16'hee72;
        src62 <= 16'hd7a0;
        src63 <= 16'h49c9;
        src64 <= 16'h8ed2;
        src65 <= 16'h114a;
        src66 <= 16'hd4aa;
        src67 <= 16'h2696;
        src68 <= 16'h8476;
        src69 <= 16'hd518;
        src70 <= 16'h5381;
        src71 <= 16'h3a45;
        src72 <= 16'hfee4;
        src73 <= 16'h7ff0;
        src74 <= 16'hb570;
        src75 <= 16'h5a4e;
        src76 <= 16'h97fd;
        src77 <= 16'hf621;
        src78 <= 16'h49ec;
        src79 <= 16'hf37e;
        src80 <= 16'h594e;
        src81 <= 16'h6575;
        src82 <= 16'h4ad5;
        src83 <= 16'h76c1;
        src84 <= 16'h737a;
        src85 <= 16'h6989;
        src86 <= 16'h7486;
        src87 <= 16'hced8;
        src88 <= 16'hc7af;
        src89 <= 16'hee80;
        src90 <= 16'hec15;
        src91 <= 16'h3752;
        src92 <= 16'h82c4;
        src93 <= 16'h5bd7;
        src94 <= 16'h199f;
        src95 <= 16'h5993;
        src96 <= 16'h98c;
        src97 <= 16'ha71c;
        src98 <= 16'hf9ec;
        src99 <= 16'hc54a;
        src100 <= 16'h8dbc;
        src101 <= 16'hd9a9;
        src102 <= 16'hac82;
        src103 <= 16'h712a;
        src104 <= 16'h934a;
        src105 <= 16'hc00a;
        src106 <= 16'he85e;
        src107 <= 16'h4a4f;
        src108 <= 16'h2b10;
        src109 <= 16'hacd6;
        src110 <= 16'hc8de;
        src111 <= 16'ha6f7;
        src112 <= 16'h2f55;
        src113 <= 16'hb234;
        src114 <= 16'h2c25;
        src115 <= 16'ha221;
        src116 <= 16'h9585;
        src117 <= 16'he091;
        src118 <= 16'h249f;
        src119 <= 16'h95cb;
        src120 <= 16'h7d7;
        src121 <= 16'h9297;
        src122 <= 16'h38c6;
        src123 <= 16'hcb43;
        src124 <= 16'h98c;
        src125 <= 16'h1960;
        src126 <= 16'h4897;
        src127 <= 16'h8f21;
        src128 <= 16'hc95e;
        src129 <= 16'hd264;
        src130 <= 16'hc5b2;
        src131 <= 16'hbd24;
        src132 <= 16'hb502;
        src133 <= 16'h9cbe;
        src134 <= 16'hb5c1;
        src135 <= 16'hae75;
        src136 <= 16'hebf1;
        src137 <= 16'hf7f5;
        src138 <= 16'h724c;
        src139 <= 16'hc408;
        src140 <= 16'hfe37;
        src141 <= 16'h15d6;
        src142 <= 16'h4b8f;
        src143 <= 16'h533c;
        src144 <= 16'h70f2;
        src145 <= 16'h65f;
        src146 <= 16'he5ec;
        src147 <= 16'hf9f3;
        src148 <= 16'hd42f;
        src149 <= 16'h9cf3;
        src150 <= 16'he271;
        src151 <= 16'h655e;
        src152 <= 16'h6c91;
        src153 <= 16'h886d;
        src154 <= 16'hc865;
        src155 <= 16'h8cc0;
        src156 <= 16'h2e0;
        src157 <= 16'h4bc5;
        src158 <= 16'h143c;
        src159 <= 16'h871;
        src160 <= 16'hf210;
        src161 <= 16'hdbb3;
        src162 <= 16'h955e;
        src163 <= 16'h7f71;
        src164 <= 16'hdc8c;
        src165 <= 16'h750;
        src166 <= 16'hb5c5;
        src167 <= 16'h86df;
        src168 <= 16'h7e55;
        src169 <= 16'ha25b;
        src170 <= 16'hd535;
        src171 <= 16'ha741;
        src172 <= 16'ha2dd;
        src173 <= 16'h3da9;
        src174 <= 16'h8c4b;
        src175 <= 16'hf26b;
        src176 <= 16'he2e2;
        src177 <= 16'h2ff4;
        src178 <= 16'h63b1;
        src179 <= 16'h63a3;
        src180 <= 16'h6963;
        src181 <= 16'h37f3;
        src182 <= 16'h2ea5;
        src183 <= 16'h60c0;
        src184 <= 16'hb054;
        exp <= 24'h63a5fe;
        #1
        src0 <= 16'h561d;
        src1 <= 16'h65fe;
        src2 <= 16'h5f73;
        src3 <= 16'h51ec;
        src4 <= 16'hc43f;
        src5 <= 16'h5ca7;
        src6 <= 16'h28ad;
        src7 <= 16'he71e;
        src8 <= 16'h6255;
        src9 <= 16'h3e5;
        src10 <= 16'h1330;
        src11 <= 16'h573f;
        src12 <= 16'he89f;
        src13 <= 16'ha35c;
        src14 <= 16'h14d1;
        src15 <= 16'h32ab;
        src16 <= 16'h19;
        src17 <= 16'h729f;
        src18 <= 16'h56f5;
        src19 <= 16'h452e;
        src20 <= 16'h8a4a;
        src21 <= 16'hf88e;
        src22 <= 16'h92ba;
        src23 <= 16'hf065;
        src24 <= 16'h1194;
        src25 <= 16'h780d;
        src26 <= 16'had97;
        src27 <= 16'hcf12;
        src28 <= 16'h555b;
        src29 <= 16'h4df4;
        src30 <= 16'hf974;
        src31 <= 16'h2d3f;
        src32 <= 16'ha0a0;
        src33 <= 16'hc86e;
        src34 <= 16'hc9eb;
        src35 <= 16'hdbf0;
        src36 <= 16'h303c;
        src37 <= 16'ha600;
        src38 <= 16'h6819;
        src39 <= 16'h1d1f;
        src40 <= 16'hba2f;
        src41 <= 16'hd921;
        src42 <= 16'h2e4a;
        src43 <= 16'hd395;
        src44 <= 16'h9587;
        src45 <= 16'h6e3;
        src46 <= 16'h983a;
        src47 <= 16'h2e34;
        src48 <= 16'h2829;
        src49 <= 16'h33e6;
        src50 <= 16'hceb1;
        src51 <= 16'h37df;
        src52 <= 16'hf771;
        src53 <= 16'hcae2;
        src54 <= 16'h7733;
        src55 <= 16'hae05;
        src56 <= 16'he781;
        src57 <= 16'h3b51;
        src58 <= 16'h4731;
        src59 <= 16'h6fce;
        src60 <= 16'hdb4c;
        src61 <= 16'h25bc;
        src62 <= 16'h42ea;
        src63 <= 16'h2493;
        src64 <= 16'hb950;
        src65 <= 16'hb6be;
        src66 <= 16'h3a28;
        src67 <= 16'hc6dc;
        src68 <= 16'h2a62;
        src69 <= 16'hfdc0;
        src70 <= 16'h9687;
        src71 <= 16'h52a8;
        src72 <= 16'h1c7f;
        src73 <= 16'hde96;
        src74 <= 16'hc6a4;
        src75 <= 16'h5d19;
        src76 <= 16'h9afb;
        src77 <= 16'h5c54;
        src78 <= 16'h417;
        src79 <= 16'hc0ec;
        src80 <= 16'hd50c;
        src81 <= 16'he5a0;
        src82 <= 16'h61e;
        src83 <= 16'hbe5c;
        src84 <= 16'hc323;
        src85 <= 16'h45ed;
        src86 <= 16'hc10;
        src87 <= 16'hf82;
        src88 <= 16'h23b9;
        src89 <= 16'h95a0;
        src90 <= 16'he6fd;
        src91 <= 16'ha3f;
        src92 <= 16'hc494;
        src93 <= 16'h9d57;
        src94 <= 16'h3606;
        src95 <= 16'h4ce9;
        src96 <= 16'hf151;
        src97 <= 16'h4674;
        src98 <= 16'hced6;
        src99 <= 16'had9a;
        src100 <= 16'hb469;
        src101 <= 16'h1b81;
        src102 <= 16'h9233;
        src103 <= 16'h2e73;
        src104 <= 16'h8016;
        src105 <= 16'he6ea;
        src106 <= 16'hfc2c;
        src107 <= 16'h8ab8;
        src108 <= 16'h1e18;
        src109 <= 16'he426;
        src110 <= 16'h3b63;
        src111 <= 16'hdc77;
        src112 <= 16'hcc1b;
        src113 <= 16'h5846;
        src114 <= 16'h5bc7;
        src115 <= 16'ha93e;
        src116 <= 16'h62c2;
        src117 <= 16'hb6fc;
        src118 <= 16'h7999;
        src119 <= 16'h1ffa;
        src120 <= 16'h7e9f;
        src121 <= 16'hef2;
        src122 <= 16'h909f;
        src123 <= 16'h43f6;
        src124 <= 16'h5a1b;
        src125 <= 16'h21fa;
        src126 <= 16'h6df9;
        src127 <= 16'h2a64;
        src128 <= 16'h987b;
        src129 <= 16'ha3b4;
        src130 <= 16'h7d37;
        src131 <= 16'h2cfb;
        src132 <= 16'hdc67;
        src133 <= 16'h5cee;
        src134 <= 16'h97bf;
        src135 <= 16'h6c4b;
        src136 <= 16'h149b;
        src137 <= 16'he9af;
        src138 <= 16'h10fb;
        src139 <= 16'hb995;
        src140 <= 16'hb08c;
        src141 <= 16'h2516;
        src142 <= 16'h1dbf;
        src143 <= 16'h3e2;
        src144 <= 16'h279;
        src145 <= 16'h9d75;
        src146 <= 16'h8320;
        src147 <= 16'hf511;
        src148 <= 16'h2f8f;
        src149 <= 16'h55d9;
        src150 <= 16'h4a04;
        src151 <= 16'hf59a;
        src152 <= 16'hb943;
        src153 <= 16'h77a0;
        src154 <= 16'h31a4;
        src155 <= 16'h8088;
        src156 <= 16'haac3;
        src157 <= 16'hf3f1;
        src158 <= 16'hbe76;
        src159 <= 16'h28f3;
        src160 <= 16'h870;
        src161 <= 16'ha5fa;
        src162 <= 16'h4c9c;
        src163 <= 16'h7e67;
        src164 <= 16'h40ee;
        src165 <= 16'h3ff;
        src166 <= 16'h5f28;
        src167 <= 16'hd78f;
        src168 <= 16'hb849;
        src169 <= 16'h26b2;
        src170 <= 16'h3ea3;
        src171 <= 16'ha93b;
        src172 <= 16'hcf9c;
        src173 <= 16'hcb08;
        src174 <= 16'h2b25;
        src175 <= 16'hdf5b;
        src176 <= 16'h8709;
        src177 <= 16'hf174;
        src178 <= 16'hdb2e;
        src179 <= 16'h6a74;
        src180 <= 16'h6eee;
        src181 <= 16'h6554;
        src182 <= 16'h983e;
        src183 <= 16'h43ac;
        src184 <= 16'h844b;
        exp <= 24'h58c4ed;
        #1
        src0 <= 16'hb7f0;
        src1 <= 16'hecb3;
        src2 <= 16'h361;
        src3 <= 16'h2c6f;
        src4 <= 16'h13b6;
        src5 <= 16'h3af3;
        src6 <= 16'h1ac2;
        src7 <= 16'h5f40;
        src8 <= 16'hd02c;
        src9 <= 16'ha3d9;
        src10 <= 16'h84b4;
        src11 <= 16'h25a0;
        src12 <= 16'hf427;
        src13 <= 16'h732a;
        src14 <= 16'he274;
        src15 <= 16'h4efe;
        src16 <= 16'h9687;
        src17 <= 16'ha366;
        src18 <= 16'ha182;
        src19 <= 16'he2fc;
        src20 <= 16'h2276;
        src21 <= 16'h1311;
        src22 <= 16'hbd1e;
        src23 <= 16'h53f7;
        src24 <= 16'h3449;
        src25 <= 16'h558e;
        src26 <= 16'h3845;
        src27 <= 16'h60c2;
        src28 <= 16'h279e;
        src29 <= 16'hbd40;
        src30 <= 16'h2f15;
        src31 <= 16'hd8c4;
        src32 <= 16'h5196;
        src33 <= 16'h9208;
        src34 <= 16'h8cd4;
        src35 <= 16'h48;
        src36 <= 16'h50ff;
        src37 <= 16'h9951;
        src38 <= 16'hb9ab;
        src39 <= 16'hfcb3;
        src40 <= 16'h216c;
        src41 <= 16'h1d19;
        src42 <= 16'hfbd3;
        src43 <= 16'headb;
        src44 <= 16'h1238;
        src45 <= 16'h2d1a;
        src46 <= 16'hc428;
        src47 <= 16'hd7c2;
        src48 <= 16'h346f;
        src49 <= 16'hb8ca;
        src50 <= 16'h7d71;
        src51 <= 16'h1f4f;
        src52 <= 16'h4acc;
        src53 <= 16'h1c56;
        src54 <= 16'h43df;
        src55 <= 16'he5cd;
        src56 <= 16'h3281;
        src57 <= 16'hd8e4;
        src58 <= 16'hfe62;
        src59 <= 16'h5389;
        src60 <= 16'h143e;
        src61 <= 16'hb6a0;
        src62 <= 16'h42e9;
        src63 <= 16'h51b;
        src64 <= 16'he929;
        src65 <= 16'h7b71;
        src66 <= 16'h99ba;
        src67 <= 16'h68b2;
        src68 <= 16'h4d3f;
        src69 <= 16'he33f;
        src70 <= 16'h5b43;
        src71 <= 16'hf7b2;
        src72 <= 16'h3d42;
        src73 <= 16'h3d16;
        src74 <= 16'h2a96;
        src75 <= 16'he1a3;
        src76 <= 16'h6473;
        src77 <= 16'ha877;
        src78 <= 16'h64d0;
        src79 <= 16'h4c7a;
        src80 <= 16'h6769;
        src81 <= 16'h60f8;
        src82 <= 16'he462;
        src83 <= 16'he9d4;
        src84 <= 16'he32b;
        src85 <= 16'he474;
        src86 <= 16'h6543;
        src87 <= 16'h5ca1;
        src88 <= 16'h5ef1;
        src89 <= 16'he789;
        src90 <= 16'h7993;
        src91 <= 16'h6e0c;
        src92 <= 16'h6491;
        src93 <= 16'h3360;
        src94 <= 16'h7e54;
        src95 <= 16'h94da;
        src96 <= 16'h77d5;
        src97 <= 16'hece2;
        src98 <= 16'hb056;
        src99 <= 16'h6c23;
        src100 <= 16'h31e0;
        src101 <= 16'hfbe2;
        src102 <= 16'h910;
        src103 <= 16'hfa8f;
        src104 <= 16'hc382;
        src105 <= 16'h217d;
        src106 <= 16'h5a13;
        src107 <= 16'h5c04;
        src108 <= 16'hd540;
        src109 <= 16'h89d2;
        src110 <= 16'h7943;
        src111 <= 16'hc838;
        src112 <= 16'hbc11;
        src113 <= 16'h568e;
        src114 <= 16'h84fb;
        src115 <= 16'hfd47;
        src116 <= 16'hb717;
        src117 <= 16'h36dd;
        src118 <= 16'h12eb;
        src119 <= 16'hfd8c;
        src120 <= 16'h4d67;
        src121 <= 16'h3965;
        src122 <= 16'h264f;
        src123 <= 16'h3982;
        src124 <= 16'h7f92;
        src125 <= 16'hda07;
        src126 <= 16'h4c50;
        src127 <= 16'he52f;
        src128 <= 16'h5079;
        src129 <= 16'hc80b;
        src130 <= 16'h3d42;
        src131 <= 16'h1a95;
        src132 <= 16'hda2e;
        src133 <= 16'h1eda;
        src134 <= 16'hc6d0;
        src135 <= 16'h84e;
        src136 <= 16'hfaf5;
        src137 <= 16'hccc;
        src138 <= 16'h2e5c;
        src139 <= 16'h1c3e;
        src140 <= 16'h311d;
        src141 <= 16'hc9c4;
        src142 <= 16'h915;
        src143 <= 16'h8e45;
        src144 <= 16'h2c74;
        src145 <= 16'h7727;
        src146 <= 16'h3dc2;
        src147 <= 16'h1671;
        src148 <= 16'h206b;
        src149 <= 16'h12c2;
        src150 <= 16'h228e;
        src151 <= 16'had88;
        src152 <= 16'hd9c8;
        src153 <= 16'h94a5;
        src154 <= 16'h4836;
        src155 <= 16'h88b7;
        src156 <= 16'h721f;
        src157 <= 16'h59a7;
        src158 <= 16'he893;
        src159 <= 16'h2447;
        src160 <= 16'hfea7;
        src161 <= 16'h903f;
        src162 <= 16'h31ce;
        src163 <= 16'h4541;
        src164 <= 16'he4bb;
        src165 <= 16'h85c5;
        src166 <= 16'h8ede;
        src167 <= 16'hb0c4;
        src168 <= 16'haa19;
        src169 <= 16'hb177;
        src170 <= 16'hea77;
        src171 <= 16'h36fa;
        src172 <= 16'h51cd;
        src173 <= 16'h18a;
        src174 <= 16'h78a5;
        src175 <= 16'hcd48;
        src176 <= 16'hd5ef;
        src177 <= 16'h33dd;
        src178 <= 16'h49f1;
        src179 <= 16'h78f3;
        src180 <= 16'h2f72;
        src181 <= 16'h5d11;
        src182 <= 16'h9568;
        src183 <= 16'hac62;
        src184 <= 16'hf6b1;
        exp <= 24'h58a997;
        #1
        src0 <= 16'h975d;
        src1 <= 16'he4a1;
        src2 <= 16'hb5a7;
        src3 <= 16'h901f;
        src4 <= 16'h85cb;
        src5 <= 16'h1a93;
        src6 <= 16'h33fc;
        src7 <= 16'hb85f;
        src8 <= 16'h6f28;
        src9 <= 16'ha744;
        src10 <= 16'hddb2;
        src11 <= 16'hbcf7;
        src12 <= 16'he05a;
        src13 <= 16'hf4bd;
        src14 <= 16'hbdea;
        src15 <= 16'haabe;
        src16 <= 16'h354;
        src17 <= 16'h166a;
        src18 <= 16'hcbcb;
        src19 <= 16'heed8;
        src20 <= 16'h9743;
        src21 <= 16'h36b;
        src22 <= 16'h7c8f;
        src23 <= 16'hf0c8;
        src24 <= 16'h7a62;
        src25 <= 16'h654c;
        src26 <= 16'h77d;
        src27 <= 16'h406e;
        src28 <= 16'hb17;
        src29 <= 16'h9874;
        src30 <= 16'h9d6b;
        src31 <= 16'h3b4b;
        src32 <= 16'h665;
        src33 <= 16'hed74;
        src34 <= 16'h3c0e;
        src35 <= 16'h3a39;
        src36 <= 16'hb5d3;
        src37 <= 16'hd532;
        src38 <= 16'hf5be;
        src39 <= 16'h1f94;
        src40 <= 16'hfddf;
        src41 <= 16'h32b6;
        src42 <= 16'h3211;
        src43 <= 16'h6da1;
        src44 <= 16'h6183;
        src45 <= 16'heb21;
        src46 <= 16'h96be;
        src47 <= 16'h1169;
        src48 <= 16'h9f2c;
        src49 <= 16'ha58e;
        src50 <= 16'he02d;
        src51 <= 16'h11c3;
        src52 <= 16'hf753;
        src53 <= 16'h5e59;
        src54 <= 16'hafb1;
        src55 <= 16'hc32a;
        src56 <= 16'h6e38;
        src57 <= 16'h6ab9;
        src58 <= 16'h6c8e;
        src59 <= 16'h9c2c;
        src60 <= 16'hb7d6;
        src61 <= 16'h6c21;
        src62 <= 16'h1a58;
        src63 <= 16'h4d27;
        src64 <= 16'h33f7;
        src65 <= 16'hed3a;
        src66 <= 16'h7942;
        src67 <= 16'h2d40;
        src68 <= 16'h45e8;
        src69 <= 16'hce58;
        src70 <= 16'h2874;
        src71 <= 16'he83a;
        src72 <= 16'hbf4f;
        src73 <= 16'h4f5;
        src74 <= 16'h1fcc;
        src75 <= 16'ha3be;
        src76 <= 16'h1710;
        src77 <= 16'ha0f9;
        src78 <= 16'h291a;
        src79 <= 16'he2ec;
        src80 <= 16'h3932;
        src81 <= 16'h4e07;
        src82 <= 16'h42be;
        src83 <= 16'h899b;
        src84 <= 16'hf04d;
        src85 <= 16'h9b5b;
        src86 <= 16'h512f;
        src87 <= 16'h2b3e;
        src88 <= 16'hafbd;
        src89 <= 16'hb8c0;
        src90 <= 16'hcc04;
        src91 <= 16'h17fb;
        src92 <= 16'h4ca8;
        src93 <= 16'hdb93;
        src94 <= 16'hb11c;
        src95 <= 16'h3b62;
        src96 <= 16'h21b;
        src97 <= 16'h297f;
        src98 <= 16'h1a2b;
        src99 <= 16'h5593;
        src100 <= 16'hbda1;
        src101 <= 16'h9db;
        src102 <= 16'h7ba0;
        src103 <= 16'hc3c0;
        src104 <= 16'h1ffe;
        src105 <= 16'h3cb2;
        src106 <= 16'h223;
        src107 <= 16'haad6;
        src108 <= 16'h7676;
        src109 <= 16'h74ba;
        src110 <= 16'h70ce;
        src111 <= 16'h8987;
        src112 <= 16'h5bdc;
        src113 <= 16'ha6fc;
        src114 <= 16'h2e8e;
        src115 <= 16'h29c1;
        src116 <= 16'h5ccb;
        src117 <= 16'hdc1c;
        src118 <= 16'h9f12;
        src119 <= 16'h408f;
        src120 <= 16'hac72;
        src121 <= 16'h1994;
        src122 <= 16'hde47;
        src123 <= 16'hd975;
        src124 <= 16'heca5;
        src125 <= 16'hfc22;
        src126 <= 16'hea27;
        src127 <= 16'hbea1;
        src128 <= 16'hfc66;
        src129 <= 16'hbc87;
        src130 <= 16'h6e51;
        src131 <= 16'heb97;
        src132 <= 16'h1790;
        src133 <= 16'heb7;
        src134 <= 16'h3440;
        src135 <= 16'hf3ae;
        src136 <= 16'hfe49;
        src137 <= 16'h1384;
        src138 <= 16'h44b0;
        src139 <= 16'heb4b;
        src140 <= 16'h61ea;
        src141 <= 16'h9fbe;
        src142 <= 16'h252b;
        src143 <= 16'h3ccd;
        src144 <= 16'hc685;
        src145 <= 16'hed1e;
        src146 <= 16'h2a1d;
        src147 <= 16'h733e;
        src148 <= 16'heeb5;
        src149 <= 16'h41e4;
        src150 <= 16'hfe52;
        src151 <= 16'hf4b7;
        src152 <= 16'hae5c;
        src153 <= 16'h22db;
        src154 <= 16'hc6e9;
        src155 <= 16'hb772;
        src156 <= 16'haa0c;
        src157 <= 16'h9093;
        src158 <= 16'h295b;
        src159 <= 16'hc1ec;
        src160 <= 16'ha29d;
        src161 <= 16'h1cc0;
        src162 <= 16'hae80;
        src163 <= 16'h8757;
        src164 <= 16'hd160;
        src165 <= 16'h132e;
        src166 <= 16'h5018;
        src167 <= 16'h5502;
        src168 <= 16'hfcc;
        src169 <= 16'h7865;
        src170 <= 16'h439b;
        src171 <= 16'h2212;
        src172 <= 16'h7e61;
        src173 <= 16'hc877;
        src174 <= 16'h7b8e;
        src175 <= 16'hedc;
        src176 <= 16'h75e6;
        src177 <= 16'hbf4b;
        src178 <= 16'h7575;
        src179 <= 16'h5780;
        src180 <= 16'ha811;
        src181 <= 16'h607a;
        src182 <= 16'h370d;
        src183 <= 16'he1d4;
        src184 <= 16'h8f55;
        exp <= 24'h5be495;
        #1
        src0 <= 16'h8656;
        src1 <= 16'h8718;
        src2 <= 16'h855c;
        src3 <= 16'hc1ae;
        src4 <= 16'h5cc5;
        src5 <= 16'h6593;
        src6 <= 16'h8022;
        src7 <= 16'hf59d;
        src8 <= 16'h21a8;
        src9 <= 16'h3369;
        src10 <= 16'hb81a;
        src11 <= 16'hc7;
        src12 <= 16'hd7ad;
        src13 <= 16'hc89c;
        src14 <= 16'ha7fb;
        src15 <= 16'heec2;
        src16 <= 16'hbc1e;
        src17 <= 16'hca06;
        src18 <= 16'h920e;
        src19 <= 16'h1283;
        src20 <= 16'h2c28;
        src21 <= 16'h300c;
        src22 <= 16'he127;
        src23 <= 16'hcaf7;
        src24 <= 16'h5bb9;
        src25 <= 16'h83f5;
        src26 <= 16'h6452;
        src27 <= 16'h9a6e;
        src28 <= 16'h303e;
        src29 <= 16'hbd2f;
        src30 <= 16'h7d49;
        src31 <= 16'h8b88;
        src32 <= 16'h1a9b;
        src33 <= 16'h5be5;
        src34 <= 16'hcd8f;
        src35 <= 16'h26de;
        src36 <= 16'ha37c;
        src37 <= 16'h7c54;
        src38 <= 16'h9af;
        src39 <= 16'h8463;
        src40 <= 16'h8a84;
        src41 <= 16'hf6a;
        src42 <= 16'h952c;
        src43 <= 16'hb493;
        src44 <= 16'h9ddf;
        src45 <= 16'h6e22;
        src46 <= 16'hbae8;
        src47 <= 16'hf9ed;
        src48 <= 16'h5213;
        src49 <= 16'h785d;
        src50 <= 16'h66fe;
        src51 <= 16'hd8;
        src52 <= 16'h7750;
        src53 <= 16'h3ab8;
        src54 <= 16'h9a85;
        src55 <= 16'h8309;
        src56 <= 16'h8a2a;
        src57 <= 16'h7ebb;
        src58 <= 16'h5346;
        src59 <= 16'hd8f9;
        src60 <= 16'hbc5a;
        src61 <= 16'h3c73;
        src62 <= 16'h6966;
        src63 <= 16'h2d70;
        src64 <= 16'h805e;
        src65 <= 16'h94;
        src66 <= 16'h739e;
        src67 <= 16'hcb21;
        src68 <= 16'hee0d;
        src69 <= 16'hd7e7;
        src70 <= 16'h4288;
        src71 <= 16'hf44f;
        src72 <= 16'he07f;
        src73 <= 16'h3dac;
        src74 <= 16'h46b5;
        src75 <= 16'h47c8;
        src76 <= 16'hb7d5;
        src77 <= 16'h730c;
        src78 <= 16'had07;
        src79 <= 16'he03a;
        src80 <= 16'he254;
        src81 <= 16'hc1c9;
        src82 <= 16'h560d;
        src83 <= 16'hfdbb;
        src84 <= 16'h751c;
        src85 <= 16'hfddb;
        src86 <= 16'h8935;
        src87 <= 16'h80ea;
        src88 <= 16'h36ef;
        src89 <= 16'h9622;
        src90 <= 16'hcfee;
        src91 <= 16'hc3c6;
        src92 <= 16'he6d3;
        src93 <= 16'h11c1;
        src94 <= 16'hb078;
        src95 <= 16'h3826;
        src96 <= 16'h8f86;
        src97 <= 16'hed38;
        src98 <= 16'hbbde;
        src99 <= 16'hbd72;
        src100 <= 16'h7c22;
        src101 <= 16'h6152;
        src102 <= 16'hbb2d;
        src103 <= 16'h9524;
        src104 <= 16'hc803;
        src105 <= 16'ha9d3;
        src106 <= 16'hfd6a;
        src107 <= 16'h4945;
        src108 <= 16'hbd02;
        src109 <= 16'haf29;
        src110 <= 16'hbfc5;
        src111 <= 16'h38f8;
        src112 <= 16'hf249;
        src113 <= 16'hab05;
        src114 <= 16'h7dc2;
        src115 <= 16'h50f1;
        src116 <= 16'h2db;
        src117 <= 16'h6091;
        src118 <= 16'hbf2f;
        src119 <= 16'h9b11;
        src120 <= 16'hcbf;
        src121 <= 16'h524;
        src122 <= 16'h325b;
        src123 <= 16'hb406;
        src124 <= 16'h3217;
        src125 <= 16'h144;
        src126 <= 16'hf538;
        src127 <= 16'ha4fc;
        src128 <= 16'h6786;
        src129 <= 16'h934f;
        src130 <= 16'h19c1;
        src131 <= 16'hecc1;
        src132 <= 16'hb9a1;
        src133 <= 16'h4c78;
        src134 <= 16'h2214;
        src135 <= 16'h4285;
        src136 <= 16'h4f01;
        src137 <= 16'h506f;
        src138 <= 16'h8110;
        src139 <= 16'h2c53;
        src140 <= 16'hb55b;
        src141 <= 16'h5522;
        src142 <= 16'h235a;
        src143 <= 16'h3c3;
        src144 <= 16'h7af1;
        src145 <= 16'h1f34;
        src146 <= 16'hbb70;
        src147 <= 16'h32ba;
        src148 <= 16'h9e61;
        src149 <= 16'h6d8f;
        src150 <= 16'hc838;
        src151 <= 16'h14b5;
        src152 <= 16'hac7c;
        src153 <= 16'h9710;
        src154 <= 16'h6e49;
        src155 <= 16'h59e8;
        src156 <= 16'hc9ed;
        src157 <= 16'h4a62;
        src158 <= 16'h3a04;
        src159 <= 16'he9d8;
        src160 <= 16'h600b;
        src161 <= 16'hc6ae;
        src162 <= 16'h151d;
        src163 <= 16'ha954;
        src164 <= 16'h163c;
        src165 <= 16'h9f37;
        src166 <= 16'h23cd;
        src167 <= 16'h727;
        src168 <= 16'h24f8;
        src169 <= 16'h1140;
        src170 <= 16'h4fcf;
        src171 <= 16'h3162;
        src172 <= 16'h9b9;
        src173 <= 16'haf40;
        src174 <= 16'h4943;
        src175 <= 16'hd601;
        src176 <= 16'h9563;
        src177 <= 16'hddd6;
        src178 <= 16'hdc07;
        src179 <= 16'hef5d;
        src180 <= 16'h4e39;
        src181 <= 16'hc62c;
        src182 <= 16'h23cb;
        src183 <= 16'h6545;
        src184 <= 16'hc736;
        exp <= 24'h5bfe30;
        #1
        src0 <= 16'hceb;
        src1 <= 16'hc5a5;
        src2 <= 16'hb940;
        src3 <= 16'h4492;
        src4 <= 16'hd378;
        src5 <= 16'h673d;
        src6 <= 16'h4108;
        src7 <= 16'hee74;
        src8 <= 16'h8885;
        src9 <= 16'hf51;
        src10 <= 16'h4e18;
        src11 <= 16'h5578;
        src12 <= 16'h2b4a;
        src13 <= 16'hae6b;
        src14 <= 16'h53b4;
        src15 <= 16'hd3b5;
        src16 <= 16'h91f7;
        src17 <= 16'hcd70;
        src18 <= 16'hd740;
        src19 <= 16'h5800;
        src20 <= 16'h4e19;
        src21 <= 16'hf049;
        src22 <= 16'hc63d;
        src23 <= 16'h7177;
        src24 <= 16'hd049;
        src25 <= 16'h9c24;
        src26 <= 16'h4790;
        src27 <= 16'hef6d;
        src28 <= 16'he7e6;
        src29 <= 16'hbc14;
        src30 <= 16'h91cd;
        src31 <= 16'ha955;
        src32 <= 16'hc4f0;
        src33 <= 16'h73fe;
        src34 <= 16'h749f;
        src35 <= 16'h6d9c;
        src36 <= 16'h283b;
        src37 <= 16'h991e;
        src38 <= 16'h6d10;
        src39 <= 16'hbe3a;
        src40 <= 16'h15c3;
        src41 <= 16'h98a4;
        src42 <= 16'h1ce9;
        src43 <= 16'h6536;
        src44 <= 16'h18a9;
        src45 <= 16'h7b7d;
        src46 <= 16'ha063;
        src47 <= 16'h3db1;
        src48 <= 16'hc6dc;
        src49 <= 16'h4641;
        src50 <= 16'h3d69;
        src51 <= 16'h7d32;
        src52 <= 16'h1286;
        src53 <= 16'h25c0;
        src54 <= 16'h60ef;
        src55 <= 16'h845a;
        src56 <= 16'hc667;
        src57 <= 16'hae0c;
        src58 <= 16'h4ba6;
        src59 <= 16'h5ee9;
        src60 <= 16'h256c;
        src61 <= 16'ha8ef;
        src62 <= 16'h4c7f;
        src63 <= 16'h9739;
        src64 <= 16'h2894;
        src65 <= 16'hcbfd;
        src66 <= 16'h15da;
        src67 <= 16'hf9fa;
        src68 <= 16'h975e;
        src69 <= 16'h4e83;
        src70 <= 16'hb87f;
        src71 <= 16'h733e;
        src72 <= 16'hf29;
        src73 <= 16'hf910;
        src74 <= 16'h8728;
        src75 <= 16'hb7f7;
        src76 <= 16'he698;
        src77 <= 16'he273;
        src78 <= 16'ha00a;
        src79 <= 16'h8ff1;
        src80 <= 16'hae3e;
        src81 <= 16'h5de7;
        src82 <= 16'h72f1;
        src83 <= 16'h87c0;
        src84 <= 16'h82e;
        src85 <= 16'h6bb1;
        src86 <= 16'h5f68;
        src87 <= 16'h5cfb;
        src88 <= 16'h6ce7;
        src89 <= 16'h5108;
        src90 <= 16'hedfc;
        src91 <= 16'h59ba;
        src92 <= 16'h3d40;
        src93 <= 16'hdf0b;
        src94 <= 16'h96b5;
        src95 <= 16'hada2;
        src96 <= 16'h12a7;
        src97 <= 16'ha27a;
        src98 <= 16'hfcc6;
        src99 <= 16'hdcc5;
        src100 <= 16'h4aff;
        src101 <= 16'h1efc;
        src102 <= 16'he3da;
        src103 <= 16'h45e7;
        src104 <= 16'hb2c;
        src105 <= 16'hf397;
        src106 <= 16'h2c20;
        src107 <= 16'h2c97;
        src108 <= 16'h807d;
        src109 <= 16'h47e7;
        src110 <= 16'hcd7;
        src111 <= 16'hadad;
        src112 <= 16'h925b;
        src113 <= 16'hd165;
        src114 <= 16'hce6b;
        src115 <= 16'ha7c;
        src116 <= 16'h9ef4;
        src117 <= 16'h9a72;
        src118 <= 16'h75cd;
        src119 <= 16'h57b;
        src120 <= 16'h4cb4;
        src121 <= 16'hb7a7;
        src122 <= 16'h74cc;
        src123 <= 16'h2392;
        src124 <= 16'hdf79;
        src125 <= 16'hee56;
        src126 <= 16'h8f7b;
        src127 <= 16'hecbf;
        src128 <= 16'h2744;
        src129 <= 16'hc1bb;
        src130 <= 16'hea1c;
        src131 <= 16'h40ea;
        src132 <= 16'h2046;
        src133 <= 16'h9521;
        src134 <= 16'h86a1;
        src135 <= 16'h2ae7;
        src136 <= 16'h23a0;
        src137 <= 16'h9379;
        src138 <= 16'hd968;
        src139 <= 16'hf3db;
        src140 <= 16'h6ee8;
        src141 <= 16'h141c;
        src142 <= 16'hfb50;
        src143 <= 16'ha535;
        src144 <= 16'h50b0;
        src145 <= 16'h9dd3;
        src146 <= 16'h2512;
        src147 <= 16'h2c89;
        src148 <= 16'he1ec;
        src149 <= 16'ha5c3;
        src150 <= 16'hbcf1;
        src151 <= 16'h283e;
        src152 <= 16'hc09f;
        src153 <= 16'ha823;
        src154 <= 16'h3f1c;
        src155 <= 16'h3a58;
        src156 <= 16'hde40;
        src157 <= 16'hccb0;
        src158 <= 16'hb1b2;
        src159 <= 16'h2d6e;
        src160 <= 16'h4a05;
        src161 <= 16'h8202;
        src162 <= 16'h3f63;
        src163 <= 16'h7c91;
        src164 <= 16'hbc0a;
        src165 <= 16'hf301;
        src166 <= 16'hf4da;
        src167 <= 16'h169b;
        src168 <= 16'he799;
        src169 <= 16'h6039;
        src170 <= 16'h3f48;
        src171 <= 16'h150a;
        src172 <= 16'h4f56;
        src173 <= 16'hb41c;
        src174 <= 16'h90a5;
        src175 <= 16'h8496;
        src176 <= 16'h45fb;
        src177 <= 16'h428a;
        src178 <= 16'hee4f;
        src179 <= 16'hee62;
        src180 <= 16'h8ce6;
        src181 <= 16'hfb83;
        src182 <= 16'h9ec2;
        src183 <= 16'h121f;
        src184 <= 16'hb26e;
        exp <= 24'h5dac38;
        #1
        src0 <= 16'hc28b;
        src1 <= 16'hb693;
        src2 <= 16'haf6a;
        src3 <= 16'h37db;
        src4 <= 16'h9b05;
        src5 <= 16'he841;
        src6 <= 16'heed;
        src7 <= 16'hdfc7;
        src8 <= 16'hbeec;
        src9 <= 16'h7f5c;
        src10 <= 16'hd6d8;
        src11 <= 16'hcebb;
        src12 <= 16'h9589;
        src13 <= 16'ha149;
        src14 <= 16'h7f46;
        src15 <= 16'he773;
        src16 <= 16'hc95;
        src17 <= 16'hc914;
        src18 <= 16'h6bdf;
        src19 <= 16'h7a22;
        src20 <= 16'h818d;
        src21 <= 16'hf38;
        src22 <= 16'he237;
        src23 <= 16'hbf28;
        src24 <= 16'h93e2;
        src25 <= 16'hdf9e;
        src26 <= 16'h18a7;
        src27 <= 16'hf4d9;
        src28 <= 16'h84c9;
        src29 <= 16'h64f5;
        src30 <= 16'h6ab0;
        src31 <= 16'hcf54;
        src32 <= 16'haf36;
        src33 <= 16'h6dcf;
        src34 <= 16'h4513;
        src35 <= 16'h499b;
        src36 <= 16'h63cb;
        src37 <= 16'h90f6;
        src38 <= 16'h16a8;
        src39 <= 16'h7694;
        src40 <= 16'h984;
        src41 <= 16'h1f0d;
        src42 <= 16'hba7e;
        src43 <= 16'h29b3;
        src44 <= 16'h52a5;
        src45 <= 16'h57e7;
        src46 <= 16'ha6a7;
        src47 <= 16'hd7d6;
        src48 <= 16'hb650;
        src49 <= 16'hff97;
        src50 <= 16'hc0f5;
        src51 <= 16'h7115;
        src52 <= 16'hf7d9;
        src53 <= 16'hb283;
        src54 <= 16'hdfa6;
        src55 <= 16'h817a;
        src56 <= 16'h1d00;
        src57 <= 16'h13bb;
        src58 <= 16'h8c0f;
        src59 <= 16'h523;
        src60 <= 16'h405e;
        src61 <= 16'haa83;
        src62 <= 16'hec5c;
        src63 <= 16'h4824;
        src64 <= 16'h247;
        src65 <= 16'h51d2;
        src66 <= 16'h2321;
        src67 <= 16'h8e64;
        src68 <= 16'h639b;
        src69 <= 16'hf3eb;
        src70 <= 16'h2dfc;
        src71 <= 16'h9bd5;
        src72 <= 16'h1fd2;
        src73 <= 16'h75d;
        src74 <= 16'h444;
        src75 <= 16'h67ee;
        src76 <= 16'h9741;
        src77 <= 16'h4a14;
        src78 <= 16'h3159;
        src79 <= 16'hebce;
        src80 <= 16'hd5c6;
        src81 <= 16'hd13e;
        src82 <= 16'h297e;
        src83 <= 16'h5ae5;
        src84 <= 16'h44dd;
        src85 <= 16'h7b24;
        src86 <= 16'h8f64;
        src87 <= 16'h463e;
        src88 <= 16'h81f3;
        src89 <= 16'hd7f0;
        src90 <= 16'h9a5a;
        src91 <= 16'h55bf;
        src92 <= 16'h8bdd;
        src93 <= 16'h665f;
        src94 <= 16'h28ee;
        src95 <= 16'h44a5;
        src96 <= 16'h152;
        src97 <= 16'h396b;
        src98 <= 16'hf3f9;
        src99 <= 16'h8fff;
        src100 <= 16'hae26;
        src101 <= 16'h64fa;
        src102 <= 16'h9506;
        src103 <= 16'hb4f3;
        src104 <= 16'hd00;
        src105 <= 16'hc04e;
        src106 <= 16'h67b1;
        src107 <= 16'h305c;
        src108 <= 16'h327b;
        src109 <= 16'h8bd3;
        src110 <= 16'ha4a3;
        src111 <= 16'h556;
        src112 <= 16'h459f;
        src113 <= 16'h7df;
        src114 <= 16'h5f23;
        src115 <= 16'h7377;
        src116 <= 16'h3e9e;
        src117 <= 16'hadf9;
        src118 <= 16'h3f61;
        src119 <= 16'hce7f;
        src120 <= 16'h89e3;
        src121 <= 16'h8c45;
        src122 <= 16'he9b6;
        src123 <= 16'hc55b;
        src124 <= 16'h8873;
        src125 <= 16'hcd1b;
        src126 <= 16'h89cf;
        src127 <= 16'hfced;
        src128 <= 16'hc22e;
        src129 <= 16'h4f1;
        src130 <= 16'h3ae4;
        src131 <= 16'hda20;
        src132 <= 16'h53e1;
        src133 <= 16'h3d93;
        src134 <= 16'h1db0;
        src135 <= 16'hc868;
        src136 <= 16'h1c9;
        src137 <= 16'h2ea7;
        src138 <= 16'h29c0;
        src139 <= 16'h3af4;
        src140 <= 16'hfa5;
        src141 <= 16'h4907;
        src142 <= 16'h746f;
        src143 <= 16'h2529;
        src144 <= 16'hb027;
        src145 <= 16'hea85;
        src146 <= 16'h6cc8;
        src147 <= 16'hc01d;
        src148 <= 16'h95e5;
        src149 <= 16'hb88f;
        src150 <= 16'hdde6;
        src151 <= 16'h426f;
        src152 <= 16'h9f83;
        src153 <= 16'h7e56;
        src154 <= 16'h1cf0;
        src155 <= 16'h86d8;
        src156 <= 16'h4d1b;
        src157 <= 16'h2d8;
        src158 <= 16'h12ac;
        src159 <= 16'hc367;
        src160 <= 16'h50e9;
        src161 <= 16'hd510;
        src162 <= 16'h511e;
        src163 <= 16'hfd51;
        src164 <= 16'h8e9b;
        src165 <= 16'hdce8;
        src166 <= 16'h187a;
        src167 <= 16'h138f;
        src168 <= 16'h6922;
        src169 <= 16'h7c03;
        src170 <= 16'hce6b;
        src171 <= 16'h57aa;
        src172 <= 16'h8276;
        src173 <= 16'h7cc4;
        src174 <= 16'h5187;
        src175 <= 16'hc151;
        src176 <= 16'hc01;
        src177 <= 16'h73ce;
        src178 <= 16'h745;
        src179 <= 16'h490c;
        src180 <= 16'hb0a5;
        src181 <= 16'h1b6a;
        src182 <= 16'hdd50;
        src183 <= 16'hb820;
        src184 <= 16'h9279;
        exp <= 24'h57ce22;
        #1
        src0 <= 16'h5f8e;
        src1 <= 16'hbec0;
        src2 <= 16'h149c;
        src3 <= 16'h474c;
        src4 <= 16'hf820;
        src5 <= 16'hc3b1;
        src6 <= 16'he063;
        src7 <= 16'h72e1;
        src8 <= 16'h8e19;
        src9 <= 16'h1b5f;
        src10 <= 16'h792e;
        src11 <= 16'hd916;
        src12 <= 16'hc1fc;
        src13 <= 16'h92f2;
        src14 <= 16'h6746;
        src15 <= 16'h5d69;
        src16 <= 16'hac88;
        src17 <= 16'ha32e;
        src18 <= 16'h6f0d;
        src19 <= 16'h675a;
        src20 <= 16'h69af;
        src21 <= 16'hd524;
        src22 <= 16'h5b19;
        src23 <= 16'h7469;
        src24 <= 16'hafc9;
        src25 <= 16'h30c9;
        src26 <= 16'h9315;
        src27 <= 16'h9e87;
        src28 <= 16'hebdb;
        src29 <= 16'hf13a;
        src30 <= 16'hf27a;
        src31 <= 16'ha1bc;
        src32 <= 16'had2c;
        src33 <= 16'hbde3;
        src34 <= 16'h7d77;
        src35 <= 16'h989d;
        src36 <= 16'ha50f;
        src37 <= 16'ha5d6;
        src38 <= 16'h6f5;
        src39 <= 16'ha039;
        src40 <= 16'hb21e;
        src41 <= 16'ha1f8;
        src42 <= 16'h4745;
        src43 <= 16'h5e81;
        src44 <= 16'h3652;
        src45 <= 16'h3fe8;
        src46 <= 16'h9727;
        src47 <= 16'h9d12;
        src48 <= 16'h6964;
        src49 <= 16'h345d;
        src50 <= 16'h2647;
        src51 <= 16'h4717;
        src52 <= 16'hee70;
        src53 <= 16'h1db5;
        src54 <= 16'hff96;
        src55 <= 16'h512c;
        src56 <= 16'h716f;
        src57 <= 16'hbad7;
        src58 <= 16'h97aa;
        src59 <= 16'h4ba;
        src60 <= 16'he852;
        src61 <= 16'h1696;
        src62 <= 16'h2bc2;
        src63 <= 16'h4aa;
        src64 <= 16'hd844;
        src65 <= 16'ha47d;
        src66 <= 16'h88e6;
        src67 <= 16'he117;
        src68 <= 16'h1db4;
        src69 <= 16'h245c;
        src70 <= 16'h36f;
        src71 <= 16'ha183;
        src72 <= 16'hf65a;
        src73 <= 16'h5413;
        src74 <= 16'h1271;
        src75 <= 16'ha460;
        src76 <= 16'hbdd2;
        src77 <= 16'h507c;
        src78 <= 16'haa8d;
        src79 <= 16'hdae8;
        src80 <= 16'ha8f4;
        src81 <= 16'ha89d;
        src82 <= 16'hc4f1;
        src83 <= 16'h7961;
        src84 <= 16'h761b;
        src85 <= 16'h6821;
        src86 <= 16'h1aee;
        src87 <= 16'h480d;
        src88 <= 16'hc0fa;
        src89 <= 16'h2242;
        src90 <= 16'heae3;
        src91 <= 16'h4221;
        src92 <= 16'he7cb;
        src93 <= 16'h5f67;
        src94 <= 16'hc814;
        src95 <= 16'hccad;
        src96 <= 16'h8e5;
        src97 <= 16'h3987;
        src98 <= 16'h5ad7;
        src99 <= 16'h939;
        src100 <= 16'h84f8;
        src101 <= 16'h3424;
        src102 <= 16'h6734;
        src103 <= 16'h5134;
        src104 <= 16'h7c3c;
        src105 <= 16'ha3a5;
        src106 <= 16'ha96e;
        src107 <= 16'h377;
        src108 <= 16'hccbf;
        src109 <= 16'h1d26;
        src110 <= 16'h2f3a;
        src111 <= 16'h45bc;
        src112 <= 16'h2409;
        src113 <= 16'hce59;
        src114 <= 16'h4d3d;
        src115 <= 16'h6ee3;
        src116 <= 16'h5df9;
        src117 <= 16'h75e5;
        src118 <= 16'hb80;
        src119 <= 16'hf452;
        src120 <= 16'hfcc;
        src121 <= 16'h5e47;
        src122 <= 16'ha096;
        src123 <= 16'h582e;
        src124 <= 16'hc11b;
        src125 <= 16'h5cd8;
        src126 <= 16'h33ac;
        src127 <= 16'hd7c3;
        src128 <= 16'h7e73;
        src129 <= 16'h5344;
        src130 <= 16'h4d3a;
        src131 <= 16'h90ac;
        src132 <= 16'hb8e8;
        src133 <= 16'hed84;
        src134 <= 16'h944c;
        src135 <= 16'h931e;
        src136 <= 16'h991a;
        src137 <= 16'h4f5d;
        src138 <= 16'h8468;
        src139 <= 16'h9cf9;
        src140 <= 16'hd0e9;
        src141 <= 16'hc92b;
        src142 <= 16'hf8d1;
        src143 <= 16'hb50b;
        src144 <= 16'hb2d6;
        src145 <= 16'h8f1d;
        src146 <= 16'hc5b0;
        src147 <= 16'h7646;
        src148 <= 16'h2fde;
        src149 <= 16'h3c5c;
        src150 <= 16'h6a4;
        src151 <= 16'ha163;
        src152 <= 16'hc222;
        src153 <= 16'he423;
        src154 <= 16'h4487;
        src155 <= 16'h64b5;
        src156 <= 16'h801a;
        src157 <= 16'hce21;
        src158 <= 16'he35b;
        src159 <= 16'hec69;
        src160 <= 16'h8541;
        src161 <= 16'heb36;
        src162 <= 16'hc6eb;
        src163 <= 16'ha6e7;
        src164 <= 16'hef64;
        src165 <= 16'h2d68;
        src166 <= 16'hbaf4;
        src167 <= 16'hb413;
        src168 <= 16'h3f45;
        src169 <= 16'h66a8;
        src170 <= 16'h2e6d;
        src171 <= 16'h15bc;
        src172 <= 16'h1a7a;
        src173 <= 16'h96ae;
        src174 <= 16'h6f50;
        src175 <= 16'hb9;
        src176 <= 16'hf3ba;
        src177 <= 16'h4c30;
        src178 <= 16'h11e4;
        src179 <= 16'hbba6;
        src180 <= 16'h6df7;
        src181 <= 16'hfd7;
        src182 <= 16'hd5e6;
        src183 <= 16'hf13b;
        src184 <= 16'ha905;
        exp <= 24'h5d83e2;
        #1
        src0 <= 16'h4bb9;
        src1 <= 16'h265c;
        src2 <= 16'h710f;
        src3 <= 16'h1edd;
        src4 <= 16'h7046;
        src5 <= 16'hb945;
        src6 <= 16'h775c;
        src7 <= 16'ha303;
        src8 <= 16'hbe81;
        src9 <= 16'h727;
        src10 <= 16'hc11;
        src11 <= 16'h8058;
        src12 <= 16'h3b91;
        src13 <= 16'h8543;
        src14 <= 16'hb45;
        src15 <= 16'h7be7;
        src16 <= 16'hec54;
        src17 <= 16'h75ed;
        src18 <= 16'hb2d4;
        src19 <= 16'h9a6d;
        src20 <= 16'h69d9;
        src21 <= 16'hd0da;
        src22 <= 16'h8511;
        src23 <= 16'hfe1e;
        src24 <= 16'he1d8;
        src25 <= 16'he3e4;
        src26 <= 16'h50db;
        src27 <= 16'h37c;
        src28 <= 16'hb865;
        src29 <= 16'h20c2;
        src30 <= 16'h14ee;
        src31 <= 16'h6606;
        src32 <= 16'ha00b;
        src33 <= 16'hf58e;
        src34 <= 16'h87af;
        src35 <= 16'h41dd;
        src36 <= 16'h7786;
        src37 <= 16'he878;
        src38 <= 16'h359d;
        src39 <= 16'hb63f;
        src40 <= 16'h650f;
        src41 <= 16'ha9cd;
        src42 <= 16'hc855;
        src43 <= 16'h5db5;
        src44 <= 16'h5d74;
        src45 <= 16'h353f;
        src46 <= 16'h3f2f;
        src47 <= 16'ha21d;
        src48 <= 16'h7c2f;
        src49 <= 16'h644f;
        src50 <= 16'he405;
        src51 <= 16'h4af8;
        src52 <= 16'h6942;
        src53 <= 16'h2dfd;
        src54 <= 16'h2df7;
        src55 <= 16'hcd71;
        src56 <= 16'hb503;
        src57 <= 16'hb8db;
        src58 <= 16'h951d;
        src59 <= 16'ha383;
        src60 <= 16'hf0f4;
        src61 <= 16'h796a;
        src62 <= 16'h9055;
        src63 <= 16'h1bc9;
        src64 <= 16'h5d23;
        src65 <= 16'hbec8;
        src66 <= 16'h1381;
        src67 <= 16'hc513;
        src68 <= 16'h62e4;
        src69 <= 16'h2e94;
        src70 <= 16'hfca;
        src71 <= 16'h6772;
        src72 <= 16'hb37f;
        src73 <= 16'h46fb;
        src74 <= 16'h36c6;
        src75 <= 16'h4ac6;
        src76 <= 16'h190;
        src77 <= 16'h6dbc;
        src78 <= 16'h3220;
        src79 <= 16'h440;
        src80 <= 16'h76b4;
        src81 <= 16'hdf21;
        src82 <= 16'hf7ab;
        src83 <= 16'h1158;
        src84 <= 16'hd2ed;
        src85 <= 16'h82ef;
        src86 <= 16'hcffc;
        src87 <= 16'hfc1a;
        src88 <= 16'h4867;
        src89 <= 16'h13bb;
        src90 <= 16'ha2b3;
        src91 <= 16'h452;
        src92 <= 16'h1710;
        src93 <= 16'hccef;
        src94 <= 16'he9aa;
        src95 <= 16'hb217;
        src96 <= 16'h20cd;
        src97 <= 16'h28d5;
        src98 <= 16'hbf12;
        src99 <= 16'hc659;
        src100 <= 16'h462c;
        src101 <= 16'hb33d;
        src102 <= 16'h5f10;
        src103 <= 16'he380;
        src104 <= 16'h65ff;
        src105 <= 16'h24ad;
        src106 <= 16'h4879;
        src107 <= 16'h3141;
        src108 <= 16'h4e4f;
        src109 <= 16'hd195;
        src110 <= 16'habc6;
        src111 <= 16'h7523;
        src112 <= 16'hfd06;
        src113 <= 16'hd8ea;
        src114 <= 16'h3b68;
        src115 <= 16'h2d59;
        src116 <= 16'hecad;
        src117 <= 16'h78b2;
        src118 <= 16'hd4b5;
        src119 <= 16'h497c;
        src120 <= 16'h3c08;
        src121 <= 16'hdf1e;
        src122 <= 16'hee6d;
        src123 <= 16'hd2d9;
        src124 <= 16'hf182;
        src125 <= 16'hfd29;
        src126 <= 16'h89d0;
        src127 <= 16'h73c3;
        src128 <= 16'hb087;
        src129 <= 16'h3ae;
        src130 <= 16'h8346;
        src131 <= 16'hd572;
        src132 <= 16'hbf13;
        src133 <= 16'h1af7;
        src134 <= 16'h5add;
        src135 <= 16'hb2ea;
        src136 <= 16'h128f;
        src137 <= 16'hd78e;
        src138 <= 16'hdfee;
        src139 <= 16'ha227;
        src140 <= 16'hac18;
        src141 <= 16'hde1a;
        src142 <= 16'h876c;
        src143 <= 16'hd883;
        src144 <= 16'hb4c;
        src145 <= 16'h2886;
        src146 <= 16'ha177;
        src147 <= 16'hc564;
        src148 <= 16'haa2c;
        src149 <= 16'hfcb7;
        src150 <= 16'hbbd7;
        src151 <= 16'hae1d;
        src152 <= 16'hc75b;
        src153 <= 16'hf0c2;
        src154 <= 16'hd19b;
        src155 <= 16'h416f;
        src156 <= 16'h6265;
        src157 <= 16'hab4d;
        src158 <= 16'h4dc1;
        src159 <= 16'hf8e8;
        src160 <= 16'h9b0f;
        src161 <= 16'h5a82;
        src162 <= 16'he2a3;
        src163 <= 16'h669d;
        src164 <= 16'h4c36;
        src165 <= 16'hfd42;
        src166 <= 16'h3aa2;
        src167 <= 16'hbe28;
        src168 <= 16'h49fb;
        src169 <= 16'he5ce;
        src170 <= 16'h3e74;
        src171 <= 16'h3a83;
        src172 <= 16'h805e;
        src173 <= 16'hde80;
        src174 <= 16'ha58a;
        src175 <= 16'h3a17;
        src176 <= 16'hf55;
        src177 <= 16'ha19f;
        src178 <= 16'h14cd;
        src179 <= 16'haff0;
        src180 <= 16'h7905;
        src181 <= 16'h9a5;
        src182 <= 16'h2e44;
        src183 <= 16'h4c09;
        src184 <= 16'h3c5a;
        exp <= 24'h5d99b3;
        #1
        src0 <= 16'h1e83;
        src1 <= 16'hd7ba;
        src2 <= 16'h7696;
        src3 <= 16'h2a;
        src4 <= 16'h16c1;
        src5 <= 16'h5654;
        src6 <= 16'h54cd;
        src7 <= 16'h98eb;
        src8 <= 16'h7ec7;
        src9 <= 16'he27b;
        src10 <= 16'hfeb4;
        src11 <= 16'hb8b0;
        src12 <= 16'hb2fa;
        src13 <= 16'h8891;
        src14 <= 16'hdd5;
        src15 <= 16'hf2aa;
        src16 <= 16'hc7ae;
        src17 <= 16'hd5da;
        src18 <= 16'h9860;
        src19 <= 16'h914c;
        src20 <= 16'hf773;
        src21 <= 16'hbcc4;
        src22 <= 16'hcc6c;
        src23 <= 16'h32de;
        src24 <= 16'h6ace;
        src25 <= 16'h1e6d;
        src26 <= 16'heefd;
        src27 <= 16'h99fe;
        src28 <= 16'h82e;
        src29 <= 16'hb139;
        src30 <= 16'h5867;
        src31 <= 16'h7b2e;
        src32 <= 16'h9a1e;
        src33 <= 16'h9d52;
        src34 <= 16'hc97f;
        src35 <= 16'h1230;
        src36 <= 16'h6913;
        src37 <= 16'h1033;
        src38 <= 16'h6aa2;
        src39 <= 16'h2a54;
        src40 <= 16'h699a;
        src41 <= 16'h5126;
        src42 <= 16'h1732;
        src43 <= 16'h2155;
        src44 <= 16'hd153;
        src45 <= 16'h2877;
        src46 <= 16'heec7;
        src47 <= 16'h3b47;
        src48 <= 16'h65b5;
        src49 <= 16'h7b35;
        src50 <= 16'hd6ef;
        src51 <= 16'h10a9;
        src52 <= 16'h8fe8;
        src53 <= 16'hf087;
        src54 <= 16'h26;
        src55 <= 16'hdc2c;
        src56 <= 16'hba5a;
        src57 <= 16'h6491;
        src58 <= 16'hc0e5;
        src59 <= 16'hae0f;
        src60 <= 16'h77c5;
        src61 <= 16'hdc26;
        src62 <= 16'h4e0f;
        src63 <= 16'h2623;
        src64 <= 16'hdc2a;
        src65 <= 16'hb149;
        src66 <= 16'habe8;
        src67 <= 16'h457;
        src68 <= 16'h4b89;
        src69 <= 16'h95e7;
        src70 <= 16'h360a;
        src71 <= 16'hae47;
        src72 <= 16'hb8d;
        src73 <= 16'h80e8;
        src74 <= 16'hf31b;
        src75 <= 16'h2642;
        src76 <= 16'h7935;
        src77 <= 16'h9a05;
        src78 <= 16'hb472;
        src79 <= 16'hf8f0;
        src80 <= 16'hc8ab;
        src81 <= 16'h74b9;
        src82 <= 16'haa24;
        src83 <= 16'h6d;
        src84 <= 16'h4ab7;
        src85 <= 16'hdf22;
        src86 <= 16'h3d12;
        src87 <= 16'h82a3;
        src88 <= 16'h7c23;
        src89 <= 16'h7db6;
        src90 <= 16'h1995;
        src91 <= 16'h7014;
        src92 <= 16'h4ced;
        src93 <= 16'h4ba5;
        src94 <= 16'hd05d;
        src95 <= 16'ha228;
        src96 <= 16'hd6cf;
        src97 <= 16'h1bf2;
        src98 <= 16'hd7c5;
        src99 <= 16'h77da;
        src100 <= 16'h82ce;
        src101 <= 16'h8daa;
        src102 <= 16'h266e;
        src103 <= 16'ha005;
        src104 <= 16'h8401;
        src105 <= 16'h6610;
        src106 <= 16'hd097;
        src107 <= 16'h3a27;
        src108 <= 16'hb94e;
        src109 <= 16'hd49a;
        src110 <= 16'ha8b0;
        src111 <= 16'hcbed;
        src112 <= 16'hac4f;
        src113 <= 16'h1216;
        src114 <= 16'he8e7;
        src115 <= 16'h3fa0;
        src116 <= 16'hf8cb;
        src117 <= 16'h2a56;
        src118 <= 16'hff21;
        src119 <= 16'h785c;
        src120 <= 16'habe3;
        src121 <= 16'hb445;
        src122 <= 16'h6cb0;
        src123 <= 16'hd171;
        src124 <= 16'h650a;
        src125 <= 16'hecf2;
        src126 <= 16'hed4e;
        src127 <= 16'hc07a;
        src128 <= 16'h3679;
        src129 <= 16'hf15e;
        src130 <= 16'hee99;
        src131 <= 16'hfccf;
        src132 <= 16'hf46f;
        src133 <= 16'h4fb3;
        src134 <= 16'h69ee;
        src135 <= 16'h6bc2;
        src136 <= 16'h248d;
        src137 <= 16'hd829;
        src138 <= 16'hbeb5;
        src139 <= 16'hef3c;
        src140 <= 16'h82f0;
        src141 <= 16'h72e7;
        src142 <= 16'h5a74;
        src143 <= 16'h68ad;
        src144 <= 16'h1624;
        src145 <= 16'h26d6;
        src146 <= 16'h8b3d;
        src147 <= 16'h945d;
        src148 <= 16'h5666;
        src149 <= 16'hfa41;
        src150 <= 16'h567a;
        src151 <= 16'hf76f;
        src152 <= 16'h6c2a;
        src153 <= 16'hecfa;
        src154 <= 16'h368c;
        src155 <= 16'h7b6;
        src156 <= 16'hc9c5;
        src157 <= 16'h3a08;
        src158 <= 16'hd84a;
        src159 <= 16'he427;
        src160 <= 16'hce4;
        src161 <= 16'h9afc;
        src162 <= 16'hd190;
        src163 <= 16'h7121;
        src164 <= 16'hd261;
        src165 <= 16'h7db2;
        src166 <= 16'h2dea;
        src167 <= 16'ha00c;
        src168 <= 16'hb119;
        src169 <= 16'hd9c1;
        src170 <= 16'ha948;
        src171 <= 16'h1b2f;
        src172 <= 16'h9af3;
        src173 <= 16'h3bc3;
        src174 <= 16'h190a;
        src175 <= 16'he881;
        src176 <= 16'ha908;
        src177 <= 16'h256b;
        src178 <= 16'h758a;
        src179 <= 16'h3039;
        src180 <= 16'h10a3;
        src181 <= 16'h5d88;
        src182 <= 16'hc592;
        src183 <= 16'h2abe;
        src184 <= 16'h72f8;
        exp <= 24'h603d9a;
        #1
        src0 <= 16'h9ff7;
        src1 <= 16'hcde1;
        src2 <= 16'h1454;
        src3 <= 16'h13a1;
        src4 <= 16'hfb20;
        src5 <= 16'ha09e;
        src6 <= 16'he4c3;
        src7 <= 16'hb7b8;
        src8 <= 16'h840c;
        src9 <= 16'hadb4;
        src10 <= 16'h7c80;
        src11 <= 16'hc888;
        src12 <= 16'h64b1;
        src13 <= 16'h9969;
        src14 <= 16'h65fe;
        src15 <= 16'h84e6;
        src16 <= 16'he955;
        src17 <= 16'haa30;
        src18 <= 16'h9416;
        src19 <= 16'h346e;
        src20 <= 16'h792d;
        src21 <= 16'hd213;
        src22 <= 16'hd964;
        src23 <= 16'hfcb1;
        src24 <= 16'h10d;
        src25 <= 16'h1f6e;
        src26 <= 16'h8aa6;
        src27 <= 16'h8fa4;
        src28 <= 16'hdfe4;
        src29 <= 16'h75f1;
        src30 <= 16'hbc2c;
        src31 <= 16'he5a8;
        src32 <= 16'hc4e1;
        src33 <= 16'h394e;
        src34 <= 16'hb49e;
        src35 <= 16'h21dc;
        src36 <= 16'h7103;
        src37 <= 16'h72d6;
        src38 <= 16'ha0c4;
        src39 <= 16'hc428;
        src40 <= 16'h76aa;
        src41 <= 16'hde;
        src42 <= 16'hed08;
        src43 <= 16'hc20;
        src44 <= 16'h6d2f;
        src45 <= 16'h44ba;
        src46 <= 16'h906e;
        src47 <= 16'h70bc;
        src48 <= 16'h6f9e;
        src49 <= 16'hb0f1;
        src50 <= 16'h3464;
        src51 <= 16'h910a;
        src52 <= 16'h908a;
        src53 <= 16'h35cc;
        src54 <= 16'he582;
        src55 <= 16'h37ea;
        src56 <= 16'he2e3;
        src57 <= 16'h416d;
        src58 <= 16'ha4d1;
        src59 <= 16'h72b;
        src60 <= 16'h35e8;
        src61 <= 16'had73;
        src62 <= 16'h7855;
        src63 <= 16'h6ded;
        src64 <= 16'h5d8c;
        src65 <= 16'hc55a;
        src66 <= 16'h5de6;
        src67 <= 16'h7f80;
        src68 <= 16'h1a9b;
        src69 <= 16'h5fb1;
        src70 <= 16'h7dd0;
        src71 <= 16'h632a;
        src72 <= 16'ha403;
        src73 <= 16'h9fbe;
        src74 <= 16'h5bd5;
        src75 <= 16'h221d;
        src76 <= 16'h1f03;
        src77 <= 16'hd683;
        src78 <= 16'h51a8;
        src79 <= 16'he391;
        src80 <= 16'h4fca;
        src81 <= 16'hd28d;
        src82 <= 16'h54a1;
        src83 <= 16'h37ff;
        src84 <= 16'hfd73;
        src85 <= 16'h8852;
        src86 <= 16'h4b92;
        src87 <= 16'hf33e;
        src88 <= 16'h34f2;
        src89 <= 16'h1049;
        src90 <= 16'h43fa;
        src91 <= 16'haacb;
        src92 <= 16'h6738;
        src93 <= 16'h26ce;
        src94 <= 16'ha250;
        src95 <= 16'hc432;
        src96 <= 16'hc2f4;
        src97 <= 16'h9317;
        src98 <= 16'hcbd6;
        src99 <= 16'h4e7b;
        src100 <= 16'hb673;
        src101 <= 16'hb3d6;
        src102 <= 16'ha34;
        src103 <= 16'he1a0;
        src104 <= 16'h9a0e;
        src105 <= 16'hcabd;
        src106 <= 16'h9d6e;
        src107 <= 16'h5d8e;
        src108 <= 16'h32a5;
        src109 <= 16'ha6b0;
        src110 <= 16'h3741;
        src111 <= 16'h8878;
        src112 <= 16'h616d;
        src113 <= 16'h2165;
        src114 <= 16'hdf5a;
        src115 <= 16'h3fa0;
        src116 <= 16'ha4e1;
        src117 <= 16'hcf4d;
        src118 <= 16'hc3eb;
        src119 <= 16'he20a;
        src120 <= 16'heb5c;
        src121 <= 16'h2d11;
        src122 <= 16'hd9a1;
        src123 <= 16'h538f;
        src124 <= 16'h5f12;
        src125 <= 16'h8291;
        src126 <= 16'ha81;
        src127 <= 16'hbf0;
        src128 <= 16'ha6fa;
        src129 <= 16'h81e2;
        src130 <= 16'ha7e3;
        src131 <= 16'h4658;
        src132 <= 16'h14e4;
        src133 <= 16'hacd7;
        src134 <= 16'h3828;
        src135 <= 16'h6e41;
        src136 <= 16'ha8fd;
        src137 <= 16'hdc83;
        src138 <= 16'hc295;
        src139 <= 16'h4d57;
        src140 <= 16'h70e;
        src141 <= 16'ha1bb;
        src142 <= 16'he6e9;
        src143 <= 16'h7f5e;
        src144 <= 16'h8f19;
        src145 <= 16'h4618;
        src146 <= 16'h6088;
        src147 <= 16'h7e74;
        src148 <= 16'h5abc;
        src149 <= 16'he49d;
        src150 <= 16'h102a;
        src151 <= 16'hf02e;
        src152 <= 16'h160e;
        src153 <= 16'ha9f2;
        src154 <= 16'h7f5;
        src155 <= 16'h973b;
        src156 <= 16'h11c5;
        src157 <= 16'hc6dc;
        src158 <= 16'h57e6;
        src159 <= 16'h1386;
        src160 <= 16'h5bb1;
        src161 <= 16'hb34a;
        src162 <= 16'hd386;
        src163 <= 16'h7abb;
        src164 <= 16'h3ab5;
        src165 <= 16'h4984;
        src166 <= 16'hddf9;
        src167 <= 16'h52d2;
        src168 <= 16'he688;
        src169 <= 16'h2859;
        src170 <= 16'hf83d;
        src171 <= 16'hc96b;
        src172 <= 16'h899c;
        src173 <= 16'he51b;
        src174 <= 16'h6f0e;
        src175 <= 16'h843e;
        src176 <= 16'hccf5;
        src177 <= 16'hc0de;
        src178 <= 16'hfe38;
        src179 <= 16'h9660;
        src180 <= 16'ha88e;
        src181 <= 16'h8089;
        src182 <= 16'h3e87;
        src183 <= 16'h67a8;
        src184 <= 16'hab6f;
        exp <= 24'h5ebc35;
        #1
        src0 <= 16'hd924;
        src1 <= 16'ha201;
        src2 <= 16'h598d;
        src3 <= 16'ha659;
        src4 <= 16'ha738;
        src5 <= 16'hd7a7;
        src6 <= 16'h7b53;
        src7 <= 16'h186;
        src8 <= 16'hb79a;
        src9 <= 16'hf32b;
        src10 <= 16'hb546;
        src11 <= 16'h6758;
        src12 <= 16'h73f9;
        src13 <= 16'hdb38;
        src14 <= 16'h8f2c;
        src15 <= 16'hcd5e;
        src16 <= 16'h11f2;
        src17 <= 16'h5bf9;
        src18 <= 16'hc12d;
        src19 <= 16'h81af;
        src20 <= 16'h49ec;
        src21 <= 16'h3ccd;
        src22 <= 16'hbb50;
        src23 <= 16'hf9b;
        src24 <= 16'hfe70;
        src25 <= 16'h568c;
        src26 <= 16'ha647;
        src27 <= 16'h254a;
        src28 <= 16'hd33e;
        src29 <= 16'hc3d6;
        src30 <= 16'h57ac;
        src31 <= 16'h6035;
        src32 <= 16'h66f7;
        src33 <= 16'h9271;
        src34 <= 16'h5a89;
        src35 <= 16'hf97a;
        src36 <= 16'h9338;
        src37 <= 16'h5d8f;
        src38 <= 16'hf44b;
        src39 <= 16'hcc44;
        src40 <= 16'hcde8;
        src41 <= 16'hc512;
        src42 <= 16'ha945;
        src43 <= 16'he6c;
        src44 <= 16'h4eed;
        src45 <= 16'hfebe;
        src46 <= 16'h1447;
        src47 <= 16'h7215;
        src48 <= 16'h5ee0;
        src49 <= 16'h4e47;
        src50 <= 16'hb70d;
        src51 <= 16'hb086;
        src52 <= 16'h14c5;
        src53 <= 16'h9340;
        src54 <= 16'hd61d;
        src55 <= 16'h894a;
        src56 <= 16'h3d40;
        src57 <= 16'hbde5;
        src58 <= 16'h7439;
        src59 <= 16'h21c9;
        src60 <= 16'h51bb;
        src61 <= 16'h29a7;
        src62 <= 16'ha2fe;
        src63 <= 16'hb684;
        src64 <= 16'h54a5;
        src65 <= 16'he76b;
        src66 <= 16'hc89e;
        src67 <= 16'hfe1e;
        src68 <= 16'h653d;
        src69 <= 16'h227b;
        src70 <= 16'h785;
        src71 <= 16'h6ae7;
        src72 <= 16'h501f;
        src73 <= 16'h1e4;
        src74 <= 16'h926b;
        src75 <= 16'h7734;
        src76 <= 16'h45e8;
        src77 <= 16'h5878;
        src78 <= 16'h5e97;
        src79 <= 16'h76ed;
        src80 <= 16'h7b2f;
        src81 <= 16'h489c;
        src82 <= 16'h2c9c;
        src83 <= 16'h956e;
        src84 <= 16'hb625;
        src85 <= 16'he1d2;
        src86 <= 16'h338b;
        src87 <= 16'h7433;
        src88 <= 16'he1a2;
        src89 <= 16'ha42f;
        src90 <= 16'h59cf;
        src91 <= 16'hf420;
        src92 <= 16'h1975;
        src93 <= 16'h8973;
        src94 <= 16'h2380;
        src95 <= 16'ha78c;
        src96 <= 16'h5d4f;
        src97 <= 16'h83d2;
        src98 <= 16'h77d9;
        src99 <= 16'hfc8f;
        src100 <= 16'haf56;
        src101 <= 16'h9f9a;
        src102 <= 16'hf8d4;
        src103 <= 16'h63a5;
        src104 <= 16'h331f;
        src105 <= 16'hbb12;
        src106 <= 16'he2f0;
        src107 <= 16'h9dc;
        src108 <= 16'h1e8;
        src109 <= 16'hf791;
        src110 <= 16'ha5d5;
        src111 <= 16'h1b79;
        src112 <= 16'hd104;
        src113 <= 16'h8e2f;
        src114 <= 16'ha267;
        src115 <= 16'h676d;
        src116 <= 16'h9a88;
        src117 <= 16'h5d1;
        src118 <= 16'h4ec7;
        src119 <= 16'hd35e;
        src120 <= 16'h1027;
        src121 <= 16'h8dff;
        src122 <= 16'h1740;
        src123 <= 16'h8137;
        src124 <= 16'h2b72;
        src125 <= 16'hc358;
        src126 <= 16'h3422;
        src127 <= 16'hb331;
        src128 <= 16'h44e3;
        src129 <= 16'h6fc3;
        src130 <= 16'h891d;
        src131 <= 16'h2d9b;
        src132 <= 16'hb11d;
        src133 <= 16'hd16d;
        src134 <= 16'h329b;
        src135 <= 16'hee1d;
        src136 <= 16'h41cb;
        src137 <= 16'hac62;
        src138 <= 16'h136;
        src139 <= 16'h87c;
        src140 <= 16'ha959;
        src141 <= 16'h1fb6;
        src142 <= 16'h1569;
        src143 <= 16'hd59d;
        src144 <= 16'hdac;
        src145 <= 16'h53cb;
        src146 <= 16'hf60b;
        src147 <= 16'h48dd;
        src148 <= 16'h613f;
        src149 <= 16'h1db7;
        src150 <= 16'h9cde;
        src151 <= 16'h5baa;
        src152 <= 16'h9894;
        src153 <= 16'hd4ef;
        src154 <= 16'hd621;
        src155 <= 16'h627d;
        src156 <= 16'hab1a;
        src157 <= 16'ha9;
        src158 <= 16'h5d6c;
        src159 <= 16'h53c2;
        src160 <= 16'hdb89;
        src161 <= 16'hc391;
        src162 <= 16'h9bc6;
        src163 <= 16'ha335;
        src164 <= 16'hb521;
        src165 <= 16'ha06c;
        src166 <= 16'h3a2c;
        src167 <= 16'h897b;
        src168 <= 16'h3091;
        src169 <= 16'h9d69;
        src170 <= 16'h201a;
        src171 <= 16'h4e01;
        src172 <= 16'h68a;
        src173 <= 16'h6ac1;
        src174 <= 16'h412d;
        src175 <= 16'h4f21;
        src176 <= 16'he39f;
        src177 <= 16'hdd63;
        src178 <= 16'h803e;
        src179 <= 16'hda1f;
        src180 <= 16'hf868;
        src181 <= 16'h289e;
        src182 <= 16'h1cc2;
        src183 <= 16'h3434;
        src184 <= 16'ha282;
        exp <= 24'h5ad872;
        #1
        src0 <= 16'h9730;
        src1 <= 16'hd7d5;
        src2 <= 16'h4730;
        src3 <= 16'h59f2;
        src4 <= 16'h2952;
        src5 <= 16'hed8;
        src6 <= 16'hd602;
        src7 <= 16'hdc77;
        src8 <= 16'hfd53;
        src9 <= 16'h9cfe;
        src10 <= 16'h2981;
        src11 <= 16'he725;
        src12 <= 16'hd9bb;
        src13 <= 16'h8a5b;
        src14 <= 16'h9f7d;
        src15 <= 16'hdce;
        src16 <= 16'h4fb7;
        src17 <= 16'ha90b;
        src18 <= 16'h26d0;
        src19 <= 16'h9262;
        src20 <= 16'h55f3;
        src21 <= 16'hccec;
        src22 <= 16'haf5e;
        src23 <= 16'hb904;
        src24 <= 16'he069;
        src25 <= 16'hba10;
        src26 <= 16'h713a;
        src27 <= 16'ha976;
        src28 <= 16'h1bfd;
        src29 <= 16'h5691;
        src30 <= 16'hd4a;
        src31 <= 16'hd768;
        src32 <= 16'hd4fa;
        src33 <= 16'h6cb0;
        src34 <= 16'h15a7;
        src35 <= 16'h5045;
        src36 <= 16'h65da;
        src37 <= 16'h60bc;
        src38 <= 16'h6cd5;
        src39 <= 16'ha2b3;
        src40 <= 16'h8c35;
        src41 <= 16'h902b;
        src42 <= 16'he268;
        src43 <= 16'h7215;
        src44 <= 16'h2270;
        src45 <= 16'h4c99;
        src46 <= 16'hdd94;
        src47 <= 16'h34bb;
        src48 <= 16'h351f;
        src49 <= 16'hc492;
        src50 <= 16'hc4b6;
        src51 <= 16'h2716;
        src52 <= 16'h2c74;
        src53 <= 16'h41fa;
        src54 <= 16'h3a54;
        src55 <= 16'h271e;
        src56 <= 16'h917;
        src57 <= 16'hb596;
        src58 <= 16'h3e26;
        src59 <= 16'h339d;
        src60 <= 16'h8423;
        src61 <= 16'hb038;
        src62 <= 16'h66ca;
        src63 <= 16'h9cff;
        src64 <= 16'h3985;
        src65 <= 16'h7a56;
        src66 <= 16'h7888;
        src67 <= 16'hfb70;
        src68 <= 16'h17b7;
        src69 <= 16'h7509;
        src70 <= 16'hd725;
        src71 <= 16'ha292;
        src72 <= 16'h9b2c;
        src73 <= 16'h4ea5;
        src74 <= 16'haa2f;
        src75 <= 16'h73b1;
        src76 <= 16'h35ea;
        src77 <= 16'h4cc9;
        src78 <= 16'hb457;
        src79 <= 16'h1bf8;
        src80 <= 16'h1128;
        src81 <= 16'h6c49;
        src82 <= 16'h21cd;
        src83 <= 16'h484e;
        src84 <= 16'h4f80;
        src85 <= 16'h84d2;
        src86 <= 16'h23cc;
        src87 <= 16'h40c5;
        src88 <= 16'h92ce;
        src89 <= 16'hb3d4;
        src90 <= 16'he876;
        src91 <= 16'hbf37;
        src92 <= 16'hf70b;
        src93 <= 16'h77d3;
        src94 <= 16'ha9a3;
        src95 <= 16'h9a56;
        src96 <= 16'h9a39;
        src97 <= 16'hafd7;
        src98 <= 16'hc984;
        src99 <= 16'h8f64;
        src100 <= 16'h208e;
        src101 <= 16'ha494;
        src102 <= 16'h3852;
        src103 <= 16'hce8a;
        src104 <= 16'hfb9d;
        src105 <= 16'h15ee;
        src106 <= 16'he08b;
        src107 <= 16'hf5c6;
        src108 <= 16'h1314;
        src109 <= 16'h4add;
        src110 <= 16'hbadc;
        src111 <= 16'hc916;
        src112 <= 16'heae;
        src113 <= 16'h6582;
        src114 <= 16'hb8c3;
        src115 <= 16'hc5af;
        src116 <= 16'h6c96;
        src117 <= 16'h5126;
        src118 <= 16'hc890;
        src119 <= 16'hab82;
        src120 <= 16'h4350;
        src121 <= 16'h9a8b;
        src122 <= 16'h370e;
        src123 <= 16'hfe0b;
        src124 <= 16'h577c;
        src125 <= 16'h7c82;
        src126 <= 16'hcdde;
        src127 <= 16'h4317;
        src128 <= 16'h7971;
        src129 <= 16'h89c0;
        src130 <= 16'h2bf6;
        src131 <= 16'h498e;
        src132 <= 16'hfbaa;
        src133 <= 16'h7003;
        src134 <= 16'h836c;
        src135 <= 16'h6b54;
        src136 <= 16'h6328;
        src137 <= 16'hf66;
        src138 <= 16'hdefc;
        src139 <= 16'h66c9;
        src140 <= 16'hf86b;
        src141 <= 16'h44e9;
        src142 <= 16'h772c;
        src143 <= 16'h2e53;
        src144 <= 16'hb990;
        src145 <= 16'h39b7;
        src146 <= 16'h310;
        src147 <= 16'haef8;
        src148 <= 16'hc926;
        src149 <= 16'h7c28;
        src150 <= 16'hed0e;
        src151 <= 16'ha817;
        src152 <= 16'h3d92;
        src153 <= 16'hc582;
        src154 <= 16'h1179;
        src155 <= 16'h7896;
        src156 <= 16'h2616;
        src157 <= 16'h2b6d;
        src158 <= 16'hc76a;
        src159 <= 16'h1147;
        src160 <= 16'h833b;
        src161 <= 16'h2bd8;
        src162 <= 16'h35b1;
        src163 <= 16'h963;
        src164 <= 16'hf884;
        src165 <= 16'h484a;
        src166 <= 16'hf994;
        src167 <= 16'hf506;
        src168 <= 16'h17db;
        src169 <= 16'hb374;
        src170 <= 16'hba7b;
        src171 <= 16'he4a8;
        src172 <= 16'h5e20;
        src173 <= 16'hbec8;
        src174 <= 16'h6c1f;
        src175 <= 16'h547d;
        src176 <= 16'h9342;
        src177 <= 16'hb697;
        src178 <= 16'hfd08;
        src179 <= 16'hba87;
        src180 <= 16'h2f10;
        src181 <= 16'h583;
        src182 <= 16'h237a;
        src183 <= 16'h7d5;
        src184 <= 16'hf0ac;
        exp <= 24'h5a8b14;
        #1
        src0 <= 16'h421;
        src1 <= 16'h9936;
        src2 <= 16'h5fae;
        src3 <= 16'heef2;
        src4 <= 16'h147d;
        src5 <= 16'hb394;
        src6 <= 16'h2a36;
        src7 <= 16'ha65f;
        src8 <= 16'h47b7;
        src9 <= 16'h3ea5;
        src10 <= 16'ha907;
        src11 <= 16'hd640;
        src12 <= 16'he21e;
        src13 <= 16'h3e48;
        src14 <= 16'h99de;
        src15 <= 16'h75fa;
        src16 <= 16'hfc52;
        src17 <= 16'hb73c;
        src18 <= 16'h3449;
        src19 <= 16'heb90;
        src20 <= 16'hcce5;
        src21 <= 16'hf2bb;
        src22 <= 16'h4a37;
        src23 <= 16'h102d;
        src24 <= 16'hbf4d;
        src25 <= 16'h2d5b;
        src26 <= 16'h1d98;
        src27 <= 16'hf67d;
        src28 <= 16'haef9;
        src29 <= 16'hc4ff;
        src30 <= 16'h924d;
        src31 <= 16'h5b25;
        src32 <= 16'h18bd;
        src33 <= 16'h1ee3;
        src34 <= 16'h55c8;
        src35 <= 16'h668b;
        src36 <= 16'h68ae;
        src37 <= 16'head2;
        src38 <= 16'hdbf8;
        src39 <= 16'h64af;
        src40 <= 16'hfcfc;
        src41 <= 16'he31d;
        src42 <= 16'heed5;
        src43 <= 16'h9057;
        src44 <= 16'h6c91;
        src45 <= 16'h97f8;
        src46 <= 16'h9e78;
        src47 <= 16'h81f7;
        src48 <= 16'h22ad;
        src49 <= 16'h6ff8;
        src50 <= 16'h2358;
        src51 <= 16'h6168;
        src52 <= 16'h9fe8;
        src53 <= 16'hae16;
        src54 <= 16'he58b;
        src55 <= 16'h8f07;
        src56 <= 16'hb9d4;
        src57 <= 16'hbf16;
        src58 <= 16'he763;
        src59 <= 16'ha471;
        src60 <= 16'h199b;
        src61 <= 16'hf64b;
        src62 <= 16'h2f92;
        src63 <= 16'hef97;
        src64 <= 16'h425b;
        src65 <= 16'ha1e5;
        src66 <= 16'h7cb5;
        src67 <= 16'h2d0a;
        src68 <= 16'h974c;
        src69 <= 16'h56ab;
        src70 <= 16'h743c;
        src71 <= 16'h51d;
        src72 <= 16'h81f2;
        src73 <= 16'h89f5;
        src74 <= 16'h4601;
        src75 <= 16'hf0d5;
        src76 <= 16'h6e06;
        src77 <= 16'hdac;
        src78 <= 16'hdc08;
        src79 <= 16'h2078;
        src80 <= 16'h596e;
        src81 <= 16'h571;
        src82 <= 16'h7bea;
        src83 <= 16'h6c2d;
        src84 <= 16'hae6c;
        src85 <= 16'h5641;
        src86 <= 16'h89a2;
        src87 <= 16'h64cb;
        src88 <= 16'h84c3;
        src89 <= 16'he2fb;
        src90 <= 16'h4585;
        src91 <= 16'hbc2;
        src92 <= 16'h2f1a;
        src93 <= 16'hc321;
        src94 <= 16'hac17;
        src95 <= 16'h6b7d;
        src96 <= 16'hf91d;
        src97 <= 16'h3e03;
        src98 <= 16'hfdff;
        src99 <= 16'h57bd;
        src100 <= 16'h3aa;
        src101 <= 16'h1155;
        src102 <= 16'h6bbd;
        src103 <= 16'h257;
        src104 <= 16'hfdad;
        src105 <= 16'h9ff3;
        src106 <= 16'hf2e;
        src107 <= 16'h229b;
        src108 <= 16'h739c;
        src109 <= 16'h2b52;
        src110 <= 16'hf2af;
        src111 <= 16'h1822;
        src112 <= 16'h3bd3;
        src113 <= 16'h8fbd;
        src114 <= 16'h9439;
        src115 <= 16'h858;
        src116 <= 16'he7ad;
        src117 <= 16'h19d5;
        src118 <= 16'ha695;
        src119 <= 16'hacbe;
        src120 <= 16'h2c4c;
        src121 <= 16'h5a67;
        src122 <= 16'hbc09;
        src123 <= 16'hd7b8;
        src124 <= 16'hf2ed;
        src125 <= 16'hc51b;
        src126 <= 16'h8d14;
        src127 <= 16'h5079;
        src128 <= 16'h48ce;
        src129 <= 16'h9e8;
        src130 <= 16'he5b2;
        src131 <= 16'hb6c7;
        src132 <= 16'hf4b8;
        src133 <= 16'hb1a4;
        src134 <= 16'h54ca;
        src135 <= 16'hb16c;
        src136 <= 16'h1071;
        src137 <= 16'hf329;
        src138 <= 16'h897e;
        src139 <= 16'h873b;
        src140 <= 16'ha19f;
        src141 <= 16'h2bca;
        src142 <= 16'h39b9;
        src143 <= 16'h95cc;
        src144 <= 16'h11fe;
        src145 <= 16'hdf19;
        src146 <= 16'h45b9;
        src147 <= 16'he872;
        src148 <= 16'h4f2f;
        src149 <= 16'h3368;
        src150 <= 16'h1109;
        src151 <= 16'h5e6e;
        src152 <= 16'h42df;
        src153 <= 16'hf37c;
        src154 <= 16'ha017;
        src155 <= 16'h96b0;
        src156 <= 16'h42b2;
        src157 <= 16'hc8a;
        src158 <= 16'hff23;
        src159 <= 16'hdf82;
        src160 <= 16'hc44;
        src161 <= 16'he397;
        src162 <= 16'h3207;
        src163 <= 16'h43eb;
        src164 <= 16'h7a7d;
        src165 <= 16'h593b;
        src166 <= 16'h56ff;
        src167 <= 16'h1ac1;
        src168 <= 16'h5f14;
        src169 <= 16'ha723;
        src170 <= 16'h25dc;
        src171 <= 16'h63ae;
        src172 <= 16'h35db;
        src173 <= 16'hd2b;
        src174 <= 16'hbda6;
        src175 <= 16'hff9c;
        src176 <= 16'h3479;
        src177 <= 16'hda06;
        src178 <= 16'h251d;
        src179 <= 16'h59c2;
        src180 <= 16'h4a45;
        src181 <= 16'h4ffe;
        src182 <= 16'h310;
        src183 <= 16'h9444;
        src184 <= 16'h19ba;
        exp <= 24'h58d4b3;
        #1
        src0 <= 16'haaa3;
        src1 <= 16'h230b;
        src2 <= 16'h46e9;
        src3 <= 16'hd04d;
        src4 <= 16'hc48b;
        src5 <= 16'h9fb6;
        src6 <= 16'h2742;
        src7 <= 16'h4a37;
        src8 <= 16'h19fc;
        src9 <= 16'h246f;
        src10 <= 16'h2a40;
        src11 <= 16'h7df;
        src12 <= 16'h382b;
        src13 <= 16'h1cb3;
        src14 <= 16'h2fee;
        src15 <= 16'h6549;
        src16 <= 16'h7155;
        src17 <= 16'ha87f;
        src18 <= 16'h56a7;
        src19 <= 16'ha791;
        src20 <= 16'hf74d;
        src21 <= 16'h20c4;
        src22 <= 16'h5861;
        src23 <= 16'h5ba2;
        src24 <= 16'h285c;
        src25 <= 16'h2f5;
        src26 <= 16'h2cab;
        src27 <= 16'h69a6;
        src28 <= 16'hd316;
        src29 <= 16'hf9ad;
        src30 <= 16'h9ffb;
        src31 <= 16'h1566;
        src32 <= 16'h217b;
        src33 <= 16'hda5;
        src34 <= 16'ha72d;
        src35 <= 16'h7510;
        src36 <= 16'hb10e;
        src37 <= 16'h3d99;
        src38 <= 16'hc0e4;
        src39 <= 16'hf0c1;
        src40 <= 16'h90f8;
        src41 <= 16'h389f;
        src42 <= 16'hc84d;
        src43 <= 16'hbcf4;
        src44 <= 16'h6f3a;
        src45 <= 16'h688b;
        src46 <= 16'hc7ac;
        src47 <= 16'hcc5a;
        src48 <= 16'hc8c0;
        src49 <= 16'hb714;
        src50 <= 16'h2068;
        src51 <= 16'ha73a;
        src52 <= 16'h983f;
        src53 <= 16'h3358;
        src54 <= 16'h85c8;
        src55 <= 16'hfc8f;
        src56 <= 16'hb2cb;
        src57 <= 16'h9973;
        src58 <= 16'hc7e0;
        src59 <= 16'hf193;
        src60 <= 16'hbc75;
        src61 <= 16'h59b4;
        src62 <= 16'h4683;
        src63 <= 16'h3fbb;
        src64 <= 16'h10f9;
        src65 <= 16'hff28;
        src66 <= 16'ha99c;
        src67 <= 16'h61f0;
        src68 <= 16'h8d2f;
        src69 <= 16'h9479;
        src70 <= 16'hcdc2;
        src71 <= 16'h1d50;
        src72 <= 16'he2da;
        src73 <= 16'h9a5d;
        src74 <= 16'he569;
        src75 <= 16'h7790;
        src76 <= 16'h33f3;
        src77 <= 16'hfa70;
        src78 <= 16'h73f7;
        src79 <= 16'h5c83;
        src80 <= 16'hbfb9;
        src81 <= 16'hf902;
        src82 <= 16'hc6b7;
        src83 <= 16'h7cc3;
        src84 <= 16'hdadf;
        src85 <= 16'h579e;
        src86 <= 16'hee;
        src87 <= 16'hb65b;
        src88 <= 16'h3517;
        src89 <= 16'h7477;
        src90 <= 16'h65cc;
        src91 <= 16'h6852;
        src92 <= 16'h117;
        src93 <= 16'h3e01;
        src94 <= 16'h66a2;
        src95 <= 16'ha39c;
        src96 <= 16'h197;
        src97 <= 16'hdc29;
        src98 <= 16'ha0a8;
        src99 <= 16'ha913;
        src100 <= 16'h5b65;
        src101 <= 16'h3967;
        src102 <= 16'h57a9;
        src103 <= 16'hd5ad;
        src104 <= 16'h6be8;
        src105 <= 16'h78f3;
        src106 <= 16'h72f5;
        src107 <= 16'h498e;
        src108 <= 16'h5466;
        src109 <= 16'h8bc3;
        src110 <= 16'h47c5;
        src111 <= 16'hb0ed;
        src112 <= 16'he10b;
        src113 <= 16'hcef;
        src114 <= 16'hc7c4;
        src115 <= 16'h6855;
        src116 <= 16'h7e6d;
        src117 <= 16'h7675;
        src118 <= 16'h85cb;
        src119 <= 16'hdb64;
        src120 <= 16'h51d6;
        src121 <= 16'hc8dd;
        src122 <= 16'he510;
        src123 <= 16'h9259;
        src124 <= 16'hf5e3;
        src125 <= 16'hb353;
        src126 <= 16'h4e55;
        src127 <= 16'h9d5;
        src128 <= 16'hfb43;
        src129 <= 16'hcc93;
        src130 <= 16'hb60f;
        src131 <= 16'h264;
        src132 <= 16'h5bb;
        src133 <= 16'hb768;
        src134 <= 16'h63d0;
        src135 <= 16'h21c6;
        src136 <= 16'he473;
        src137 <= 16'h4f53;
        src138 <= 16'h84d9;
        src139 <= 16'hd4f4;
        src140 <= 16'h55ef;
        src141 <= 16'hc223;
        src142 <= 16'h2842;
        src143 <= 16'h5889;
        src144 <= 16'h5023;
        src145 <= 16'hcd2c;
        src146 <= 16'hfd19;
        src147 <= 16'h476;
        src148 <= 16'h15ab;
        src149 <= 16'hf8e6;
        src150 <= 16'h7bd2;
        src151 <= 16'h9ee;
        src152 <= 16'h883d;
        src153 <= 16'hd2d1;
        src154 <= 16'h8adb;
        src155 <= 16'h32ce;
        src156 <= 16'he743;
        src157 <= 16'h9424;
        src158 <= 16'hf9d4;
        src159 <= 16'h6683;
        src160 <= 16'h6d3e;
        src161 <= 16'h14f3;
        src162 <= 16'h8fa6;
        src163 <= 16'h9815;
        src164 <= 16'h5418;
        src165 <= 16'h23d0;
        src166 <= 16'h925b;
        src167 <= 16'h363;
        src168 <= 16'hcbca;
        src169 <= 16'h9156;
        src170 <= 16'h6635;
        src171 <= 16'h9a9;
        src172 <= 16'hdce7;
        src173 <= 16'h9397;
        src174 <= 16'hde5e;
        src175 <= 16'h8834;
        src176 <= 16'h8806;
        src177 <= 16'hfebb;
        src178 <= 16'h5942;
        src179 <= 16'h4953;
        src180 <= 16'hbb06;
        src181 <= 16'h7ff8;
        src182 <= 16'hae3f;
        src183 <= 16'h591a;
        src184 <= 16'h5902;
        exp <= 24'h5be037;
        #1
        src0 <= 16'h27ad;
        src1 <= 16'h566c;
        src2 <= 16'hb592;
        src3 <= 16'hdb2;
        src4 <= 16'h8ff7;
        src5 <= 16'h5482;
        src6 <= 16'hc10a;
        src7 <= 16'h486;
        src8 <= 16'h9e77;
        src9 <= 16'hdc11;
        src10 <= 16'h23ac;
        src11 <= 16'hc6fa;
        src12 <= 16'h772b;
        src13 <= 16'hf928;
        src14 <= 16'h6cc8;
        src15 <= 16'h619c;
        src16 <= 16'h36e3;
        src17 <= 16'h37d2;
        src18 <= 16'h836b;
        src19 <= 16'h9f52;
        src20 <= 16'h6ae7;
        src21 <= 16'haf2d;
        src22 <= 16'h7237;
        src23 <= 16'h3bd3;
        src24 <= 16'hbbf9;
        src25 <= 16'hb83;
        src26 <= 16'h4098;
        src27 <= 16'h3bd4;
        src28 <= 16'hc8a8;
        src29 <= 16'h8182;
        src30 <= 16'h3a22;
        src31 <= 16'hab35;
        src32 <= 16'h16d7;
        src33 <= 16'he219;
        src34 <= 16'hdd39;
        src35 <= 16'h43b5;
        src36 <= 16'h3276;
        src37 <= 16'he452;
        src38 <= 16'h8cdb;
        src39 <= 16'hd289;
        src40 <= 16'he8bb;
        src41 <= 16'h46a7;
        src42 <= 16'h17b9;
        src43 <= 16'ha7a0;
        src44 <= 16'h1892;
        src45 <= 16'h8d99;
        src46 <= 16'h205b;
        src47 <= 16'hd408;
        src48 <= 16'hbdbd;
        src49 <= 16'h6ee;
        src50 <= 16'h12cb;
        src51 <= 16'h84b1;
        src52 <= 16'hbb63;
        src53 <= 16'h6d51;
        src54 <= 16'h3f90;
        src55 <= 16'hadf;
        src56 <= 16'hdaa5;
        src57 <= 16'h76d7;
        src58 <= 16'he3b7;
        src59 <= 16'hda6d;
        src60 <= 16'hf4bd;
        src61 <= 16'h4c86;
        src62 <= 16'h1286;
        src63 <= 16'h72fc;
        src64 <= 16'hba9c;
        src65 <= 16'h6bac;
        src66 <= 16'h2a87;
        src67 <= 16'h9843;
        src68 <= 16'h52d3;
        src69 <= 16'hcefb;
        src70 <= 16'h13f7;
        src71 <= 16'hb7ba;
        src72 <= 16'h50b7;
        src73 <= 16'haa3;
        src74 <= 16'h90a1;
        src75 <= 16'ha1e5;
        src76 <= 16'he581;
        src77 <= 16'h3f4c;
        src78 <= 16'hd855;
        src79 <= 16'hca91;
        src80 <= 16'h30f9;
        src81 <= 16'h119f;
        src82 <= 16'hccd2;
        src83 <= 16'h37cc;
        src84 <= 16'h2076;
        src85 <= 16'h723f;
        src86 <= 16'hd2ee;
        src87 <= 16'h17e9;
        src88 <= 16'h48b8;
        src89 <= 16'h85c6;
        src90 <= 16'h53cc;
        src91 <= 16'h5b00;
        src92 <= 16'h78ba;
        src93 <= 16'hb1fd;
        src94 <= 16'hf43f;
        src95 <= 16'he106;
        src96 <= 16'hd28c;
        src97 <= 16'hc5a1;
        src98 <= 16'he658;
        src99 <= 16'h91b3;
        src100 <= 16'h1767;
        src101 <= 16'h7065;
        src102 <= 16'h3de;
        src103 <= 16'he2e0;
        src104 <= 16'hb809;
        src105 <= 16'hfd1d;
        src106 <= 16'hf14f;
        src107 <= 16'h504d;
        src108 <= 16'h5211;
        src109 <= 16'hc4a9;
        src110 <= 16'hcbba;
        src111 <= 16'h9238;
        src112 <= 16'h9bd1;
        src113 <= 16'h5165;
        src114 <= 16'hbda5;
        src115 <= 16'h37a3;
        src116 <= 16'h5886;
        src117 <= 16'h6e1f;
        src118 <= 16'h5d60;
        src119 <= 16'hea42;
        src120 <= 16'hc940;
        src121 <= 16'hee86;
        src122 <= 16'he364;
        src123 <= 16'h1110;
        src124 <= 16'h6d4d;
        src125 <= 16'h7017;
        src126 <= 16'hd9f3;
        src127 <= 16'hbed8;
        src128 <= 16'hf2f8;
        src129 <= 16'h745c;
        src130 <= 16'he1f8;
        src131 <= 16'hab1b;
        src132 <= 16'h7881;
        src133 <= 16'h36de;
        src134 <= 16'h82cb;
        src135 <= 16'h48c4;
        src136 <= 16'h4cf3;
        src137 <= 16'hdca3;
        src138 <= 16'hc364;
        src139 <= 16'h151f;
        src140 <= 16'h232;
        src141 <= 16'h5c96;
        src142 <= 16'h268c;
        src143 <= 16'h13aa;
        src144 <= 16'h2fe0;
        src145 <= 16'hf231;
        src146 <= 16'hd0d4;
        src147 <= 16'h6bcd;
        src148 <= 16'hd4fa;
        src149 <= 16'ha18a;
        src150 <= 16'h55b4;
        src151 <= 16'hc9bc;
        src152 <= 16'h6fe4;
        src153 <= 16'h1716;
        src154 <= 16'h4272;
        src155 <= 16'hab01;
        src156 <= 16'h2719;
        src157 <= 16'heb7c;
        src158 <= 16'h6f6e;
        src159 <= 16'h87fa;
        src160 <= 16'hc605;
        src161 <= 16'h65bc;
        src162 <= 16'h9d7a;
        src163 <= 16'h5506;
        src164 <= 16'hb342;
        src165 <= 16'h7b02;
        src166 <= 16'h259f;
        src167 <= 16'hdd6f;
        src168 <= 16'hd8db;
        src169 <= 16'h2a;
        src170 <= 16'ha05c;
        src171 <= 16'h5ed;
        src172 <= 16'ha98a;
        src173 <= 16'hed0d;
        src174 <= 16'hc82;
        src175 <= 16'hbdec;
        src176 <= 16'h53e0;
        src177 <= 16'hd3c7;
        src178 <= 16'ha519;
        src179 <= 16'h6352;
        src180 <= 16'h3dc0;
        src181 <= 16'hb3c1;
        src182 <= 16'h96b0;
        src183 <= 16'hec5c;
        src184 <= 16'h2edc;
        exp <= 24'h5d07ad;
        #1
        src0 <= 16'h1f7a;
        src1 <= 16'h1ba4;
        src2 <= 16'h48b7;
        src3 <= 16'h2ce7;
        src4 <= 16'h11f0;
        src5 <= 16'h2eb;
        src6 <= 16'hdcae;
        src7 <= 16'h4116;
        src8 <= 16'h530e;
        src9 <= 16'h3454;
        src10 <= 16'h1d9f;
        src11 <= 16'h5eaa;
        src12 <= 16'hd39a;
        src13 <= 16'ha2a4;
        src14 <= 16'haba9;
        src15 <= 16'hd331;
        src16 <= 16'h1015;
        src17 <= 16'hfca1;
        src18 <= 16'h9bcc;
        src19 <= 16'h8b08;
        src20 <= 16'hfc0f;
        src21 <= 16'he7ed;
        src22 <= 16'h3947;
        src23 <= 16'h4936;
        src24 <= 16'h384;
        src25 <= 16'h7aab;
        src26 <= 16'h599c;
        src27 <= 16'hd789;
        src28 <= 16'h38fb;
        src29 <= 16'hc28;
        src30 <= 16'h153;
        src31 <= 16'hd046;
        src32 <= 16'h35b2;
        src33 <= 16'h23b9;
        src34 <= 16'h9b64;
        src35 <= 16'hfee6;
        src36 <= 16'h1f0b;
        src37 <= 16'h6549;
        src38 <= 16'ha6f1;
        src39 <= 16'h22fa;
        src40 <= 16'h4ae5;
        src41 <= 16'h5999;
        src42 <= 16'hd4df;
        src43 <= 16'he09a;
        src44 <= 16'h6163;
        src45 <= 16'h76c5;
        src46 <= 16'h986e;
        src47 <= 16'h20bb;
        src48 <= 16'h7e38;
        src49 <= 16'hdbf5;
        src50 <= 16'h560d;
        src51 <= 16'h2dd5;
        src52 <= 16'ha0d8;
        src53 <= 16'h83e2;
        src54 <= 16'h3c0;
        src55 <= 16'h7b14;
        src56 <= 16'h771d;
        src57 <= 16'he971;
        src58 <= 16'hcb4f;
        src59 <= 16'h9e9;
        src60 <= 16'hf821;
        src61 <= 16'hd48e;
        src62 <= 16'hcef1;
        src63 <= 16'h2bf7;
        src64 <= 16'h2ed0;
        src65 <= 16'h8451;
        src66 <= 16'h8a44;
        src67 <= 16'h2273;
        src68 <= 16'h4e47;
        src69 <= 16'h1c17;
        src70 <= 16'h1280;
        src71 <= 16'h7f94;
        src72 <= 16'h9e41;
        src73 <= 16'h3bbe;
        src74 <= 16'h3603;
        src75 <= 16'hda8d;
        src76 <= 16'hab37;
        src77 <= 16'h5aa3;
        src78 <= 16'hbc5;
        src79 <= 16'ha055;
        src80 <= 16'h4c56;
        src81 <= 16'h95a7;
        src82 <= 16'h2027;
        src83 <= 16'hd7ba;
        src84 <= 16'h9367;
        src85 <= 16'h7f95;
        src86 <= 16'hc3b8;
        src87 <= 16'h3c0d;
        src88 <= 16'hf874;
        src89 <= 16'hf3f6;
        src90 <= 16'ha2d5;
        src91 <= 16'h2f7;
        src92 <= 16'h1a2;
        src93 <= 16'h2ea1;
        src94 <= 16'hb587;
        src95 <= 16'h26e7;
        src96 <= 16'h1c9c;
        src97 <= 16'h76fe;
        src98 <= 16'h9382;
        src99 <= 16'he80c;
        src100 <= 16'hf0d5;
        src101 <= 16'hb671;
        src102 <= 16'h8622;
        src103 <= 16'h2e6e;
        src104 <= 16'h7de6;
        src105 <= 16'h934d;
        src106 <= 16'h9e3d;
        src107 <= 16'h6e5;
        src108 <= 16'h9314;
        src109 <= 16'h5722;
        src110 <= 16'ha851;
        src111 <= 16'h6bd2;
        src112 <= 16'h9bb9;
        src113 <= 16'h7b93;
        src114 <= 16'h3ed0;
        src115 <= 16'hda85;
        src116 <= 16'hdfae;
        src117 <= 16'h8ed9;
        src118 <= 16'h5e75;
        src119 <= 16'h7a96;
        src120 <= 16'hfcd7;
        src121 <= 16'h179a;
        src122 <= 16'h1af8;
        src123 <= 16'hf83a;
        src124 <= 16'h53b4;
        src125 <= 16'hb156;
        src126 <= 16'h4b5a;
        src127 <= 16'heee7;
        src128 <= 16'hf4d4;
        src129 <= 16'he2d2;
        src130 <= 16'h8648;
        src131 <= 16'h7921;
        src132 <= 16'h56ee;
        src133 <= 16'h5b7e;
        src134 <= 16'h698f;
        src135 <= 16'h46aa;
        src136 <= 16'h2909;
        src137 <= 16'h1c50;
        src138 <= 16'hfc6f;
        src139 <= 16'hb30a;
        src140 <= 16'h823a;
        src141 <= 16'h816c;
        src142 <= 16'h24ca;
        src143 <= 16'h4c13;
        src144 <= 16'h3d34;
        src145 <= 16'h6c5;
        src146 <= 16'h3e0;
        src147 <= 16'h8571;
        src148 <= 16'h6e61;
        src149 <= 16'hdbf2;
        src150 <= 16'hde17;
        src151 <= 16'h5dc;
        src152 <= 16'h9530;
        src153 <= 16'ha564;
        src154 <= 16'hb6ee;
        src155 <= 16'h59a7;
        src156 <= 16'h1d03;
        src157 <= 16'h7901;
        src158 <= 16'hac1f;
        src159 <= 16'h6a0d;
        src160 <= 16'h8fa;
        src161 <= 16'h8ae8;
        src162 <= 16'h359d;
        src163 <= 16'h59a8;
        src164 <= 16'h93db;
        src165 <= 16'h28ef;
        src166 <= 16'h3dee;
        src167 <= 16'h9e2c;
        src168 <= 16'h11e8;
        src169 <= 16'hd6a2;
        src170 <= 16'hde76;
        src171 <= 16'h47cf;
        src172 <= 16'h35ff;
        src173 <= 16'h5d2a;
        src174 <= 16'hc095;
        src175 <= 16'h6059;
        src176 <= 16'h3b6b;
        src177 <= 16'he57c;
        src178 <= 16'h21b;
        src179 <= 16'h3894;
        src180 <= 16'he042;
        src181 <= 16'h7a9a;
        src182 <= 16'h44fe;
        src183 <= 16'h8a89;
        src184 <= 16'h7948;
        exp <= 24'h547fab;
        #1
        src0 <= 16'ha227;
        src1 <= 16'h3687;
        src2 <= 16'hee93;
        src3 <= 16'hec1d;
        src4 <= 16'hb2c4;
        src5 <= 16'h1852;
        src6 <= 16'hcd39;
        src7 <= 16'hac1f;
        src8 <= 16'h2918;
        src9 <= 16'hdca4;
        src10 <= 16'ha9d2;
        src11 <= 16'h228c;
        src12 <= 16'h19a1;
        src13 <= 16'hf182;
        src14 <= 16'h77cd;
        src15 <= 16'h2b4b;
        src16 <= 16'hdafa;
        src17 <= 16'h4997;
        src18 <= 16'h636;
        src19 <= 16'hf11c;
        src20 <= 16'h3bb;
        src21 <= 16'hf684;
        src22 <= 16'h40b5;
        src23 <= 16'hbc7c;
        src24 <= 16'hb782;
        src25 <= 16'hfd83;
        src26 <= 16'h431b;
        src27 <= 16'h4662;
        src28 <= 16'h243b;
        src29 <= 16'hd4ac;
        src30 <= 16'h1737;
        src31 <= 16'h4c18;
        src32 <= 16'h1d47;
        src33 <= 16'h17d7;
        src34 <= 16'h7092;
        src35 <= 16'hca6f;
        src36 <= 16'h4ef;
        src37 <= 16'h735b;
        src38 <= 16'ha8f6;
        src39 <= 16'h5a1f;
        src40 <= 16'he80d;
        src41 <= 16'h4b2f;
        src42 <= 16'hcdfd;
        src43 <= 16'h40d8;
        src44 <= 16'h8b76;
        src45 <= 16'hfd98;
        src46 <= 16'h902c;
        src47 <= 16'h2987;
        src48 <= 16'h99af;
        src49 <= 16'h78a3;
        src50 <= 16'hffa6;
        src51 <= 16'h7f35;
        src52 <= 16'h6a8;
        src53 <= 16'h3bed;
        src54 <= 16'h6a72;
        src55 <= 16'h1efd;
        src56 <= 16'h8dfe;
        src57 <= 16'ha685;
        src58 <= 16'h5670;
        src59 <= 16'ha5bf;
        src60 <= 16'hbd2;
        src61 <= 16'ha493;
        src62 <= 16'hf31c;
        src63 <= 16'he089;
        src64 <= 16'h77e6;
        src65 <= 16'h23c2;
        src66 <= 16'h5e23;
        src67 <= 16'h24e7;
        src68 <= 16'hf056;
        src69 <= 16'h7f7b;
        src70 <= 16'he622;
        src71 <= 16'hc5c2;
        src72 <= 16'h34bd;
        src73 <= 16'hdf1c;
        src74 <= 16'hd267;
        src75 <= 16'hfd5b;
        src76 <= 16'h1f03;
        src77 <= 16'h6f87;
        src78 <= 16'h14da;
        src79 <= 16'hf8c8;
        src80 <= 16'ha0e0;
        src81 <= 16'hd6c6;
        src82 <= 16'h782b;
        src83 <= 16'hf36;
        src84 <= 16'hba66;
        src85 <= 16'hfef5;
        src86 <= 16'h23ac;
        src87 <= 16'h998e;
        src88 <= 16'hd43c;
        src89 <= 16'h5d27;
        src90 <= 16'hca27;
        src91 <= 16'h18ea;
        src92 <= 16'h4f79;
        src93 <= 16'h83e;
        src94 <= 16'h3633;
        src95 <= 16'h8194;
        src96 <= 16'hd7c6;
        src97 <= 16'hb783;
        src98 <= 16'he06a;
        src99 <= 16'hb4a4;
        src100 <= 16'h7fd3;
        src101 <= 16'hbfa7;
        src102 <= 16'h32b7;
        src103 <= 16'h262b;
        src104 <= 16'he667;
        src105 <= 16'h987f;
        src106 <= 16'hd40c;
        src107 <= 16'hc308;
        src108 <= 16'h981b;
        src109 <= 16'h3ce4;
        src110 <= 16'hdcb1;
        src111 <= 16'h2ba9;
        src112 <= 16'h11f8;
        src113 <= 16'h782;
        src114 <= 16'h714a;
        src115 <= 16'h47c7;
        src116 <= 16'h491b;
        src117 <= 16'h6aa;
        src118 <= 16'h8b1e;
        src119 <= 16'h4b3e;
        src120 <= 16'h8c71;
        src121 <= 16'heb15;
        src122 <= 16'h69c0;
        src123 <= 16'hc428;
        src124 <= 16'h4a11;
        src125 <= 16'hd099;
        src126 <= 16'hb6bf;
        src127 <= 16'h791e;
        src128 <= 16'hd26f;
        src129 <= 16'hc0db;
        src130 <= 16'ha063;
        src131 <= 16'h1146;
        src132 <= 16'h3b15;
        src133 <= 16'haac8;
        src134 <= 16'h11f0;
        src135 <= 16'hf278;
        src136 <= 16'h82b9;
        src137 <= 16'h16ed;
        src138 <= 16'hf995;
        src139 <= 16'h6236;
        src140 <= 16'hdbf2;
        src141 <= 16'h804f;
        src142 <= 16'h78ab;
        src143 <= 16'ha71f;
        src144 <= 16'hc555;
        src145 <= 16'he0bd;
        src146 <= 16'h837c;
        src147 <= 16'h2894;
        src148 <= 16'h197b;
        src149 <= 16'h6152;
        src150 <= 16'h3305;
        src151 <= 16'h9dc9;
        src152 <= 16'h78eb;
        src153 <= 16'hff72;
        src154 <= 16'h9e52;
        src155 <= 16'h7d79;
        src156 <= 16'h9727;
        src157 <= 16'h226d;
        src158 <= 16'h6c9b;
        src159 <= 16'hb971;
        src160 <= 16'h68bc;
        src161 <= 16'h328e;
        src162 <= 16'hb6ca;
        src163 <= 16'hef11;
        src164 <= 16'hbef0;
        src165 <= 16'h3617;
        src166 <= 16'he363;
        src167 <= 16'hd30d;
        src168 <= 16'hbf92;
        src169 <= 16'h40ab;
        src170 <= 16'hf8a7;
        src171 <= 16'h1665;
        src172 <= 16'hd73f;
        src173 <= 16'h82f1;
        src174 <= 16'h774c;
        src175 <= 16'h25b6;
        src176 <= 16'ha06b;
        src177 <= 16'h2763;
        src178 <= 16'hf8b0;
        src179 <= 16'hc021;
        src180 <= 16'hefc9;
        src181 <= 16'h449c;
        src182 <= 16'h2799;
        src183 <= 16'hb509;
        src184 <= 16'hc874;
        exp <= 24'h5f9436;
        #1
        src0 <= 16'h5f88;
        src1 <= 16'h72e1;
        src2 <= 16'hf9c7;
        src3 <= 16'h65fa;
        src4 <= 16'h765f;
        src5 <= 16'h730c;
        src6 <= 16'h3c1f;
        src7 <= 16'h8e52;
        src8 <= 16'hae1d;
        src9 <= 16'h76a4;
        src10 <= 16'ha36c;
        src11 <= 16'hfeb8;
        src12 <= 16'hc35e;
        src13 <= 16'h6dd7;
        src14 <= 16'h7f88;
        src15 <= 16'hf5c0;
        src16 <= 16'hc1f8;
        src17 <= 16'h5624;
        src18 <= 16'h474b;
        src19 <= 16'hd1a6;
        src20 <= 16'h7406;
        src21 <= 16'h4dc3;
        src22 <= 16'h6aa6;
        src23 <= 16'h953d;
        src24 <= 16'he58a;
        src25 <= 16'h9562;
        src26 <= 16'h157b;
        src27 <= 16'h2d4b;
        src28 <= 16'h4746;
        src29 <= 16'h8c05;
        src30 <= 16'hefd3;
        src31 <= 16'h40de;
        src32 <= 16'hd465;
        src33 <= 16'h7025;
        src34 <= 16'hc028;
        src35 <= 16'h3893;
        src36 <= 16'h100e;
        src37 <= 16'hea3a;
        src38 <= 16'hec07;
        src39 <= 16'h7671;
        src40 <= 16'h798a;
        src41 <= 16'hf48d;
        src42 <= 16'h9132;
        src43 <= 16'hdaef;
        src44 <= 16'h6fd5;
        src45 <= 16'h7b3e;
        src46 <= 16'hc318;
        src47 <= 16'h657e;
        src48 <= 16'h383f;
        src49 <= 16'h24e5;
        src50 <= 16'h1ea0;
        src51 <= 16'hb2fe;
        src52 <= 16'h73b;
        src53 <= 16'h29b1;
        src54 <= 16'hb4e7;
        src55 <= 16'h6106;
        src56 <= 16'h2406;
        src57 <= 16'hc589;
        src58 <= 16'h6100;
        src59 <= 16'h9c56;
        src60 <= 16'hbb10;
        src61 <= 16'hb98d;
        src62 <= 16'hb32e;
        src63 <= 16'h206a;
        src64 <= 16'h4289;
        src65 <= 16'hb620;
        src66 <= 16'h447;
        src67 <= 16'h6f59;
        src68 <= 16'h62bf;
        src69 <= 16'ha3ec;
        src70 <= 16'h73cc;
        src71 <= 16'heb75;
        src72 <= 16'h187d;
        src73 <= 16'haf00;
        src74 <= 16'he74a;
        src75 <= 16'h8db5;
        src76 <= 16'h7ded;
        src77 <= 16'h506c;
        src78 <= 16'hf225;
        src79 <= 16'h9189;
        src80 <= 16'h3bd4;
        src81 <= 16'hcd03;
        src82 <= 16'h3226;
        src83 <= 16'h4194;
        src84 <= 16'hc324;
        src85 <= 16'hb761;
        src86 <= 16'h5b98;
        src87 <= 16'h7d8;
        src88 <= 16'h8004;
        src89 <= 16'hf2dd;
        src90 <= 16'h8a0;
        src91 <= 16'h8ddd;
        src92 <= 16'hc522;
        src93 <= 16'h969f;
        src94 <= 16'hd69b;
        src95 <= 16'h8d5b;
        src96 <= 16'haf5c;
        src97 <= 16'hab;
        src98 <= 16'h1360;
        src99 <= 16'hb0ec;
        src100 <= 16'h2c71;
        src101 <= 16'hd0ed;
        src102 <= 16'h78a;
        src103 <= 16'hf1c1;
        src104 <= 16'ha1f3;
        src105 <= 16'ha0c2;
        src106 <= 16'hcb83;
        src107 <= 16'h225d;
        src108 <= 16'h8abd;
        src109 <= 16'hf831;
        src110 <= 16'ha057;
        src111 <= 16'hcc59;
        src112 <= 16'hbcf0;
        src113 <= 16'h43d1;
        src114 <= 16'h3583;
        src115 <= 16'ha47;
        src116 <= 16'h9f27;
        src117 <= 16'ha39c;
        src118 <= 16'h283c;
        src119 <= 16'hdaa2;
        src120 <= 16'h5305;
        src121 <= 16'h90d1;
        src122 <= 16'h7646;
        src123 <= 16'hab1d;
        src124 <= 16'h9514;
        src125 <= 16'h6837;
        src126 <= 16'h814;
        src127 <= 16'h6c6a;
        src128 <= 16'h9d02;
        src129 <= 16'h9a09;
        src130 <= 16'hc590;
        src131 <= 16'h6931;
        src132 <= 16'hee21;
        src133 <= 16'h71f0;
        src134 <= 16'hfbac;
        src135 <= 16'h411a;
        src136 <= 16'h93f9;
        src137 <= 16'hecc9;
        src138 <= 16'h2ea1;
        src139 <= 16'ha8af;
        src140 <= 16'he2f5;
        src141 <= 16'h5b0a;
        src142 <= 16'hc831;
        src143 <= 16'h1dd6;
        src144 <= 16'h2542;
        src145 <= 16'hbb7e;
        src146 <= 16'heb9f;
        src147 <= 16'hc5e9;
        src148 <= 16'hf6f4;
        src149 <= 16'h29a8;
        src150 <= 16'h257b;
        src151 <= 16'h349;
        src152 <= 16'hd205;
        src153 <= 16'h7cc0;
        src154 <= 16'hc8c0;
        src155 <= 16'hb5a0;
        src156 <= 16'hace3;
        src157 <= 16'h47bc;
        src158 <= 16'h8436;
        src159 <= 16'h2403;
        src160 <= 16'h5045;
        src161 <= 16'ha3e6;
        src162 <= 16'hfc5f;
        src163 <= 16'h3e5a;
        src164 <= 16'h80f6;
        src165 <= 16'h3692;
        src166 <= 16'ha669;
        src167 <= 16'h9c31;
        src168 <= 16'h258b;
        src169 <= 16'hb73a;
        src170 <= 16'h715;
        src171 <= 16'hc7df;
        src172 <= 16'h8fb6;
        src173 <= 16'h2ee4;
        src174 <= 16'h3639;
        src175 <= 16'h52cc;
        src176 <= 16'h686c;
        src177 <= 16'h9311;
        src178 <= 16'h9452;
        src179 <= 16'h74c2;
        src180 <= 16'h9e1c;
        src181 <= 16'h7f34;
        src182 <= 16'hafc7;
        src183 <= 16'h25e9;
        src184 <= 16'h3855;
        exp <= 24'h5e51be;
        #1
        src0 <= 16'hface;
        src1 <= 16'hf9cf;
        src2 <= 16'hb2d6;
        src3 <= 16'h1280;
        src4 <= 16'hfa94;
        src5 <= 16'h3a95;
        src6 <= 16'h5607;
        src7 <= 16'h6101;
        src8 <= 16'h6cd0;
        src9 <= 16'hf852;
        src10 <= 16'h1b14;
        src11 <= 16'h670;
        src12 <= 16'he8e6;
        src13 <= 16'h5ee0;
        src14 <= 16'he36a;
        src15 <= 16'h1a68;
        src16 <= 16'h375b;
        src17 <= 16'h306d;
        src18 <= 16'h64af;
        src19 <= 16'h1090;
        src20 <= 16'h94aa;
        src21 <= 16'h6320;
        src22 <= 16'h1c4f;
        src23 <= 16'h271;
        src24 <= 16'h8309;
        src25 <= 16'hfc30;
        src26 <= 16'had1c;
        src27 <= 16'h1801;
        src28 <= 16'h9010;
        src29 <= 16'h12c8;
        src30 <= 16'hfb9c;
        src31 <= 16'ha9a4;
        src32 <= 16'haff;
        src33 <= 16'hbac5;
        src34 <= 16'h792b;
        src35 <= 16'hf873;
        src36 <= 16'h562f;
        src37 <= 16'h54d3;
        src38 <= 16'hc71d;
        src39 <= 16'h1509;
        src40 <= 16'h1b8f;
        src41 <= 16'h2522;
        src42 <= 16'hffec;
        src43 <= 16'hb64b;
        src44 <= 16'h10dd;
        src45 <= 16'he72e;
        src46 <= 16'h144b;
        src47 <= 16'h730c;
        src48 <= 16'hd20;
        src49 <= 16'h3b71;
        src50 <= 16'h57be;
        src51 <= 16'he262;
        src52 <= 16'h97ec;
        src53 <= 16'hba63;
        src54 <= 16'hc7b0;
        src55 <= 16'h3f6f;
        src56 <= 16'h99f7;
        src57 <= 16'h1f6e;
        src58 <= 16'h1368;
        src59 <= 16'h700f;
        src60 <= 16'h247e;
        src61 <= 16'h84da;
        src62 <= 16'h2a8e;
        src63 <= 16'hb214;
        src64 <= 16'h88ca;
        src65 <= 16'hde39;
        src66 <= 16'hb98f;
        src67 <= 16'h9bf0;
        src68 <= 16'h35ff;
        src69 <= 16'h5e10;
        src70 <= 16'h901a;
        src71 <= 16'h1cac;
        src72 <= 16'ha591;
        src73 <= 16'he170;
        src74 <= 16'hb445;
        src75 <= 16'h1aec;
        src76 <= 16'ha966;
        src77 <= 16'h62c0;
        src78 <= 16'h36fd;
        src79 <= 16'hb940;
        src80 <= 16'h496c;
        src81 <= 16'heec6;
        src82 <= 16'h3f72;
        src83 <= 16'h666a;
        src84 <= 16'h6fbb;
        src85 <= 16'ha064;
        src86 <= 16'h88d5;
        src87 <= 16'h98f6;
        src88 <= 16'hc5b;
        src89 <= 16'hb0d0;
        src90 <= 16'h9f3a;
        src91 <= 16'he822;
        src92 <= 16'he669;
        src93 <= 16'h5cba;
        src94 <= 16'h4215;
        src95 <= 16'h5ac6;
        src96 <= 16'hb42f;
        src97 <= 16'hff81;
        src98 <= 16'heb7a;
        src99 <= 16'he5;
        src100 <= 16'h2712;
        src101 <= 16'hc2fa;
        src102 <= 16'ha3;
        src103 <= 16'he2d7;
        src104 <= 16'h768c;
        src105 <= 16'h6574;
        src106 <= 16'he1c2;
        src107 <= 16'hc9a5;
        src108 <= 16'h34e9;
        src109 <= 16'hb831;
        src110 <= 16'he2f0;
        src111 <= 16'hcc40;
        src112 <= 16'h4d73;
        src113 <= 16'h46b7;
        src114 <= 16'hb358;
        src115 <= 16'hd736;
        src116 <= 16'haf38;
        src117 <= 16'h23c2;
        src118 <= 16'h8b20;
        src119 <= 16'hc708;
        src120 <= 16'ha17;
        src121 <= 16'h7f0d;
        src122 <= 16'hf792;
        src123 <= 16'h29af;
        src124 <= 16'hd528;
        src125 <= 16'h683f;
        src126 <= 16'h231a;
        src127 <= 16'h94ed;
        src128 <= 16'hf838;
        src129 <= 16'hee79;
        src130 <= 16'hcb50;
        src131 <= 16'h2f0c;
        src132 <= 16'hc54d;
        src133 <= 16'hbe74;
        src134 <= 16'h4cc3;
        src135 <= 16'h7fec;
        src136 <= 16'h1422;
        src137 <= 16'h5ffb;
        src138 <= 16'h4f12;
        src139 <= 16'hdbb7;
        src140 <= 16'h8ee9;
        src141 <= 16'h15f8;
        src142 <= 16'h2899;
        src143 <= 16'h85d6;
        src144 <= 16'hf910;
        src145 <= 16'he252;
        src146 <= 16'h166b;
        src147 <= 16'hf1f4;
        src148 <= 16'h3166;
        src149 <= 16'hc0ed;
        src150 <= 16'h84e5;
        src151 <= 16'h539;
        src152 <= 16'h9743;
        src153 <= 16'he261;
        src154 <= 16'h24e7;
        src155 <= 16'h78e;
        src156 <= 16'h5d32;
        src157 <= 16'hb5a2;
        src158 <= 16'h6399;
        src159 <= 16'hbf16;
        src160 <= 16'h9cb3;
        src161 <= 16'hefcb;
        src162 <= 16'h6ae1;
        src163 <= 16'hf69c;
        src164 <= 16'h9cae;
        src165 <= 16'h483d;
        src166 <= 16'h393f;
        src167 <= 16'h20e9;
        src168 <= 16'hf796;
        src169 <= 16'hd740;
        src170 <= 16'h28b0;
        src171 <= 16'h87a2;
        src172 <= 16'h70f9;
        src173 <= 16'h88a5;
        src174 <= 16'h9a44;
        src175 <= 16'hea5a;
        src176 <= 16'hce9f;
        src177 <= 16'hbf01;
        src178 <= 16'he082;
        src179 <= 16'he82c;
        src180 <= 16'h4498;
        src181 <= 16'h462b;
        src182 <= 16'haaad;
        src183 <= 16'hce42;
        src184 <= 16'hb39f;
        exp <= 24'h5e5718;
        #1
        src0 <= 16'h7c8e;
        src1 <= 16'h2827;
        src2 <= 16'he118;
        src3 <= 16'h49c5;
        src4 <= 16'h5d3c;
        src5 <= 16'hb32c;
        src6 <= 16'h8e84;
        src7 <= 16'h1ef;
        src8 <= 16'h96f0;
        src9 <= 16'h88a9;
        src10 <= 16'h60e4;
        src11 <= 16'h5e51;
        src12 <= 16'hfbbb;
        src13 <= 16'h593a;
        src14 <= 16'hc13c;
        src15 <= 16'h81d3;
        src16 <= 16'hbbec;
        src17 <= 16'h5e1;
        src18 <= 16'h9939;
        src19 <= 16'ha297;
        src20 <= 16'he08f;
        src21 <= 16'h4624;
        src22 <= 16'h1744;
        src23 <= 16'h66af;
        src24 <= 16'hb990;
        src25 <= 16'h227b;
        src26 <= 16'h7ef;
        src27 <= 16'hff14;
        src28 <= 16'h910b;
        src29 <= 16'ha956;
        src30 <= 16'h4164;
        src31 <= 16'h2587;
        src32 <= 16'h1f1f;
        src33 <= 16'h272a;
        src34 <= 16'h48fc;
        src35 <= 16'h55b4;
        src36 <= 16'hfa7f;
        src37 <= 16'h2f91;
        src38 <= 16'h6bb0;
        src39 <= 16'h8de5;
        src40 <= 16'h52d4;
        src41 <= 16'h17e6;
        src42 <= 16'he8f7;
        src43 <= 16'h1569;
        src44 <= 16'hd8a5;
        src45 <= 16'h2905;
        src46 <= 16'he26c;
        src47 <= 16'h9a1e;
        src48 <= 16'h6c5f;
        src49 <= 16'h505;
        src50 <= 16'h476b;
        src51 <= 16'h8729;
        src52 <= 16'h1cdf;
        src53 <= 16'h895e;
        src54 <= 16'h7b6;
        src55 <= 16'h1a62;
        src56 <= 16'hfcf2;
        src57 <= 16'h2fac;
        src58 <= 16'h1cd8;
        src59 <= 16'h69f5;
        src60 <= 16'h2f1;
        src61 <= 16'haa97;
        src62 <= 16'had53;
        src63 <= 16'h6c3f;
        src64 <= 16'hcf8f;
        src65 <= 16'hf171;
        src66 <= 16'h9c1c;
        src67 <= 16'hb9d9;
        src68 <= 16'h6bad;
        src69 <= 16'hbb75;
        src70 <= 16'h34a8;
        src71 <= 16'h89fd;
        src72 <= 16'h5a23;
        src73 <= 16'h23f;
        src74 <= 16'hb72f;
        src75 <= 16'h497c;
        src76 <= 16'h55a3;
        src77 <= 16'h31e5;
        src78 <= 16'h12d7;
        src79 <= 16'hb3d6;
        src80 <= 16'heb63;
        src81 <= 16'h7659;
        src82 <= 16'hed35;
        src83 <= 16'h347c;
        src84 <= 16'h3192;
        src85 <= 16'hfd5c;
        src86 <= 16'hf159;
        src87 <= 16'h9f56;
        src88 <= 16'h1076;
        src89 <= 16'h64ea;
        src90 <= 16'h17c9;
        src91 <= 16'h3aa1;
        src92 <= 16'h43fe;
        src93 <= 16'hb5cd;
        src94 <= 16'h741c;
        src95 <= 16'h14da;
        src96 <= 16'h90bb;
        src97 <= 16'hda3;
        src98 <= 16'h7034;
        src99 <= 16'h5169;
        src100 <= 16'hc5ea;
        src101 <= 16'hd30c;
        src102 <= 16'hd4d2;
        src103 <= 16'h55b1;
        src104 <= 16'he52a;
        src105 <= 16'h4947;
        src106 <= 16'hc37e;
        src107 <= 16'h1452;
        src108 <= 16'hfc2b;
        src109 <= 16'hec54;
        src110 <= 16'h1d8a;
        src111 <= 16'h58d7;
        src112 <= 16'h54d5;
        src113 <= 16'hb32c;
        src114 <= 16'h72c8;
        src115 <= 16'h6799;
        src116 <= 16'hdc00;
        src117 <= 16'h4fdb;
        src118 <= 16'h2894;
        src119 <= 16'h5a71;
        src120 <= 16'h531d;
        src121 <= 16'h7057;
        src122 <= 16'hfeb3;
        src123 <= 16'h9c41;
        src124 <= 16'ha03b;
        src125 <= 16'hf54a;
        src126 <= 16'hbf30;
        src127 <= 16'hf76f;
        src128 <= 16'hb869;
        src129 <= 16'he0fa;
        src130 <= 16'h3977;
        src131 <= 16'hb065;
        src132 <= 16'hfd8d;
        src133 <= 16'h464a;
        src134 <= 16'hb4e9;
        src135 <= 16'h97a5;
        src136 <= 16'h8e45;
        src137 <= 16'h4b0;
        src138 <= 16'h91a3;
        src139 <= 16'h9401;
        src140 <= 16'h636e;
        src141 <= 16'h9edf;
        src142 <= 16'h851a;
        src143 <= 16'h6ba;
        src144 <= 16'heaba;
        src145 <= 16'hd6d6;
        src146 <= 16'h7677;
        src147 <= 16'hf40d;
        src148 <= 16'h7efb;
        src149 <= 16'hb209;
        src150 <= 16'h2b5;
        src151 <= 16'hcb72;
        src152 <= 16'ha02c;
        src153 <= 16'h93da;
        src154 <= 16'h5bba;
        src155 <= 16'h1c94;
        src156 <= 16'h5c4b;
        src157 <= 16'ha8d6;
        src158 <= 16'h19a4;
        src159 <= 16'hca40;
        src160 <= 16'he46a;
        src161 <= 16'ha6bf;
        src162 <= 16'hd432;
        src163 <= 16'h56df;
        src164 <= 16'he14e;
        src165 <= 16'hb5d2;
        src166 <= 16'h538a;
        src167 <= 16'h8338;
        src168 <= 16'hcb94;
        src169 <= 16'h51b8;
        src170 <= 16'h565f;
        src171 <= 16'h3ac5;
        src172 <= 16'h8b97;
        src173 <= 16'hdeea;
        src174 <= 16'hd805;
        src175 <= 16'hf71d;
        src176 <= 16'h5c87;
        src177 <= 16'h6f97;
        src178 <= 16'h85ec;
        src179 <= 16'hfd62;
        src180 <= 16'hd5ce;
        src181 <= 16'h8336;
        src182 <= 16'h659;
        src183 <= 16'hd10a;
        src184 <= 16'h861;
        exp <= 24'h5c29e9;
        #1
        src0 <= 16'hfb47;
        src1 <= 16'h44c0;
        src2 <= 16'h243f;
        src3 <= 16'hcfba;
        src4 <= 16'hfd61;
        src5 <= 16'ha3b5;
        src6 <= 16'hde3f;
        src7 <= 16'h7149;
        src8 <= 16'he63d;
        src9 <= 16'h7691;
        src10 <= 16'hfe4;
        src11 <= 16'h421f;
        src12 <= 16'ha0e2;
        src13 <= 16'hd206;
        src14 <= 16'h3882;
        src15 <= 16'hcc33;
        src16 <= 16'hc5d6;
        src17 <= 16'h27ae;
        src18 <= 16'h185a;
        src19 <= 16'h9f51;
        src20 <= 16'hdecc;
        src21 <= 16'h6363;
        src22 <= 16'h90a6;
        src23 <= 16'h7847;
        src24 <= 16'h2c24;
        src25 <= 16'he207;
        src26 <= 16'h2040;
        src27 <= 16'h8c12;
        src28 <= 16'h5dde;
        src29 <= 16'hc2f8;
        src30 <= 16'ha030;
        src31 <= 16'hcdfb;
        src32 <= 16'h2d09;
        src33 <= 16'h7795;
        src34 <= 16'hcb1f;
        src35 <= 16'h344b;
        src36 <= 16'h5d68;
        src37 <= 16'he76d;
        src38 <= 16'h44b6;
        src39 <= 16'hb806;
        src40 <= 16'h5108;
        src41 <= 16'hfcf2;
        src42 <= 16'hd0f9;
        src43 <= 16'he0e2;
        src44 <= 16'h379f;
        src45 <= 16'he707;
        src46 <= 16'hba8d;
        src47 <= 16'heeba;
        src48 <= 16'h32a4;
        src49 <= 16'hb58;
        src50 <= 16'h8815;
        src51 <= 16'h727f;
        src52 <= 16'hf988;
        src53 <= 16'h8837;
        src54 <= 16'h7289;
        src55 <= 16'hd8b4;
        src56 <= 16'hc57b;
        src57 <= 16'hbdbf;
        src58 <= 16'h913c;
        src59 <= 16'ha720;
        src60 <= 16'hee60;
        src61 <= 16'ha0a0;
        src62 <= 16'hbb99;
        src63 <= 16'h395c;
        src64 <= 16'hcce2;
        src65 <= 16'h594;
        src66 <= 16'haa11;
        src67 <= 16'h4e44;
        src68 <= 16'h85f4;
        src69 <= 16'h4408;
        src70 <= 16'h9566;
        src71 <= 16'h8529;
        src72 <= 16'h240c;
        src73 <= 16'h8246;
        src74 <= 16'hc993;
        src75 <= 16'h6c47;
        src76 <= 16'h17fa;
        src77 <= 16'h8f64;
        src78 <= 16'h5778;
        src79 <= 16'h1a32;
        src80 <= 16'h6fd2;
        src81 <= 16'ha6e6;
        src82 <= 16'hd3b0;
        src83 <= 16'hfbdd;
        src84 <= 16'h176d;
        src85 <= 16'hbe2;
        src86 <= 16'h9dc9;
        src87 <= 16'he9a2;
        src88 <= 16'h5471;
        src89 <= 16'hbcf1;
        src90 <= 16'h407b;
        src91 <= 16'h83fe;
        src92 <= 16'hee46;
        src93 <= 16'hcb7d;
        src94 <= 16'h2b5;
        src95 <= 16'he6cf;
        src96 <= 16'h93e4;
        src97 <= 16'h3d7e;
        src98 <= 16'hbc60;
        src99 <= 16'h5b76;
        src100 <= 16'h248f;
        src101 <= 16'hfe99;
        src102 <= 16'h358e;
        src103 <= 16'h10f7;
        src104 <= 16'hb64d;
        src105 <= 16'hef83;
        src106 <= 16'h71b7;
        src107 <= 16'h2a78;
        src108 <= 16'ha035;
        src109 <= 16'he4df;
        src110 <= 16'h67b;
        src111 <= 16'h7961;
        src112 <= 16'he58;
        src113 <= 16'h3425;
        src114 <= 16'h4823;
        src115 <= 16'h665c;
        src116 <= 16'h1ea2;
        src117 <= 16'hbfec;
        src118 <= 16'hd2fa;
        src119 <= 16'h500f;
        src120 <= 16'h1101;
        src121 <= 16'h3a5f;
        src122 <= 16'h115e;
        src123 <= 16'hce6c;
        src124 <= 16'h5aa;
        src125 <= 16'hf4d;
        src126 <= 16'h7b77;
        src127 <= 16'h7a6e;
        src128 <= 16'hd534;
        src129 <= 16'h128c;
        src130 <= 16'ha6cd;
        src131 <= 16'hbbd0;
        src132 <= 16'h4943;
        src133 <= 16'hf7cd;
        src134 <= 16'hbdd9;
        src135 <= 16'h3866;
        src136 <= 16'h9031;
        src137 <= 16'h97db;
        src138 <= 16'haf32;
        src139 <= 16'h1e8a;
        src140 <= 16'h78e;
        src141 <= 16'h2e81;
        src142 <= 16'hd434;
        src143 <= 16'h82bb;
        src144 <= 16'h415d;
        src145 <= 16'hc65d;
        src146 <= 16'h2c50;
        src147 <= 16'h49b;
        src148 <= 16'hd087;
        src149 <= 16'h7512;
        src150 <= 16'hd272;
        src151 <= 16'h3ca6;
        src152 <= 16'hb8df;
        src153 <= 16'h76c3;
        src154 <= 16'h63f9;
        src155 <= 16'h28a6;
        src156 <= 16'h3980;
        src157 <= 16'hed38;
        src158 <= 16'h8dec;
        src159 <= 16'h3efb;
        src160 <= 16'h1083;
        src161 <= 16'hca10;
        src162 <= 16'hf3ee;
        src163 <= 16'h890f;
        src164 <= 16'h8784;
        src165 <= 16'hb649;
        src166 <= 16'hbbd0;
        src167 <= 16'habd5;
        src168 <= 16'h92e3;
        src169 <= 16'h2cf0;
        src170 <= 16'h579a;
        src171 <= 16'h4ec4;
        src172 <= 16'hd4df;
        src173 <= 16'hfb7b;
        src174 <= 16'h6d66;
        src175 <= 16'hc7e8;
        src176 <= 16'h74ef;
        src177 <= 16'haa02;
        src178 <= 16'hbfdc;
        src179 <= 16'h12e4;
        src180 <= 16'h566;
        src181 <= 16'h38f0;
        src182 <= 16'h4ccf;
        src183 <= 16'ha0b4;
        src184 <= 16'h2faf;
        exp <= 24'h5ce01b;
        #1
        src0 <= 16'h9520;
        src1 <= 16'h39b5;
        src2 <= 16'h8bd0;
        src3 <= 16'h372f;
        src4 <= 16'hf4f2;
        src5 <= 16'h5265;
        src6 <= 16'hc1d5;
        src7 <= 16'h8fac;
        src8 <= 16'hbd48;
        src9 <= 16'hbf0b;
        src10 <= 16'haf4d;
        src11 <= 16'h1b98;
        src12 <= 16'h974e;
        src13 <= 16'h280a;
        src14 <= 16'h33ed;
        src15 <= 16'habad;
        src16 <= 16'h931f;
        src17 <= 16'h646;
        src18 <= 16'h60dd;
        src19 <= 16'h1e5d;
        src20 <= 16'haeaa;
        src21 <= 16'hc8f3;
        src22 <= 16'h5eac;
        src23 <= 16'ha992;
        src24 <= 16'h46e9;
        src25 <= 16'h16aa;
        src26 <= 16'hd9e5;
        src27 <= 16'h1e91;
        src28 <= 16'h6f25;
        src29 <= 16'hd8f9;
        src30 <= 16'h954d;
        src31 <= 16'hb043;
        src32 <= 16'h25f7;
        src33 <= 16'h6bb8;
        src34 <= 16'h7980;
        src35 <= 16'heea6;
        src36 <= 16'hfd38;
        src37 <= 16'h75d2;
        src38 <= 16'h385f;
        src39 <= 16'had78;
        src40 <= 16'h28e4;
        src41 <= 16'hd616;
        src42 <= 16'h1205;
        src43 <= 16'h8000;
        src44 <= 16'h64f7;
        src45 <= 16'h8e62;
        src46 <= 16'h2d9f;
        src47 <= 16'hcdbd;
        src48 <= 16'h24b7;
        src49 <= 16'h88a6;
        src50 <= 16'hb220;
        src51 <= 16'hadc1;
        src52 <= 16'h2d09;
        src53 <= 16'h30dd;
        src54 <= 16'hb68c;
        src55 <= 16'hde98;
        src56 <= 16'hed8d;
        src57 <= 16'hcda0;
        src58 <= 16'h9ec2;
        src59 <= 16'h63e1;
        src60 <= 16'hf902;
        src61 <= 16'hfe54;
        src62 <= 16'h70ad;
        src63 <= 16'h24ad;
        src64 <= 16'had2b;
        src65 <= 16'h10bf;
        src66 <= 16'h15e4;
        src67 <= 16'hca20;
        src68 <= 16'h3589;
        src69 <= 16'he57d;
        src70 <= 16'hcb3c;
        src71 <= 16'h4e;
        src72 <= 16'h55f7;
        src73 <= 16'h357c;
        src74 <= 16'h96d6;
        src75 <= 16'h7626;
        src76 <= 16'hd382;
        src77 <= 16'h4873;
        src78 <= 16'h3b1f;
        src79 <= 16'hf2c;
        src80 <= 16'h1d71;
        src81 <= 16'h80c9;
        src82 <= 16'h6fdc;
        src83 <= 16'hc883;
        src84 <= 16'hff05;
        src85 <= 16'h3d89;
        src86 <= 16'hb056;
        src87 <= 16'ha219;
        src88 <= 16'h1730;
        src89 <= 16'h186e;
        src90 <= 16'h51b0;
        src91 <= 16'h3264;
        src92 <= 16'hf9d1;
        src93 <= 16'h12e8;
        src94 <= 16'hc083;
        src95 <= 16'hdb79;
        src96 <= 16'hb54b;
        src97 <= 16'h33c3;
        src98 <= 16'h303b;
        src99 <= 16'hfc04;
        src100 <= 16'hf6c2;
        src101 <= 16'h2b87;
        src102 <= 16'h6c1a;
        src103 <= 16'hdfd2;
        src104 <= 16'h7848;
        src105 <= 16'h96f6;
        src106 <= 16'h72e2;
        src107 <= 16'h8b38;
        src108 <= 16'h496d;
        src109 <= 16'h3d35;
        src110 <= 16'h285;
        src111 <= 16'h83cd;
        src112 <= 16'ha076;
        src113 <= 16'he73e;
        src114 <= 16'h3010;
        src115 <= 16'hd875;
        src116 <= 16'ha2a;
        src117 <= 16'hb06a;
        src118 <= 16'hae54;
        src119 <= 16'h5fe4;
        src120 <= 16'ha64;
        src121 <= 16'h4159;
        src122 <= 16'h9455;
        src123 <= 16'h57ed;
        src124 <= 16'hb544;
        src125 <= 16'h1aca;
        src126 <= 16'ha693;
        src127 <= 16'hc1ca;
        src128 <= 16'h1d0b;
        src129 <= 16'h2b03;
        src130 <= 16'ha7e5;
        src131 <= 16'hc31d;
        src132 <= 16'h173f;
        src133 <= 16'ha26b;
        src134 <= 16'h4fc3;
        src135 <= 16'hdcdc;
        src136 <= 16'hf140;
        src137 <= 16'h2f1;
        src138 <= 16'h4172;
        src139 <= 16'h34fb;
        src140 <= 16'h25d9;
        src141 <= 16'h5c72;
        src142 <= 16'hec05;
        src143 <= 16'h6692;
        src144 <= 16'h7068;
        src145 <= 16'h6ea5;
        src146 <= 16'h2be6;
        src147 <= 16'h5983;
        src148 <= 16'h2a09;
        src149 <= 16'hb46f;
        src150 <= 16'h21ae;
        src151 <= 16'h4a3e;
        src152 <= 16'h161f;
        src153 <= 16'hcafa;
        src154 <= 16'h86ba;
        src155 <= 16'h3ad7;
        src156 <= 16'hec37;
        src157 <= 16'heff;
        src158 <= 16'ha9b;
        src159 <= 16'h7806;
        src160 <= 16'hab31;
        src161 <= 16'hd4fb;
        src162 <= 16'h5c86;
        src163 <= 16'h8442;
        src164 <= 16'h64f0;
        src165 <= 16'h3370;
        src166 <= 16'h9126;
        src167 <= 16'h9d16;
        src168 <= 16'h48c0;
        src169 <= 16'hfd9a;
        src170 <= 16'h7dc2;
        src171 <= 16'h2676;
        src172 <= 16'h3138;
        src173 <= 16'h1de7;
        src174 <= 16'hfbf1;
        src175 <= 16'h8eb9;
        src176 <= 16'hdf6;
        src177 <= 16'hdc73;
        src178 <= 16'hea0;
        src179 <= 16'hf82a;
        src180 <= 16'h4f55;
        src181 <= 16'ha827;
        src182 <= 16'h7871;
        src183 <= 16'h35f5;
        src184 <= 16'h1e4f;
        exp <= 24'h56a023;
        #1
        src0 <= 16'hb930;
        src1 <= 16'hfa44;
        src2 <= 16'hee59;
        src3 <= 16'h42e0;
        src4 <= 16'hc9cd;
        src5 <= 16'hf353;
        src6 <= 16'hb84a;
        src7 <= 16'he040;
        src8 <= 16'hbe02;
        src9 <= 16'h8da3;
        src10 <= 16'h620d;
        src11 <= 16'h5fb1;
        src12 <= 16'h431;
        src13 <= 16'h5e9d;
        src14 <= 16'hc2c3;
        src15 <= 16'h2822;
        src16 <= 16'h5412;
        src17 <= 16'hb1de;
        src18 <= 16'h8447;
        src19 <= 16'h1820;
        src20 <= 16'h8c8f;
        src21 <= 16'h405a;
        src22 <= 16'h4e8f;
        src23 <= 16'h510f;
        src24 <= 16'h4d8a;
        src25 <= 16'h5153;
        src26 <= 16'haab;
        src27 <= 16'h31f0;
        src28 <= 16'h3b86;
        src29 <= 16'h9ebd;
        src30 <= 16'he272;
        src31 <= 16'h23d4;
        src32 <= 16'hb4eb;
        src33 <= 16'hb7e5;
        src34 <= 16'h222e;
        src35 <= 16'hf4a5;
        src36 <= 16'hd5f3;
        src37 <= 16'h4c0d;
        src38 <= 16'h3190;
        src39 <= 16'h2259;
        src40 <= 16'hb8b5;
        src41 <= 16'hea8b;
        src42 <= 16'h3b83;
        src43 <= 16'h53a2;
        src44 <= 16'h578d;
        src45 <= 16'hf77;
        src46 <= 16'hd52e;
        src47 <= 16'h3228;
        src48 <= 16'hb3cb;
        src49 <= 16'h715a;
        src50 <= 16'h4bdf;
        src51 <= 16'h6981;
        src52 <= 16'h1707;
        src53 <= 16'hc073;
        src54 <= 16'h2397;
        src55 <= 16'h1e88;
        src56 <= 16'h82d1;
        src57 <= 16'h9eb8;
        src58 <= 16'h367e;
        src59 <= 16'h5de2;
        src60 <= 16'h28cd;
        src61 <= 16'h2514;
        src62 <= 16'hfd89;
        src63 <= 16'hebb1;
        src64 <= 16'hfe5d;
        src65 <= 16'h21bc;
        src66 <= 16'he27d;
        src67 <= 16'h8ae1;
        src68 <= 16'h1c31;
        src69 <= 16'h7e37;
        src70 <= 16'hf0d7;
        src71 <= 16'h8699;
        src72 <= 16'h499e;
        src73 <= 16'h6acd;
        src74 <= 16'h2611;
        src75 <= 16'h40a0;
        src76 <= 16'h8ff;
        src77 <= 16'h6107;
        src78 <= 16'h6be9;
        src79 <= 16'h73b9;
        src80 <= 16'h419b;
        src81 <= 16'hf607;
        src82 <= 16'h47d2;
        src83 <= 16'h2ff1;
        src84 <= 16'h921f;
        src85 <= 16'h8953;
        src86 <= 16'h27bc;
        src87 <= 16'h681b;
        src88 <= 16'hcd69;
        src89 <= 16'hd07;
        src90 <= 16'h716e;
        src91 <= 16'h911c;
        src92 <= 16'h142c;
        src93 <= 16'h4c98;
        src94 <= 16'h823f;
        src95 <= 16'h47c3;
        src96 <= 16'h1ac2;
        src97 <= 16'hdecf;
        src98 <= 16'hcc4d;
        src99 <= 16'h67bb;
        src100 <= 16'ha4f1;
        src101 <= 16'h3aef;
        src102 <= 16'hc67d;
        src103 <= 16'h1756;
        src104 <= 16'h33cc;
        src105 <= 16'h70a7;
        src106 <= 16'h337;
        src107 <= 16'h3ea0;
        src108 <= 16'h2928;
        src109 <= 16'heb4a;
        src110 <= 16'h9944;
        src111 <= 16'h8a37;
        src112 <= 16'h253b;
        src113 <= 16'h6944;
        src114 <= 16'hbf;
        src115 <= 16'h2d9;
        src116 <= 16'hebae;
        src117 <= 16'h9b9c;
        src118 <= 16'h9aaf;
        src119 <= 16'ha4eb;
        src120 <= 16'h75fa;
        src121 <= 16'h4c6e;
        src122 <= 16'h4d48;
        src123 <= 16'h35f6;
        src124 <= 16'h524b;
        src125 <= 16'hb89e;
        src126 <= 16'h2f90;
        src127 <= 16'h9aa1;
        src128 <= 16'hfd98;
        src129 <= 16'hb878;
        src130 <= 16'h220a;
        src131 <= 16'h27b6;
        src132 <= 16'h46a;
        src133 <= 16'h7828;
        src134 <= 16'h2d41;
        src135 <= 16'hb072;
        src136 <= 16'h6aae;
        src137 <= 16'h4dbd;
        src138 <= 16'hae45;
        src139 <= 16'h349e;
        src140 <= 16'ha297;
        src141 <= 16'h75c9;
        src142 <= 16'hdbf5;
        src143 <= 16'hae30;
        src144 <= 16'h708d;
        src145 <= 16'hbbe3;
        src146 <= 16'hf530;
        src147 <= 16'ha569;
        src148 <= 16'h6616;
        src149 <= 16'h1506;
        src150 <= 16'h3cb;
        src151 <= 16'hcdb1;
        src152 <= 16'h6190;
        src153 <= 16'h922e;
        src154 <= 16'h2397;
        src155 <= 16'h638c;
        src156 <= 16'h1fff;
        src157 <= 16'h5056;
        src158 <= 16'hac6a;
        src159 <= 16'h1fa3;
        src160 <= 16'hc81a;
        src161 <= 16'h7b8f;
        src162 <= 16'he4b;
        src163 <= 16'h6ea0;
        src164 <= 16'hdd2c;
        src165 <= 16'hee6e;
        src166 <= 16'h17a0;
        src167 <= 16'hd408;
        src168 <= 16'h586c;
        src169 <= 16'h5ad6;
        src170 <= 16'hdb5e;
        src171 <= 16'h5ca6;
        src172 <= 16'h8450;
        src173 <= 16'h2528;
        src174 <= 16'h6632;
        src175 <= 16'hc9a3;
        src176 <= 16'h19ae;
        src177 <= 16'h31b6;
        src178 <= 16'h348d;
        src179 <= 16'he205;
        src180 <= 16'h884a;
        src181 <= 16'h1cc1;
        src182 <= 16'h2947;
        src183 <= 16'h9feb;
        src184 <= 16'h5912;
        exp <= 24'h5287f2;
        #1
        src0 <= 16'h501a;
        src1 <= 16'h9e4d;
        src2 <= 16'h9d47;
        src3 <= 16'hd831;
        src4 <= 16'hb617;
        src5 <= 16'h6189;
        src6 <= 16'h77a2;
        src7 <= 16'hb81e;
        src8 <= 16'hb65;
        src9 <= 16'hd954;
        src10 <= 16'had30;
        src11 <= 16'he17a;
        src12 <= 16'h3d84;
        src13 <= 16'h6ef0;
        src14 <= 16'hca46;
        src15 <= 16'hbccd;
        src16 <= 16'h84b7;
        src17 <= 16'hda6b;
        src18 <= 16'h12d6;
        src19 <= 16'hb5f2;
        src20 <= 16'h7a86;
        src21 <= 16'h7d34;
        src22 <= 16'h4ecf;
        src23 <= 16'h1404;
        src24 <= 16'h4637;
        src25 <= 16'h8a3d;
        src26 <= 16'hc5c9;
        src27 <= 16'h5b67;
        src28 <= 16'h5618;
        src29 <= 16'he495;
        src30 <= 16'h1fc0;
        src31 <= 16'h61e8;
        src32 <= 16'hcce4;
        src33 <= 16'hdeda;
        src34 <= 16'h9df0;
        src35 <= 16'h6568;
        src36 <= 16'h5955;
        src37 <= 16'h1178;
        src38 <= 16'h9e7a;
        src39 <= 16'h9cdb;
        src40 <= 16'h99;
        src41 <= 16'h98e3;
        src42 <= 16'h4821;
        src43 <= 16'hfec1;
        src44 <= 16'ha076;
        src45 <= 16'hb170;
        src46 <= 16'h8db6;
        src47 <= 16'hd9ff;
        src48 <= 16'hc8f5;
        src49 <= 16'hb2fb;
        src50 <= 16'h368f;
        src51 <= 16'h62fc;
        src52 <= 16'hd7e1;
        src53 <= 16'hb444;
        src54 <= 16'h6f88;
        src55 <= 16'hbbcd;
        src56 <= 16'h33d5;
        src57 <= 16'h8f59;
        src58 <= 16'he5dd;
        src59 <= 16'h127;
        src60 <= 16'h22e5;
        src61 <= 16'h24ba;
        src62 <= 16'h1f3e;
        src63 <= 16'h580e;
        src64 <= 16'h3928;
        src65 <= 16'h53c;
        src66 <= 16'hd6d4;
        src67 <= 16'h1384;
        src68 <= 16'hcd5c;
        src69 <= 16'ha00b;
        src70 <= 16'ha970;
        src71 <= 16'hebfe;
        src72 <= 16'hffb8;
        src73 <= 16'hce3d;
        src74 <= 16'h5294;
        src75 <= 16'heef9;
        src76 <= 16'haa05;
        src77 <= 16'h27ea;
        src78 <= 16'h1961;
        src79 <= 16'h70f5;
        src80 <= 16'h3a8b;
        src81 <= 16'hd971;
        src82 <= 16'h35a5;
        src83 <= 16'h9afe;
        src84 <= 16'h2c93;
        src85 <= 16'h192;
        src86 <= 16'h60a7;
        src87 <= 16'hfe9c;
        src88 <= 16'hc7f7;
        src89 <= 16'he6b8;
        src90 <= 16'hb68e;
        src91 <= 16'h7d8a;
        src92 <= 16'ha5ae;
        src93 <= 16'h6daf;
        src94 <= 16'hadd9;
        src95 <= 16'h36d3;
        src96 <= 16'h32f4;
        src97 <= 16'h87d1;
        src98 <= 16'hf717;
        src99 <= 16'h26a1;
        src100 <= 16'h4f1f;
        src101 <= 16'hd5b1;
        src102 <= 16'hd922;
        src103 <= 16'h9e79;
        src104 <= 16'h960f;
        src105 <= 16'h42;
        src106 <= 16'hb781;
        src107 <= 16'hae70;
        src108 <= 16'habc0;
        src109 <= 16'hcf4e;
        src110 <= 16'hd8d9;
        src111 <= 16'h8790;
        src112 <= 16'ha9fe;
        src113 <= 16'h1e99;
        src114 <= 16'h4d68;
        src115 <= 16'h1c1b;
        src116 <= 16'hae5f;
        src117 <= 16'h991c;
        src118 <= 16'ha043;
        src119 <= 16'h6852;
        src120 <= 16'h9f37;
        src121 <= 16'h75aa;
        src122 <= 16'h4193;
        src123 <= 16'h1e4f;
        src124 <= 16'hc857;
        src125 <= 16'h2d17;
        src126 <= 16'h4c5b;
        src127 <= 16'hbce4;
        src128 <= 16'h13;
        src129 <= 16'h63ac;
        src130 <= 16'h95c5;
        src131 <= 16'h1027;
        src132 <= 16'h4d02;
        src133 <= 16'he8fd;
        src134 <= 16'hef7d;
        src135 <= 16'hca4c;
        src136 <= 16'h146;
        src137 <= 16'hef4f;
        src138 <= 16'h58a3;
        src139 <= 16'hb64e;
        src140 <= 16'h3eec;
        src141 <= 16'he4e7;
        src142 <= 16'h191b;
        src143 <= 16'hab64;
        src144 <= 16'ha045;
        src145 <= 16'h8478;
        src146 <= 16'hdb19;
        src147 <= 16'h2e65;
        src148 <= 16'h5f70;
        src149 <= 16'h7b0b;
        src150 <= 16'hcc91;
        src151 <= 16'h229;
        src152 <= 16'h8670;
        src153 <= 16'h56d7;
        src154 <= 16'h3a20;
        src155 <= 16'h941a;
        src156 <= 16'h6d74;
        src157 <= 16'hab8e;
        src158 <= 16'hab0c;
        src159 <= 16'h7afe;
        src160 <= 16'he119;
        src161 <= 16'h217b;
        src162 <= 16'heec9;
        src163 <= 16'ha349;
        src164 <= 16'hec;
        src165 <= 16'haa71;
        src166 <= 16'h3628;
        src167 <= 16'h589f;
        src168 <= 16'hfe01;
        src169 <= 16'hed9b;
        src170 <= 16'h6520;
        src171 <= 16'haff8;
        src172 <= 16'h54c9;
        src173 <= 16'h6e78;
        src174 <= 16'hcf;
        src175 <= 16'he35c;
        src176 <= 16'h6b0a;
        src177 <= 16'hf671;
        src178 <= 16'hba87;
        src179 <= 16'h18e8;
        src180 <= 16'h8ab2;
        src181 <= 16'hb481;
        src182 <= 16'h9ccc;
        src183 <= 16'hc8c9;
        src184 <= 16'h350d;
        exp <= 24'h5ef737;
        #1
        src0 <= 16'h2142;
        src1 <= 16'h7bef;
        src2 <= 16'hb9f5;
        src3 <= 16'h1f4c;
        src4 <= 16'he618;
        src5 <= 16'h7ac5;
        src6 <= 16'hf4f;
        src7 <= 16'hc328;
        src8 <= 16'h8d6a;
        src9 <= 16'h6018;
        src10 <= 16'ha3bf;
        src11 <= 16'h3a5f;
        src12 <= 16'h26d8;
        src13 <= 16'h54f5;
        src14 <= 16'h16c6;
        src15 <= 16'ha737;
        src16 <= 16'hbfbc;
        src17 <= 16'h5b13;
        src18 <= 16'h7f1e;
        src19 <= 16'h6db7;
        src20 <= 16'h6173;
        src21 <= 16'h6b50;
        src22 <= 16'h31c1;
        src23 <= 16'he0d4;
        src24 <= 16'h2f6c;
        src25 <= 16'h2d84;
        src26 <= 16'ha8dd;
        src27 <= 16'h670d;
        src28 <= 16'h626c;
        src29 <= 16'h927e;
        src30 <= 16'h848a;
        src31 <= 16'h6661;
        src32 <= 16'h9e7f;
        src33 <= 16'h4505;
        src34 <= 16'h6e61;
        src35 <= 16'hda77;
        src36 <= 16'hbc3b;
        src37 <= 16'h72c0;
        src38 <= 16'ha08b;
        src39 <= 16'hff0f;
        src40 <= 16'h8808;
        src41 <= 16'hcf45;
        src42 <= 16'hc64c;
        src43 <= 16'he1aa;
        src44 <= 16'h33d6;
        src45 <= 16'hc0a8;
        src46 <= 16'h854f;
        src47 <= 16'h24e3;
        src48 <= 16'hf3fe;
        src49 <= 16'hc8e0;
        src50 <= 16'ha7b8;
        src51 <= 16'h50a5;
        src52 <= 16'he7d7;
        src53 <= 16'h3f5e;
        src54 <= 16'hb7f3;
        src55 <= 16'h3f2d;
        src56 <= 16'hc2aa;
        src57 <= 16'h2160;
        src58 <= 16'hb7ed;
        src59 <= 16'hc4f9;
        src60 <= 16'hcada;
        src61 <= 16'hee8;
        src62 <= 16'h210e;
        src63 <= 16'h5bc;
        src64 <= 16'h2778;
        src65 <= 16'h74f6;
        src66 <= 16'he8cb;
        src67 <= 16'hece6;
        src68 <= 16'haef2;
        src69 <= 16'h23d;
        src70 <= 16'h775a;
        src71 <= 16'hc615;
        src72 <= 16'he00b;
        src73 <= 16'hf704;
        src74 <= 16'h165f;
        src75 <= 16'hdb4d;
        src76 <= 16'h4e6b;
        src77 <= 16'h3f2e;
        src78 <= 16'h7448;
        src79 <= 16'h1055;
        src80 <= 16'h2a26;
        src81 <= 16'hfdb8;
        src82 <= 16'h7d97;
        src83 <= 16'h3b50;
        src84 <= 16'h3902;
        src85 <= 16'ha8f5;
        src86 <= 16'h17d2;
        src87 <= 16'hd36d;
        src88 <= 16'hec5a;
        src89 <= 16'he845;
        src90 <= 16'h5574;
        src91 <= 16'h8db8;
        src92 <= 16'heee6;
        src93 <= 16'ha807;
        src94 <= 16'h55c6;
        src95 <= 16'h6759;
        src96 <= 16'hea83;
        src97 <= 16'h9f3e;
        src98 <= 16'h57ec;
        src99 <= 16'h64b;
        src100 <= 16'hfd51;
        src101 <= 16'h7230;
        src102 <= 16'h5b2d;
        src103 <= 16'he1f0;
        src104 <= 16'hf0d1;
        src105 <= 16'h4608;
        src106 <= 16'hcac0;
        src107 <= 16'h4291;
        src108 <= 16'h1fcf;
        src109 <= 16'h1fcf;
        src110 <= 16'h42c1;
        src111 <= 16'h24a;
        src112 <= 16'h8a66;
        src113 <= 16'h64d3;
        src114 <= 16'h5a8e;
        src115 <= 16'h7ba9;
        src116 <= 16'h2bf;
        src117 <= 16'h9c41;
        src118 <= 16'h7ede;
        src119 <= 16'hf6a8;
        src120 <= 16'h12c0;
        src121 <= 16'h60a5;
        src122 <= 16'h4545;
        src123 <= 16'hdb50;
        src124 <= 16'hf31c;
        src125 <= 16'hb82e;
        src126 <= 16'h3487;
        src127 <= 16'h3813;
        src128 <= 16'h7c08;
        src129 <= 16'hc248;
        src130 <= 16'h9573;
        src131 <= 16'h1c47;
        src132 <= 16'hfd04;
        src133 <= 16'hcdf2;
        src134 <= 16'h18f4;
        src135 <= 16'h4c0c;
        src136 <= 16'h1b56;
        src137 <= 16'hf25e;
        src138 <= 16'h89e4;
        src139 <= 16'h739a;
        src140 <= 16'hb5f5;
        src141 <= 16'h5430;
        src142 <= 16'hc6c5;
        src143 <= 16'hb9a2;
        src144 <= 16'hf0d8;
        src145 <= 16'h63a0;
        src146 <= 16'h5c73;
        src147 <= 16'hf00f;
        src148 <= 16'h752d;
        src149 <= 16'hb20f;
        src150 <= 16'h59b;
        src151 <= 16'hf7c2;
        src152 <= 16'h2e5c;
        src153 <= 16'h1ae9;
        src154 <= 16'h4179;
        src155 <= 16'hf338;
        src156 <= 16'h39e7;
        src157 <= 16'hb6c4;
        src158 <= 16'hd164;
        src159 <= 16'hc7db;
        src160 <= 16'h2efc;
        src161 <= 16'h489d;
        src162 <= 16'h423f;
        src163 <= 16'h1d78;
        src164 <= 16'h3678;
        src165 <= 16'hb4e6;
        src166 <= 16'h643f;
        src167 <= 16'h6016;
        src168 <= 16'ha24;
        src169 <= 16'h6d38;
        src170 <= 16'h2b6c;
        src171 <= 16'ha842;
        src172 <= 16'ha536;
        src173 <= 16'h8e31;
        src174 <= 16'h45cd;
        src175 <= 16'h3a78;
        src176 <= 16'hcf3b;
        src177 <= 16'h85e4;
        src178 <= 16'hc313;
        src179 <= 16'h2af3;
        src180 <= 16'hd696;
        src181 <= 16'hea49;
        src182 <= 16'h16e5;
        src183 <= 16'h4349;
        src184 <= 16'ha71f;
        exp <= 24'h5b97c3;
        #1
        src0 <= 16'h6b62;
        src1 <= 16'hda3b;
        src2 <= 16'h1794;
        src3 <= 16'hbb34;
        src4 <= 16'hee6b;
        src5 <= 16'h2626;
        src6 <= 16'hf745;
        src7 <= 16'he747;
        src8 <= 16'hfd1c;
        src9 <= 16'h5497;
        src10 <= 16'h120d;
        src11 <= 16'ha297;
        src12 <= 16'heb87;
        src13 <= 16'hf356;
        src14 <= 16'h6c44;
        src15 <= 16'hce91;
        src16 <= 16'h7d3;
        src17 <= 16'h3571;
        src18 <= 16'hade1;
        src19 <= 16'h3f1a;
        src20 <= 16'h22cf;
        src21 <= 16'h756a;
        src22 <= 16'h11df;
        src23 <= 16'hd5f2;
        src24 <= 16'h8453;
        src25 <= 16'h8647;
        src26 <= 16'hd6f9;
        src27 <= 16'hb03d;
        src28 <= 16'he819;
        src29 <= 16'hcaca;
        src30 <= 16'h97a9;
        src31 <= 16'h81c7;
        src32 <= 16'h6a02;
        src33 <= 16'h21d4;
        src34 <= 16'hd446;
        src35 <= 16'h6a80;
        src36 <= 16'h21a9;
        src37 <= 16'h27f7;
        src38 <= 16'h473a;
        src39 <= 16'h86c4;
        src40 <= 16'hc0e8;
        src41 <= 16'h1464;
        src42 <= 16'hfb48;
        src43 <= 16'hd9ff;
        src44 <= 16'h7528;
        src45 <= 16'h2f4a;
        src46 <= 16'h98a2;
        src47 <= 16'he28a;
        src48 <= 16'h6ca7;
        src49 <= 16'h9e05;
        src50 <= 16'h71af;
        src51 <= 16'h6946;
        src52 <= 16'h34cc;
        src53 <= 16'hdc2d;
        src54 <= 16'hcd45;
        src55 <= 16'h48f9;
        src56 <= 16'hefc6;
        src57 <= 16'h32ee;
        src58 <= 16'h6224;
        src59 <= 16'h8f3;
        src60 <= 16'h9630;
        src61 <= 16'hbf0a;
        src62 <= 16'h58bd;
        src63 <= 16'h2bec;
        src64 <= 16'h17be;
        src65 <= 16'h4308;
        src66 <= 16'h14f8;
        src67 <= 16'h6284;
        src68 <= 16'he9c8;
        src69 <= 16'hc4e0;
        src70 <= 16'h509d;
        src71 <= 16'h3fb6;
        src72 <= 16'h656d;
        src73 <= 16'hcfdd;
        src74 <= 16'hd373;
        src75 <= 16'h2dcf;
        src76 <= 16'h3ca6;
        src77 <= 16'h4b95;
        src78 <= 16'h43a3;
        src79 <= 16'h4948;
        src80 <= 16'hfc90;
        src81 <= 16'h5cf8;
        src82 <= 16'hbbed;
        src83 <= 16'h47ea;
        src84 <= 16'hb2eb;
        src85 <= 16'hb08b;
        src86 <= 16'ha480;
        src87 <= 16'h83d;
        src88 <= 16'h28c2;
        src89 <= 16'h4b38;
        src90 <= 16'h6900;
        src91 <= 16'h762d;
        src92 <= 16'h72f9;
        src93 <= 16'hc339;
        src94 <= 16'h5cf1;
        src95 <= 16'h670e;
        src96 <= 16'hbf8e;
        src97 <= 16'h3290;
        src98 <= 16'h987;
        src99 <= 16'h17eb;
        src100 <= 16'hfc4e;
        src101 <= 16'h828f;
        src102 <= 16'hb813;
        src103 <= 16'he2a1;
        src104 <= 16'h642d;
        src105 <= 16'hc320;
        src106 <= 16'hc56d;
        src107 <= 16'hcdaf;
        src108 <= 16'h8737;
        src109 <= 16'h6959;
        src110 <= 16'h87cb;
        src111 <= 16'h4f80;
        src112 <= 16'hff64;
        src113 <= 16'h3155;
        src114 <= 16'h4e55;
        src115 <= 16'h824;
        src116 <= 16'h873e;
        src117 <= 16'h105c;
        src118 <= 16'h3431;
        src119 <= 16'h8332;
        src120 <= 16'h6870;
        src121 <= 16'hb957;
        src122 <= 16'h1ff7;
        src123 <= 16'h32f;
        src124 <= 16'h938c;
        src125 <= 16'hd09;
        src126 <= 16'h3f10;
        src127 <= 16'ha36b;
        src128 <= 16'hfb9b;
        src129 <= 16'h8760;
        src130 <= 16'hf4ea;
        src131 <= 16'he3ac;
        src132 <= 16'hb5a5;
        src133 <= 16'h9424;
        src134 <= 16'hfce5;
        src135 <= 16'h38bd;
        src136 <= 16'h7bef;
        src137 <= 16'hab6b;
        src138 <= 16'h35b4;
        src139 <= 16'hc544;
        src140 <= 16'ha166;
        src141 <= 16'habdc;
        src142 <= 16'h2776;
        src143 <= 16'h267e;
        src144 <= 16'h1063;
        src145 <= 16'h9152;
        src146 <= 16'h9152;
        src147 <= 16'ha875;
        src148 <= 16'h3b;
        src149 <= 16'hf5fc;
        src150 <= 16'hddb2;
        src151 <= 16'h9094;
        src152 <= 16'hc1c6;
        src153 <= 16'h5edc;
        src154 <= 16'h2a79;
        src155 <= 16'h694;
        src156 <= 16'h6323;
        src157 <= 16'h6b60;
        src158 <= 16'h399c;
        src159 <= 16'hb024;
        src160 <= 16'h3d2;
        src161 <= 16'h576c;
        src162 <= 16'h6665;
        src163 <= 16'h3f67;
        src164 <= 16'h114e;
        src165 <= 16'ha73a;
        src166 <= 16'hb0d7;
        src167 <= 16'h4ce5;
        src168 <= 16'hf132;
        src169 <= 16'hb3ce;
        src170 <= 16'heebe;
        src171 <= 16'h22a4;
        src172 <= 16'he0fb;
        src173 <= 16'h7762;
        src174 <= 16'h1643;
        src175 <= 16'ha181;
        src176 <= 16'hb1a6;
        src177 <= 16'h3c65;
        src178 <= 16'hb153;
        src179 <= 16'hdf0a;
        src180 <= 16'h7fc8;
        src181 <= 16'h1c24;
        src182 <= 16'h159b;
        src183 <= 16'h91ff;
        src184 <= 16'hca11;
        exp <= 24'h5aa691;
        #1
        src0 <= 16'hb61e;
        src1 <= 16'h48a8;
        src2 <= 16'h3579;
        src3 <= 16'h7827;
        src4 <= 16'ha9fa;
        src5 <= 16'hc0f1;
        src6 <= 16'hc7e5;
        src7 <= 16'h697c;
        src8 <= 16'h311b;
        src9 <= 16'h5bc1;
        src10 <= 16'h3c94;
        src11 <= 16'h4dd5;
        src12 <= 16'h26fd;
        src13 <= 16'h63bc;
        src14 <= 16'hd21e;
        src15 <= 16'hba6f;
        src16 <= 16'hd02e;
        src17 <= 16'he6bc;
        src18 <= 16'h9b03;
        src19 <= 16'ha917;
        src20 <= 16'h82b4;
        src21 <= 16'h179f;
        src22 <= 16'hddad;
        src23 <= 16'h86d7;
        src24 <= 16'h116d;
        src25 <= 16'h2b16;
        src26 <= 16'h1f74;
        src27 <= 16'he13;
        src28 <= 16'h7277;
        src29 <= 16'hcb3b;
        src30 <= 16'hd718;
        src31 <= 16'h57c0;
        src32 <= 16'head;
        src33 <= 16'hf5d1;
        src34 <= 16'hee0b;
        src35 <= 16'h3680;
        src36 <= 16'h8ac8;
        src37 <= 16'h5caa;
        src38 <= 16'h5c4f;
        src39 <= 16'hf690;
        src40 <= 16'h1a1d;
        src41 <= 16'hc7a;
        src42 <= 16'hc62e;
        src43 <= 16'hda0;
        src44 <= 16'hbfec;
        src45 <= 16'h45a9;
        src46 <= 16'hb11b;
        src47 <= 16'h8813;
        src48 <= 16'h35c4;
        src49 <= 16'h93ff;
        src50 <= 16'h5c96;
        src51 <= 16'h99ce;
        src52 <= 16'hfbd9;
        src53 <= 16'h9298;
        src54 <= 16'hd183;
        src55 <= 16'h200;
        src56 <= 16'h97b6;
        src57 <= 16'hedf8;
        src58 <= 16'hba46;
        src59 <= 16'h5665;
        src60 <= 16'h25ac;
        src61 <= 16'h9087;
        src62 <= 16'hb244;
        src63 <= 16'h115b;
        src64 <= 16'h8f7f;
        src65 <= 16'h33bf;
        src66 <= 16'hd83d;
        src67 <= 16'h201;
        src68 <= 16'hbab2;
        src69 <= 16'h1b0c;
        src70 <= 16'h6e6a;
        src71 <= 16'hacd8;
        src72 <= 16'h9dc7;
        src73 <= 16'h9e7a;
        src74 <= 16'h5ba4;
        src75 <= 16'h90f0;
        src76 <= 16'h3737;
        src77 <= 16'hd4b4;
        src78 <= 16'h943a;
        src79 <= 16'h3d58;
        src80 <= 16'h7a6b;
        src81 <= 16'h1837;
        src82 <= 16'h6970;
        src83 <= 16'hcb7b;
        src84 <= 16'hf4a3;
        src85 <= 16'h10cb;
        src86 <= 16'h3f9b;
        src87 <= 16'h2754;
        src88 <= 16'hb39d;
        src89 <= 16'h4360;
        src90 <= 16'hbd8e;
        src91 <= 16'hddbe;
        src92 <= 16'h1a69;
        src93 <= 16'hd85b;
        src94 <= 16'h856b;
        src95 <= 16'hb634;
        src96 <= 16'h1ea7;
        src97 <= 16'he263;
        src98 <= 16'ha6c7;
        src99 <= 16'hf4e2;
        src100 <= 16'hd9d3;
        src101 <= 16'h9c92;
        src102 <= 16'h12ed;
        src103 <= 16'h153e;
        src104 <= 16'h89ff;
        src105 <= 16'h4c42;
        src106 <= 16'h4f91;
        src107 <= 16'h6c65;
        src108 <= 16'headd;
        src109 <= 16'h497b;
        src110 <= 16'hdd4b;
        src111 <= 16'h1f37;
        src112 <= 16'h1331;
        src113 <= 16'h1f7d;
        src114 <= 16'hb3d9;
        src115 <= 16'hd9ca;
        src116 <= 16'h221c;
        src117 <= 16'h3613;
        src118 <= 16'habf3;
        src119 <= 16'h7be3;
        src120 <= 16'ha158;
        src121 <= 16'ha203;
        src122 <= 16'h28a;
        src123 <= 16'h7835;
        src124 <= 16'haef6;
        src125 <= 16'h232c;
        src126 <= 16'h1e3b;
        src127 <= 16'hfb33;
        src128 <= 16'h27ed;
        src129 <= 16'hb7b6;
        src130 <= 16'h598a;
        src131 <= 16'hb7c0;
        src132 <= 16'hc427;
        src133 <= 16'h2cba;
        src134 <= 16'h4736;
        src135 <= 16'h753b;
        src136 <= 16'hfa11;
        src137 <= 16'h127e;
        src138 <= 16'h6a02;
        src139 <= 16'hdfe3;
        src140 <= 16'he86f;
        src141 <= 16'h15de;
        src142 <= 16'h7514;
        src143 <= 16'h6fe4;
        src144 <= 16'hcd22;
        src145 <= 16'hf5a5;
        src146 <= 16'hcc8;
        src147 <= 16'h72c6;
        src148 <= 16'hf95e;
        src149 <= 16'h1c3b;
        src150 <= 16'h71ae;
        src151 <= 16'hde26;
        src152 <= 16'h5de;
        src153 <= 16'h2d7a;
        src154 <= 16'hd4a8;
        src155 <= 16'h71fc;
        src156 <= 16'h5939;
        src157 <= 16'h1133;
        src158 <= 16'hc7bc;
        src159 <= 16'h40b7;
        src160 <= 16'h184a;
        src161 <= 16'h401c;
        src162 <= 16'ha11b;
        src163 <= 16'h2f2a;
        src164 <= 16'h381b;
        src165 <= 16'hdca8;
        src166 <= 16'hbd49;
        src167 <= 16'heec;
        src168 <= 16'h7007;
        src169 <= 16'h365;
        src170 <= 16'h5705;
        src171 <= 16'h1503;
        src172 <= 16'hf7a1;
        src173 <= 16'hdb9c;
        src174 <= 16'h8871;
        src175 <= 16'h307f;
        src176 <= 16'h9d8c;
        src177 <= 16'h8780;
        src178 <= 16'h4068;
        src179 <= 16'ha8aa;
        src180 <= 16'h84a;
        src181 <= 16'h934b;
        src182 <= 16'hd44c;
        src183 <= 16'h4831;
        src184 <= 16'hf8d;
        exp <= 24'h573fc2;
        #1
        src0 <= 16'hd862;
        src1 <= 16'h1b88;
        src2 <= 16'h973c;
        src3 <= 16'hdda3;
        src4 <= 16'h6df6;
        src5 <= 16'hdc3f;
        src6 <= 16'h2bfd;
        src7 <= 16'h52bc;
        src8 <= 16'h4aba;
        src9 <= 16'h7ed2;
        src10 <= 16'he029;
        src11 <= 16'hacec;
        src12 <= 16'haf15;
        src13 <= 16'h9627;
        src14 <= 16'h7821;
        src15 <= 16'hc829;
        src16 <= 16'h194a;
        src17 <= 16'h9d27;
        src18 <= 16'h474a;
        src19 <= 16'hf779;
        src20 <= 16'h6316;
        src21 <= 16'h545d;
        src22 <= 16'hb8a9;
        src23 <= 16'h1694;
        src24 <= 16'h414d;
        src25 <= 16'h6d96;
        src26 <= 16'h70b5;
        src27 <= 16'h51ba;
        src28 <= 16'h7018;
        src29 <= 16'h5278;
        src30 <= 16'h42e5;
        src31 <= 16'ha96a;
        src32 <= 16'h3cb5;
        src33 <= 16'h5da6;
        src34 <= 16'h3846;
        src35 <= 16'h7ea3;
        src36 <= 16'hb661;
        src37 <= 16'hee26;
        src38 <= 16'h863a;
        src39 <= 16'ha51;
        src40 <= 16'hd569;
        src41 <= 16'h57cc;
        src42 <= 16'h2326;
        src43 <= 16'hbf3e;
        src44 <= 16'h2965;
        src45 <= 16'h2d12;
        src46 <= 16'h3ac9;
        src47 <= 16'h3d88;
        src48 <= 16'hc882;
        src49 <= 16'h8762;
        src50 <= 16'h81ea;
        src51 <= 16'hc477;
        src52 <= 16'h4db8;
        src53 <= 16'h4661;
        src54 <= 16'h766a;
        src55 <= 16'h438e;
        src56 <= 16'hb6a4;
        src57 <= 16'h7f4c;
        src58 <= 16'h117d;
        src59 <= 16'hd010;
        src60 <= 16'h35e3;
        src61 <= 16'hfa19;
        src62 <= 16'h4506;
        src63 <= 16'hca86;
        src64 <= 16'h2679;
        src65 <= 16'h92da;
        src66 <= 16'h8c7b;
        src67 <= 16'h21a5;
        src68 <= 16'hfa82;
        src69 <= 16'hcaca;
        src70 <= 16'h2e7;
        src71 <= 16'h82f0;
        src72 <= 16'h6450;
        src73 <= 16'haaca;
        src74 <= 16'hb352;
        src75 <= 16'h8086;
        src76 <= 16'hbab5;
        src77 <= 16'hd1ff;
        src78 <= 16'hc9f9;
        src79 <= 16'ha2a8;
        src80 <= 16'hb359;
        src81 <= 16'h7db0;
        src82 <= 16'he57f;
        src83 <= 16'hfbb6;
        src84 <= 16'h3464;
        src85 <= 16'hb4f5;
        src86 <= 16'h9719;
        src87 <= 16'h9d05;
        src88 <= 16'h9c3c;
        src89 <= 16'hdc96;
        src90 <= 16'h143a;
        src91 <= 16'h9512;
        src92 <= 16'he067;
        src93 <= 16'h5f7b;
        src94 <= 16'hea43;
        src95 <= 16'h35e1;
        src96 <= 16'h1b92;
        src97 <= 16'h2999;
        src98 <= 16'he878;
        src99 <= 16'h14b2;
        src100 <= 16'h3d39;
        src101 <= 16'had67;
        src102 <= 16'hec25;
        src103 <= 16'h5131;
        src104 <= 16'h85e8;
        src105 <= 16'h92d8;
        src106 <= 16'hc1d9;
        src107 <= 16'h4599;
        src108 <= 16'h9b10;
        src109 <= 16'h9f7f;
        src110 <= 16'h5fe9;
        src111 <= 16'h9579;
        src112 <= 16'h698c;
        src113 <= 16'hc427;
        src114 <= 16'h5bef;
        src115 <= 16'h5fc9;
        src116 <= 16'h216a;
        src117 <= 16'h389e;
        src118 <= 16'hff66;
        src119 <= 16'h785e;
        src120 <= 16'h627c;
        src121 <= 16'hc13d;
        src122 <= 16'h3c5b;
        src123 <= 16'hcadb;
        src124 <= 16'h6a7e;
        src125 <= 16'h90ee;
        src126 <= 16'hfe21;
        src127 <= 16'h823e;
        src128 <= 16'h6eda;
        src129 <= 16'h7ea9;
        src130 <= 16'h3511;
        src131 <= 16'h6b19;
        src132 <= 16'hd4d7;
        src133 <= 16'h6f41;
        src134 <= 16'ha8e4;
        src135 <= 16'h6200;
        src136 <= 16'h6dd1;
        src137 <= 16'h2cf4;
        src138 <= 16'hbc57;
        src139 <= 16'ha662;
        src140 <= 16'h3f26;
        src141 <= 16'h64a8;
        src142 <= 16'h9548;
        src143 <= 16'h8cad;
        src144 <= 16'hf4aa;
        src145 <= 16'he0cb;
        src146 <= 16'hccde;
        src147 <= 16'hb163;
        src148 <= 16'hab20;
        src149 <= 16'h2a49;
        src150 <= 16'h813f;
        src151 <= 16'h2752;
        src152 <= 16'he9cb;
        src153 <= 16'hb846;
        src154 <= 16'hd026;
        src155 <= 16'h2c8b;
        src156 <= 16'h899c;
        src157 <= 16'h338e;
        src158 <= 16'h6c7d;
        src159 <= 16'hf5d1;
        src160 <= 16'h1161;
        src161 <= 16'h1c55;
        src162 <= 16'h498e;
        src163 <= 16'h9c4f;
        src164 <= 16'h2e45;
        src165 <= 16'h6b94;
        src166 <= 16'he103;
        src167 <= 16'h4d76;
        src168 <= 16'h3edb;
        src169 <= 16'h303b;
        src170 <= 16'h8a3;
        src171 <= 16'hba61;
        src172 <= 16'hc88e;
        src173 <= 16'h2d01;
        src174 <= 16'h9fbd;
        src175 <= 16'h5c7d;
        src176 <= 16'h4054;
        src177 <= 16'hbdf5;
        src178 <= 16'hc9e;
        src179 <= 16'ha46f;
        src180 <= 16'h975;
        src181 <= 16'h6175;
        src182 <= 16'h88fd;
        src183 <= 16'hb1a6;
        src184 <= 16'hdf3f;
        exp <= 24'h5c6ad8;
        #1
        src0 <= 16'hdc1d;
        src1 <= 16'h13ce;
        src2 <= 16'hf0f7;
        src3 <= 16'hf213;
        src4 <= 16'hd8bd;
        src5 <= 16'he1c5;
        src6 <= 16'h1782;
        src7 <= 16'he564;
        src8 <= 16'hbba8;
        src9 <= 16'hf567;
        src10 <= 16'h6862;
        src11 <= 16'h5755;
        src12 <= 16'ha3aa;
        src13 <= 16'h773a;
        src14 <= 16'h5a66;
        src15 <= 16'haf53;
        src16 <= 16'h8e22;
        src17 <= 16'he422;
        src18 <= 16'h6a46;
        src19 <= 16'he6ba;
        src20 <= 16'hbbc;
        src21 <= 16'hbe47;
        src22 <= 16'h100a;
        src23 <= 16'hd993;
        src24 <= 16'h8742;
        src25 <= 16'hd3cd;
        src26 <= 16'h26e5;
        src27 <= 16'hc97b;
        src28 <= 16'h4e5f;
        src29 <= 16'h322d;
        src30 <= 16'h2e56;
        src31 <= 16'h9090;
        src32 <= 16'h2585;
        src33 <= 16'h3db6;
        src34 <= 16'h4145;
        src35 <= 16'h3fc7;
        src36 <= 16'h5713;
        src37 <= 16'h3bbf;
        src38 <= 16'h9e74;
        src39 <= 16'hde8b;
        src40 <= 16'h6b51;
        src41 <= 16'h9118;
        src42 <= 16'h219d;
        src43 <= 16'he448;
        src44 <= 16'hbd35;
        src45 <= 16'h8ff6;
        src46 <= 16'ha8f7;
        src47 <= 16'h4c0f;
        src48 <= 16'heb56;
        src49 <= 16'h66b7;
        src50 <= 16'h3915;
        src51 <= 16'ha9ff;
        src52 <= 16'hd658;
        src53 <= 16'h78c1;
        src54 <= 16'hdf4d;
        src55 <= 16'h5633;
        src56 <= 16'h4b49;
        src57 <= 16'h114e;
        src58 <= 16'h83dd;
        src59 <= 16'h764f;
        src60 <= 16'hd1d5;
        src61 <= 16'hcdd2;
        src62 <= 16'h4ebe;
        src63 <= 16'h91a0;
        src64 <= 16'h13c0;
        src65 <= 16'h862;
        src66 <= 16'hbff4;
        src67 <= 16'h1203;
        src68 <= 16'h93ab;
        src69 <= 16'h4670;
        src70 <= 16'h9137;
        src71 <= 16'h30e4;
        src72 <= 16'h642e;
        src73 <= 16'he32b;
        src74 <= 16'h7b8e;
        src75 <= 16'h6424;
        src76 <= 16'h2eee;
        src77 <= 16'h5cd3;
        src78 <= 16'hb54b;
        src79 <= 16'hc121;
        src80 <= 16'h6a64;
        src81 <= 16'h1aac;
        src82 <= 16'hd251;
        src83 <= 16'h260a;
        src84 <= 16'h5e7f;
        src85 <= 16'h5b2c;
        src86 <= 16'ha804;
        src87 <= 16'h2ed;
        src88 <= 16'hb199;
        src89 <= 16'hf736;
        src90 <= 16'h91c7;
        src91 <= 16'h8b96;
        src92 <= 16'h6fe6;
        src93 <= 16'he300;
        src94 <= 16'h227c;
        src95 <= 16'h41bc;
        src96 <= 16'h8706;
        src97 <= 16'hf901;
        src98 <= 16'h9487;
        src99 <= 16'h244c;
        src100 <= 16'h2ecc;
        src101 <= 16'h342a;
        src102 <= 16'h98ee;
        src103 <= 16'ha37f;
        src104 <= 16'h3890;
        src105 <= 16'h8f33;
        src106 <= 16'h8ad4;
        src107 <= 16'h8486;
        src108 <= 16'hcc7f;
        src109 <= 16'h7f47;
        src110 <= 16'h6a41;
        src111 <= 16'h6eba;
        src112 <= 16'hfc97;
        src113 <= 16'hae8e;
        src114 <= 16'h28b2;
        src115 <= 16'h2c5f;
        src116 <= 16'h8207;
        src117 <= 16'h6277;
        src118 <= 16'h4b12;
        src119 <= 16'hba0a;
        src120 <= 16'h3412;
        src121 <= 16'haa39;
        src122 <= 16'h8464;
        src123 <= 16'h701;
        src124 <= 16'h5eac;
        src125 <= 16'hdba4;
        src126 <= 16'h4681;
        src127 <= 16'h9858;
        src128 <= 16'h4417;
        src129 <= 16'h4ddf;
        src130 <= 16'h9349;
        src131 <= 16'h79a7;
        src132 <= 16'h34db;
        src133 <= 16'ha18c;
        src134 <= 16'he1;
        src135 <= 16'h7b7f;
        src136 <= 16'h49b2;
        src137 <= 16'h9df8;
        src138 <= 16'h943d;
        src139 <= 16'hc12a;
        src140 <= 16'hef44;
        src141 <= 16'h9d59;
        src142 <= 16'hfc55;
        src143 <= 16'h3b31;
        src144 <= 16'h301b;
        src145 <= 16'hba3c;
        src146 <= 16'hb620;
        src147 <= 16'hd8c5;
        src148 <= 16'hf853;
        src149 <= 16'h6d02;
        src150 <= 16'hb55;
        src151 <= 16'hcd5f;
        src152 <= 16'hd2c1;
        src153 <= 16'h291d;
        src154 <= 16'h6ea4;
        src155 <= 16'hea97;
        src156 <= 16'h57ca;
        src157 <= 16'hbe81;
        src158 <= 16'h6e75;
        src159 <= 16'h5b6c;
        src160 <= 16'heeea;
        src161 <= 16'ha56;
        src162 <= 16'hfe0f;
        src163 <= 16'h94aa;
        src164 <= 16'h6665;
        src165 <= 16'h16d8;
        src166 <= 16'hc736;
        src167 <= 16'h4595;
        src168 <= 16'hbd2e;
        src169 <= 16'h1738;
        src170 <= 16'h2b8a;
        src171 <= 16'h20f4;
        src172 <= 16'hd939;
        src173 <= 16'h174a;
        src174 <= 16'h8fbc;
        src175 <= 16'h9daf;
        src176 <= 16'h942d;
        src177 <= 16'h13b7;
        src178 <= 16'hd081;
        src179 <= 16'h3c3c;
        src180 <= 16'h31b3;
        src181 <= 16'hba50;
        src182 <= 16'h3b45;
        src183 <= 16'h6b1e;
        src184 <= 16'h5ed;
        exp <= 24'h5abf6c;
        #1
        src0 <= 16'h5868;
        src1 <= 16'h4b4;
        src2 <= 16'h5529;
        src3 <= 16'h9993;
        src4 <= 16'h4a2f;
        src5 <= 16'h5245;
        src6 <= 16'hedf8;
        src7 <= 16'h3dab;
        src8 <= 16'h991a;
        src9 <= 16'h1fd;
        src10 <= 16'h3220;
        src11 <= 16'h1c07;
        src12 <= 16'hab01;
        src13 <= 16'hd64f;
        src14 <= 16'hbc50;
        src15 <= 16'hf241;
        src16 <= 16'h664;
        src17 <= 16'h12d;
        src18 <= 16'hc437;
        src19 <= 16'h940d;
        src20 <= 16'hefcd;
        src21 <= 16'hbc6e;
        src22 <= 16'h8ece;
        src23 <= 16'he75e;
        src24 <= 16'h7685;
        src25 <= 16'h94b;
        src26 <= 16'hff74;
        src27 <= 16'h84b1;
        src28 <= 16'hfa3e;
        src29 <= 16'h6fb1;
        src30 <= 16'h6daf;
        src31 <= 16'ha4e5;
        src32 <= 16'hcee8;
        src33 <= 16'h8b35;
        src34 <= 16'h166d;
        src35 <= 16'h3af;
        src36 <= 16'hf191;
        src37 <= 16'h73ba;
        src38 <= 16'h803d;
        src39 <= 16'h631d;
        src40 <= 16'h259d;
        src41 <= 16'he7f1;
        src42 <= 16'hfb8f;
        src43 <= 16'he2a2;
        src44 <= 16'h1678;
        src45 <= 16'hc0fb;
        src46 <= 16'h8d45;
        src47 <= 16'hd8cd;
        src48 <= 16'hd169;
        src49 <= 16'h6a45;
        src50 <= 16'hf297;
        src51 <= 16'ha900;
        src52 <= 16'h3951;
        src53 <= 16'h1ca2;
        src54 <= 16'h6bd5;
        src55 <= 16'hcf2f;
        src56 <= 16'h7063;
        src57 <= 16'he58f;
        src58 <= 16'h390c;
        src59 <= 16'h94ee;
        src60 <= 16'h372b;
        src61 <= 16'h2ff3;
        src62 <= 16'h773;
        src63 <= 16'hdd58;
        src64 <= 16'h5a07;
        src65 <= 16'h8514;
        src66 <= 16'hd24c;
        src67 <= 16'hea73;
        src68 <= 16'h8b43;
        src69 <= 16'h6a0d;
        src70 <= 16'h8111;
        src71 <= 16'h318b;
        src72 <= 16'h3315;
        src73 <= 16'h8ffc;
        src74 <= 16'h34a1;
        src75 <= 16'h4e01;
        src76 <= 16'h1a62;
        src77 <= 16'hfba9;
        src78 <= 16'h98b0;
        src79 <= 16'hd402;
        src80 <= 16'hf01;
        src81 <= 16'h4e0e;
        src82 <= 16'h3246;
        src83 <= 16'h6ea8;
        src84 <= 16'hcdaf;
        src85 <= 16'hce06;
        src86 <= 16'ha8da;
        src87 <= 16'h70bb;
        src88 <= 16'hb0ed;
        src89 <= 16'h3064;
        src90 <= 16'h8024;
        src91 <= 16'hf280;
        src92 <= 16'h60c;
        src93 <= 16'hc0dc;
        src94 <= 16'hab66;
        src95 <= 16'hb26d;
        src96 <= 16'h8531;
        src97 <= 16'hb50f;
        src98 <= 16'h76ca;
        src99 <= 16'h34bf;
        src100 <= 16'hb1e;
        src101 <= 16'h73a8;
        src102 <= 16'h398b;
        src103 <= 16'h6edc;
        src104 <= 16'h9a09;
        src105 <= 16'h7572;
        src106 <= 16'h1973;
        src107 <= 16'h705f;
        src108 <= 16'h2395;
        src109 <= 16'haa5a;
        src110 <= 16'h260f;
        src111 <= 16'h7478;
        src112 <= 16'h62a;
        src113 <= 16'haba5;
        src114 <= 16'hbec;
        src115 <= 16'h38c6;
        src116 <= 16'hdcd1;
        src117 <= 16'h7fe0;
        src118 <= 16'h5efb;
        src119 <= 16'ha71;
        src120 <= 16'h612d;
        src121 <= 16'h440d;
        src122 <= 16'h66b7;
        src123 <= 16'hcf5;
        src124 <= 16'hdb9f;
        src125 <= 16'ha62d;
        src126 <= 16'h3c01;
        src127 <= 16'h6ca1;
        src128 <= 16'hf8f3;
        src129 <= 16'ha87b;
        src130 <= 16'hdf9;
        src131 <= 16'h1e73;
        src132 <= 16'hd29;
        src133 <= 16'h3d14;
        src134 <= 16'h2b2d;
        src135 <= 16'had28;
        src136 <= 16'h926f;
        src137 <= 16'h79e9;
        src138 <= 16'hce45;
        src139 <= 16'h2cda;
        src140 <= 16'hc4e;
        src141 <= 16'h249c;
        src142 <= 16'h961;
        src143 <= 16'h15ab;
        src144 <= 16'h748e;
        src145 <= 16'hd9d6;
        src146 <= 16'ha52c;
        src147 <= 16'h66ac;
        src148 <= 16'ha809;
        src149 <= 16'h93ab;
        src150 <= 16'ha094;
        src151 <= 16'h2598;
        src152 <= 16'h35c9;
        src153 <= 16'hebf;
        src154 <= 16'he45b;
        src155 <= 16'h4d53;
        src156 <= 16'h5748;
        src157 <= 16'h3cbd;
        src158 <= 16'hf028;
        src159 <= 16'hb6e8;
        src160 <= 16'hd9b4;
        src161 <= 16'hc8cd;
        src162 <= 16'hd102;
        src163 <= 16'hf3ef;
        src164 <= 16'hf99f;
        src165 <= 16'hec86;
        src166 <= 16'hb4b9;
        src167 <= 16'h51eb;
        src168 <= 16'ha799;
        src169 <= 16'h1986;
        src170 <= 16'h350c;
        src171 <= 16'h7b79;
        src172 <= 16'hcdcd;
        src173 <= 16'h336a;
        src174 <= 16'ha515;
        src175 <= 16'h971;
        src176 <= 16'h7d44;
        src177 <= 16'h352;
        src178 <= 16'hc065;
        src179 <= 16'hebd7;
        src180 <= 16'hb6e;
        src181 <= 16'h4b9c;
        src182 <= 16'he6bc;
        src183 <= 16'hae5b;
        src184 <= 16'h9205;
        exp <= 24'h58aaa1;
        #1
        src0 <= 16'hd48c;
        src1 <= 16'hf922;
        src2 <= 16'h1019;
        src3 <= 16'h7529;
        src4 <= 16'hfc42;
        src5 <= 16'h3da9;
        src6 <= 16'ha8ed;
        src7 <= 16'h3fa0;
        src8 <= 16'hdcd2;
        src9 <= 16'hb38a;
        src10 <= 16'hf7f8;
        src11 <= 16'hca6;
        src12 <= 16'h8fcc;
        src13 <= 16'h3d6a;
        src14 <= 16'hdb8;
        src15 <= 16'hbccb;
        src16 <= 16'h4719;
        src17 <= 16'hb38c;
        src18 <= 16'hf6c2;
        src19 <= 16'h8708;
        src20 <= 16'h8692;
        src21 <= 16'h6ae2;
        src22 <= 16'h973f;
        src23 <= 16'h50f7;
        src24 <= 16'hc56a;
        src25 <= 16'h32fb;
        src26 <= 16'h88f2;
        src27 <= 16'he85a;
        src28 <= 16'hb252;
        src29 <= 16'hdbf9;
        src30 <= 16'h2def;
        src31 <= 16'hb491;
        src32 <= 16'h14a1;
        src33 <= 16'h866c;
        src34 <= 16'hb90a;
        src35 <= 16'hf926;
        src36 <= 16'hfd97;
        src37 <= 16'hdd18;
        src38 <= 16'h4dbb;
        src39 <= 16'hf4e0;
        src40 <= 16'heed4;
        src41 <= 16'h512a;
        src42 <= 16'h6e95;
        src43 <= 16'hb8bf;
        src44 <= 16'h59e;
        src45 <= 16'ha592;
        src46 <= 16'h9991;
        src47 <= 16'h9ea9;
        src48 <= 16'h6f99;
        src49 <= 16'h72ea;
        src50 <= 16'he095;
        src51 <= 16'hc400;
        src52 <= 16'hfb92;
        src53 <= 16'he136;
        src54 <= 16'h4147;
        src55 <= 16'hb1a2;
        src56 <= 16'he2d7;
        src57 <= 16'hd6a2;
        src58 <= 16'h3dfb;
        src59 <= 16'h502a;
        src60 <= 16'h4098;
        src61 <= 16'h85f5;
        src62 <= 16'h801a;
        src63 <= 16'h4831;
        src64 <= 16'h352b;
        src65 <= 16'h7f4f;
        src66 <= 16'ha2f;
        src67 <= 16'h46d8;
        src68 <= 16'h7cc9;
        src69 <= 16'hfc73;
        src70 <= 16'h1be3;
        src71 <= 16'h10b6;
        src72 <= 16'he795;
        src73 <= 16'h2e39;
        src74 <= 16'hfacc;
        src75 <= 16'he5b9;
        src76 <= 16'h241e;
        src77 <= 16'h728d;
        src78 <= 16'hb33b;
        src79 <= 16'h4c25;
        src80 <= 16'hf4fa;
        src81 <= 16'h502d;
        src82 <= 16'h76d2;
        src83 <= 16'ha14a;
        src84 <= 16'h6909;
        src85 <= 16'h38cc;
        src86 <= 16'h67b9;
        src87 <= 16'h3907;
        src88 <= 16'h628b;
        src89 <= 16'h577;
        src90 <= 16'h5322;
        src91 <= 16'h2c4d;
        src92 <= 16'h124e;
        src93 <= 16'h5f6e;
        src94 <= 16'hd48b;
        src95 <= 16'h83fb;
        src96 <= 16'h9050;
        src97 <= 16'hb36f;
        src98 <= 16'h2356;
        src99 <= 16'hb17a;
        src100 <= 16'hea97;
        src101 <= 16'h2c59;
        src102 <= 16'h6d89;
        src103 <= 16'hfba1;
        src104 <= 16'hb9ee;
        src105 <= 16'h7ec1;
        src106 <= 16'hf176;
        src107 <= 16'ha442;
        src108 <= 16'h7213;
        src109 <= 16'hb3c8;
        src110 <= 16'hd3d2;
        src111 <= 16'hd8dd;
        src112 <= 16'h3961;
        src113 <= 16'hf35d;
        src114 <= 16'hf4ab;
        src115 <= 16'hb825;
        src116 <= 16'hcc46;
        src117 <= 16'ha60c;
        src118 <= 16'hf161;
        src119 <= 16'h9bd4;
        src120 <= 16'hdc4f;
        src121 <= 16'h548c;
        src122 <= 16'h10ea;
        src123 <= 16'h1ff0;
        src124 <= 16'h9640;
        src125 <= 16'hbe5f;
        src126 <= 16'h4f5a;
        src127 <= 16'h6ff0;
        src128 <= 16'h62ac;
        src129 <= 16'hc002;
        src130 <= 16'h2f23;
        src131 <= 16'h1a15;
        src132 <= 16'h2f7f;
        src133 <= 16'h919b;
        src134 <= 16'h300;
        src135 <= 16'h9662;
        src136 <= 16'hef46;
        src137 <= 16'hb2c4;
        src138 <= 16'h9d3b;
        src139 <= 16'hf4d;
        src140 <= 16'h4e6e;
        src141 <= 16'h79d5;
        src142 <= 16'hf215;
        src143 <= 16'hce4c;
        src144 <= 16'hf791;
        src145 <= 16'h4393;
        src146 <= 16'he511;
        src147 <= 16'h631d;
        src148 <= 16'h6462;
        src149 <= 16'ha16f;
        src150 <= 16'hd56e;
        src151 <= 16'h516e;
        src152 <= 16'h9963;
        src153 <= 16'h8ab;
        src154 <= 16'hea52;
        src155 <= 16'h314f;
        src156 <= 16'hb983;
        src157 <= 16'h1c03;
        src158 <= 16'h7a9f;
        src159 <= 16'h56b4;
        src160 <= 16'h7ae1;
        src161 <= 16'h780;
        src162 <= 16'h922c;
        src163 <= 16'hd70b;
        src164 <= 16'h7f0c;
        src165 <= 16'h3877;
        src166 <= 16'h99b7;
        src167 <= 16'hda96;
        src168 <= 16'h49d2;
        src169 <= 16'hf438;
        src170 <= 16'hf96;
        src171 <= 16'h17de;
        src172 <= 16'hf2e9;
        src173 <= 16'h5973;
        src174 <= 16'hfa34;
        src175 <= 16'h10d6;
        src176 <= 16'h3880;
        src177 <= 16'h69c9;
        src178 <= 16'h4b5b;
        src179 <= 16'hc0df;
        src180 <= 16'hc7ec;
        src181 <= 16'h9f0;
        src182 <= 16'h2d94;
        src183 <= 16'hbaeb;
        src184 <= 16'he07a;
        exp <= 24'h619281;
        #1
        src0 <= 16'h2c8c;
        src1 <= 16'h4730;
        src2 <= 16'ha96e;
        src3 <= 16'h5da2;
        src4 <= 16'hedde;
        src5 <= 16'hf6b3;
        src6 <= 16'h86ea;
        src7 <= 16'h883c;
        src8 <= 16'hb54a;
        src9 <= 16'h8708;
        src10 <= 16'hd9d3;
        src11 <= 16'h8d23;
        src12 <= 16'h2b78;
        src13 <= 16'h8ffa;
        src14 <= 16'h990b;
        src15 <= 16'h109a;
        src16 <= 16'h5fe4;
        src17 <= 16'h793d;
        src18 <= 16'hc2f1;
        src19 <= 16'hba0f;
        src20 <= 16'hecb5;
        src21 <= 16'hc4ca;
        src22 <= 16'hc11f;
        src23 <= 16'h36e2;
        src24 <= 16'h9d11;
        src25 <= 16'h1e42;
        src26 <= 16'h11ca;
        src27 <= 16'h235d;
        src28 <= 16'h9a63;
        src29 <= 16'hb799;
        src30 <= 16'hfab5;
        src31 <= 16'h3722;
        src32 <= 16'h77ea;
        src33 <= 16'h4408;
        src34 <= 16'h4e0d;
        src35 <= 16'h508c;
        src36 <= 16'h9bf0;
        src37 <= 16'hd595;
        src38 <= 16'h39bc;
        src39 <= 16'heaed;
        src40 <= 16'h4fc;
        src41 <= 16'h8f51;
        src42 <= 16'hb2e3;
        src43 <= 16'h7a49;
        src44 <= 16'hbdcd;
        src45 <= 16'h90c0;
        src46 <= 16'h4564;
        src47 <= 16'h27c1;
        src48 <= 16'hfa64;
        src49 <= 16'h31fc;
        src50 <= 16'h21d2;
        src51 <= 16'h3d6d;
        src52 <= 16'h74dd;
        src53 <= 16'hda1e;
        src54 <= 16'h17c7;
        src55 <= 16'h1e2b;
        src56 <= 16'h52a5;
        src57 <= 16'h94a5;
        src58 <= 16'h5fea;
        src59 <= 16'h191e;
        src60 <= 16'h636e;
        src61 <= 16'he574;
        src62 <= 16'h8659;
        src63 <= 16'h1e6e;
        src64 <= 16'hebad;
        src65 <= 16'h6451;
        src66 <= 16'h11ba;
        src67 <= 16'he182;
        src68 <= 16'ha39;
        src69 <= 16'h53bb;
        src70 <= 16'hb583;
        src71 <= 16'he765;
        src72 <= 16'habdd;
        src73 <= 16'h7b15;
        src74 <= 16'he662;
        src75 <= 16'hd7e2;
        src76 <= 16'h4f92;
        src77 <= 16'h232c;
        src78 <= 16'hebd0;
        src79 <= 16'hd63e;
        src80 <= 16'h9812;
        src81 <= 16'h4cdd;
        src82 <= 16'hba01;
        src83 <= 16'h41db;
        src84 <= 16'hd315;
        src85 <= 16'h5f8e;
        src86 <= 16'h9c8a;
        src87 <= 16'hde28;
        src88 <= 16'h6269;
        src89 <= 16'hb3a;
        src90 <= 16'h67af;
        src91 <= 16'h9df5;
        src92 <= 16'hf025;
        src93 <= 16'hd27f;
        src94 <= 16'h6879;
        src95 <= 16'h1f22;
        src96 <= 16'h646;
        src97 <= 16'h1f20;
        src98 <= 16'hca2b;
        src99 <= 16'h500c;
        src100 <= 16'h1be6;
        src101 <= 16'hef3d;
        src102 <= 16'h96cf;
        src103 <= 16'h5498;
        src104 <= 16'hff6d;
        src105 <= 16'h885b;
        src106 <= 16'hce50;
        src107 <= 16'hd391;
        src108 <= 16'h7f;
        src109 <= 16'h9cc9;
        src110 <= 16'he70e;
        src111 <= 16'h837a;
        src112 <= 16'hfeb2;
        src113 <= 16'h1f04;
        src114 <= 16'hd76;
        src115 <= 16'h9eeb;
        src116 <= 16'h1a0e;
        src117 <= 16'ha9f3;
        src118 <= 16'h3564;
        src119 <= 16'he421;
        src120 <= 16'hd29c;
        src121 <= 16'hf326;
        src122 <= 16'hccfc;
        src123 <= 16'hd53c;
        src124 <= 16'hce80;
        src125 <= 16'hbaaa;
        src126 <= 16'h762;
        src127 <= 16'h74b5;
        src128 <= 16'h3e29;
        src129 <= 16'hca10;
        src130 <= 16'h8d97;
        src131 <= 16'hc189;
        src132 <= 16'h4403;
        src133 <= 16'h8634;
        src134 <= 16'hae8;
        src135 <= 16'h96e5;
        src136 <= 16'h556d;
        src137 <= 16'h4648;
        src138 <= 16'hb3bf;
        src139 <= 16'hb64;
        src140 <= 16'hbfc0;
        src141 <= 16'h53b7;
        src142 <= 16'h9254;
        src143 <= 16'h928a;
        src144 <= 16'h36d6;
        src145 <= 16'h2ebf;
        src146 <= 16'h3d8a;
        src147 <= 16'he71b;
        src148 <= 16'h5d6b;
        src149 <= 16'h3578;
        src150 <= 16'h9702;
        src151 <= 16'hcb26;
        src152 <= 16'h98c0;
        src153 <= 16'he335;
        src154 <= 16'haa12;
        src155 <= 16'h2700;
        src156 <= 16'h2683;
        src157 <= 16'h69f2;
        src158 <= 16'h6c98;
        src159 <= 16'he850;
        src160 <= 16'hcad0;
        src161 <= 16'he33e;
        src162 <= 16'h7e6;
        src163 <= 16'hbc2c;
        src164 <= 16'hc5c5;
        src165 <= 16'h92d5;
        src166 <= 16'h4886;
        src167 <= 16'h75a8;
        src168 <= 16'hbf95;
        src169 <= 16'h8187;
        src170 <= 16'h339;
        src171 <= 16'h821a;
        src172 <= 16'he8a9;
        src173 <= 16'hb59f;
        src174 <= 16'h9c69;
        src175 <= 16'h41e1;
        src176 <= 16'h84a;
        src177 <= 16'h29b0;
        src178 <= 16'hb991;
        src179 <= 16'h2eb3;
        src180 <= 16'heafc;
        src181 <= 16'h45b9;
        src182 <= 16'h27cc;
        src183 <= 16'h24d1;
        src184 <= 16'h9138;
        exp <= 24'h5cd455;
        #1
        src0 <= 16'hef2f;
        src1 <= 16'ha92f;
        src2 <= 16'hdc3b;
        src3 <= 16'hc774;
        src4 <= 16'h48ad;
        src5 <= 16'h17ad;
        src6 <= 16'hb5b8;
        src7 <= 16'h862e;
        src8 <= 16'h463d;
        src9 <= 16'h9e83;
        src10 <= 16'h76f6;
        src11 <= 16'hd63;
        src12 <= 16'h6957;
        src13 <= 16'hf59a;
        src14 <= 16'h5adb;
        src15 <= 16'hb8c9;
        src16 <= 16'h4b87;
        src17 <= 16'hbd1c;
        src18 <= 16'h30db;
        src19 <= 16'hbb79;
        src20 <= 16'hac9f;
        src21 <= 16'hf07e;
        src22 <= 16'h4ef5;
        src23 <= 16'h1cac;
        src24 <= 16'h7f9f;
        src25 <= 16'h17d7;
        src26 <= 16'h5e97;
        src27 <= 16'hd458;
        src28 <= 16'h720b;
        src29 <= 16'h7b3a;
        src30 <= 16'h1021;
        src31 <= 16'h375e;
        src32 <= 16'hda19;
        src33 <= 16'h34e8;
        src34 <= 16'hed7f;
        src35 <= 16'h5eee;
        src36 <= 16'ha75e;
        src37 <= 16'h3039;
        src38 <= 16'hd4b6;
        src39 <= 16'hed2b;
        src40 <= 16'h24d3;
        src41 <= 16'h9071;
        src42 <= 16'hb050;
        src43 <= 16'hd73b;
        src44 <= 16'hd236;
        src45 <= 16'h8f22;
        src46 <= 16'hd0c;
        src47 <= 16'h56f7;
        src48 <= 16'h8e85;
        src49 <= 16'h1292;
        src50 <= 16'he9e6;
        src51 <= 16'heb4e;
        src52 <= 16'h3908;
        src53 <= 16'h3e3d;
        src54 <= 16'hbe5;
        src55 <= 16'he1d;
        src56 <= 16'haf6a;
        src57 <= 16'h520c;
        src58 <= 16'h761f;
        src59 <= 16'he9b8;
        src60 <= 16'hd9c0;
        src61 <= 16'h2472;
        src62 <= 16'h575d;
        src63 <= 16'hb3f7;
        src64 <= 16'heaf6;
        src65 <= 16'h9c1;
        src66 <= 16'h25d5;
        src67 <= 16'h59a6;
        src68 <= 16'h8f24;
        src69 <= 16'hd4cd;
        src70 <= 16'h3da5;
        src71 <= 16'ha560;
        src72 <= 16'h4a4b;
        src73 <= 16'h5d9d;
        src74 <= 16'h1350;
        src75 <= 16'hb0e3;
        src76 <= 16'h1856;
        src77 <= 16'h8e94;
        src78 <= 16'h51b9;
        src79 <= 16'h22fa;
        src80 <= 16'h3dc8;
        src81 <= 16'h6dd8;
        src82 <= 16'hd9ac;
        src83 <= 16'he75;
        src84 <= 16'h45f2;
        src85 <= 16'hc20d;
        src86 <= 16'he896;
        src87 <= 16'h5937;
        src88 <= 16'h5662;
        src89 <= 16'hc692;
        src90 <= 16'h953e;
        src91 <= 16'hf1eb;
        src92 <= 16'hd780;
        src93 <= 16'h49bc;
        src94 <= 16'hd485;
        src95 <= 16'hb9e9;
        src96 <= 16'hbd3e;
        src97 <= 16'h99c0;
        src98 <= 16'h52a2;
        src99 <= 16'h91ed;
        src100 <= 16'h2939;
        src101 <= 16'h9115;
        src102 <= 16'hf42b;
        src103 <= 16'h5751;
        src104 <= 16'h7fbe;
        src105 <= 16'h6d83;
        src106 <= 16'h3829;
        src107 <= 16'h3b88;
        src108 <= 16'h43f7;
        src109 <= 16'h6083;
        src110 <= 16'h27e;
        src111 <= 16'he0dc;
        src112 <= 16'ha38b;
        src113 <= 16'hb9b2;
        src114 <= 16'h6e0e;
        src115 <= 16'hf092;
        src116 <= 16'h75e4;
        src117 <= 16'h3cf6;
        src118 <= 16'ha447;
        src119 <= 16'hf674;
        src120 <= 16'h5d48;
        src121 <= 16'h8d0a;
        src122 <= 16'h14f0;
        src123 <= 16'h1794;
        src124 <= 16'h35b;
        src125 <= 16'h826a;
        src126 <= 16'h91e2;
        src127 <= 16'h94e6;
        src128 <= 16'h42e0;
        src129 <= 16'had72;
        src130 <= 16'h8efa;
        src131 <= 16'hada2;
        src132 <= 16'h1f0e;
        src133 <= 16'he294;
        src134 <= 16'hd380;
        src135 <= 16'h5b35;
        src136 <= 16'hd611;
        src137 <= 16'h63fb;
        src138 <= 16'h35ee;
        src139 <= 16'hf671;
        src140 <= 16'hd72;
        src141 <= 16'h5be6;
        src142 <= 16'h2165;
        src143 <= 16'h70e6;
        src144 <= 16'hca04;
        src145 <= 16'haece;
        src146 <= 16'h2377;
        src147 <= 16'hc5cc;
        src148 <= 16'h7e0a;
        src149 <= 16'ha1e4;
        src150 <= 16'he162;
        src151 <= 16'hdf78;
        src152 <= 16'h55f;
        src153 <= 16'h6014;
        src154 <= 16'h2d69;
        src155 <= 16'h2723;
        src156 <= 16'h26bd;
        src157 <= 16'h450a;
        src158 <= 16'hca33;
        src159 <= 16'h9d5c;
        src160 <= 16'hdeae;
        src161 <= 16'h306e;
        src162 <= 16'h8ac2;
        src163 <= 16'h772a;
        src164 <= 16'h3699;
        src165 <= 16'h9bed;
        src166 <= 16'hcf8a;
        src167 <= 16'h7914;
        src168 <= 16'h9383;
        src169 <= 16'hb218;
        src170 <= 16'h900b;
        src171 <= 16'h1035;
        src172 <= 16'h4598;
        src173 <= 16'h8e1b;
        src174 <= 16'h154;
        src175 <= 16'hfa2a;
        src176 <= 16'h1c16;
        src177 <= 16'hf600;
        src178 <= 16'hd576;
        src179 <= 16'hf058;
        src180 <= 16'h930b;
        src181 <= 16'hc761;
        src182 <= 16'he71d;
        src183 <= 16'h9624;
        src184 <= 16'he5b0;
        exp <= 24'h5c8b72;
        #1
        src0 <= 16'hdc7b;
        src1 <= 16'h363b;
        src2 <= 16'h474b;
        src3 <= 16'hd1b2;
        src4 <= 16'hac10;
        src5 <= 16'h4af5;
        src6 <= 16'hc9b3;
        src7 <= 16'h7ea0;
        src8 <= 16'hbb5b;
        src9 <= 16'h1346;
        src10 <= 16'h33de;
        src11 <= 16'hd4f2;
        src12 <= 16'h65f6;
        src13 <= 16'hfe91;
        src14 <= 16'h53e0;
        src15 <= 16'h582e;
        src16 <= 16'h54b0;
        src17 <= 16'hfba9;
        src18 <= 16'hbf22;
        src19 <= 16'hd11a;
        src20 <= 16'h8643;
        src21 <= 16'h267c;
        src22 <= 16'h9b85;
        src23 <= 16'hab34;
        src24 <= 16'hab80;
        src25 <= 16'hc883;
        src26 <= 16'h4cf;
        src27 <= 16'h816e;
        src28 <= 16'h7919;
        src29 <= 16'h790e;
        src30 <= 16'hb2e4;
        src31 <= 16'hc730;
        src32 <= 16'h39ca;
        src33 <= 16'h7360;
        src34 <= 16'hd9ea;
        src35 <= 16'h20;
        src36 <= 16'hcbf3;
        src37 <= 16'h7437;
        src38 <= 16'hc12d;
        src39 <= 16'h3b5e;
        src40 <= 16'hdf40;
        src41 <= 16'h91c;
        src42 <= 16'hbda8;
        src43 <= 16'h40cf;
        src44 <= 16'h3526;
        src45 <= 16'h5bd2;
        src46 <= 16'hf7a2;
        src47 <= 16'hf13a;
        src48 <= 16'h57f9;
        src49 <= 16'h1d49;
        src50 <= 16'h5f69;
        src51 <= 16'h715d;
        src52 <= 16'h2563;
        src53 <= 16'h4212;
        src54 <= 16'hde35;
        src55 <= 16'h24a1;
        src56 <= 16'hae23;
        src57 <= 16'he491;
        src58 <= 16'hed99;
        src59 <= 16'hac25;
        src60 <= 16'hc67f;
        src61 <= 16'h403d;
        src62 <= 16'he06c;
        src63 <= 16'hf5ee;
        src64 <= 16'ha27;
        src65 <= 16'hf66f;
        src66 <= 16'h1cdb;
        src67 <= 16'h50e7;
        src68 <= 16'h86c;
        src69 <= 16'h5f03;
        src70 <= 16'h94f0;
        src71 <= 16'h54a5;
        src72 <= 16'hd2c7;
        src73 <= 16'hbb0f;
        src74 <= 16'h6fd7;
        src75 <= 16'h9d4a;
        src76 <= 16'h56bf;
        src77 <= 16'h80c9;
        src78 <= 16'h19bc;
        src79 <= 16'hefb5;
        src80 <= 16'h669c;
        src81 <= 16'h2615;
        src82 <= 16'hc50;
        src83 <= 16'hd64d;
        src84 <= 16'h547e;
        src85 <= 16'h1c7b;
        src86 <= 16'h1a31;
        src87 <= 16'h5179;
        src88 <= 16'h7a6f;
        src89 <= 16'ha389;
        src90 <= 16'h6f5d;
        src91 <= 16'hadd7;
        src92 <= 16'hec3d;
        src93 <= 16'h8e31;
        src94 <= 16'h523c;
        src95 <= 16'h5a1c;
        src96 <= 16'h4dfa;
        src97 <= 16'hf286;
        src98 <= 16'h37a9;
        src99 <= 16'hcc38;
        src100 <= 16'heea7;
        src101 <= 16'h8642;
        src102 <= 16'h8221;
        src103 <= 16'h4a76;
        src104 <= 16'h68f1;
        src105 <= 16'h1f37;
        src106 <= 16'h350;
        src107 <= 16'he9e9;
        src108 <= 16'h4091;
        src109 <= 16'h8b70;
        src110 <= 16'h786c;
        src111 <= 16'h5b65;
        src112 <= 16'h6512;
        src113 <= 16'h6365;
        src114 <= 16'h1231;
        src115 <= 16'hd74e;
        src116 <= 16'h87eb;
        src117 <= 16'he20b;
        src118 <= 16'h6734;
        src119 <= 16'h7550;
        src120 <= 16'hd421;
        src121 <= 16'h943e;
        src122 <= 16'h2f1b;
        src123 <= 16'hc3b;
        src124 <= 16'h8891;
        src125 <= 16'hb7d9;
        src126 <= 16'hde9c;
        src127 <= 16'h289a;
        src128 <= 16'hcced;
        src129 <= 16'hc9cd;
        src130 <= 16'hc996;
        src131 <= 16'habcf;
        src132 <= 16'ha60a;
        src133 <= 16'h6424;
        src134 <= 16'h40ed;
        src135 <= 16'hb6a4;
        src136 <= 16'h3e6c;
        src137 <= 16'h2ad3;
        src138 <= 16'h9c66;
        src139 <= 16'h6106;
        src140 <= 16'h4375;
        src141 <= 16'hb16b;
        src142 <= 16'h9440;
        src143 <= 16'hf82;
        src144 <= 16'h8d81;
        src145 <= 16'h382e;
        src146 <= 16'heea9;
        src147 <= 16'hff8e;
        src148 <= 16'hb26b;
        src149 <= 16'h4539;
        src150 <= 16'h4eff;
        src151 <= 16'h6207;
        src152 <= 16'h17;
        src153 <= 16'h6e53;
        src154 <= 16'hbd3d;
        src155 <= 16'h9a92;
        src156 <= 16'h1f28;
        src157 <= 16'h9b6;
        src158 <= 16'h25a8;
        src159 <= 16'ha5b8;
        src160 <= 16'hc867;
        src161 <= 16'h5c98;
        src162 <= 16'h8a0b;
        src163 <= 16'hf46c;
        src164 <= 16'h33f3;
        src165 <= 16'hcea7;
        src166 <= 16'h25f6;
        src167 <= 16'h988c;
        src168 <= 16'hb40c;
        src169 <= 16'h2c05;
        src170 <= 16'he989;
        src171 <= 16'h8c4a;
        src172 <= 16'h6f82;
        src173 <= 16'h9753;
        src174 <= 16'hc474;
        src175 <= 16'hf546;
        src176 <= 16'hbde0;
        src177 <= 16'h9483;
        src178 <= 16'h5f4e;
        src179 <= 16'h5705;
        src180 <= 16'h33b2;
        src181 <= 16'h82d8;
        src182 <= 16'hfe;
        src183 <= 16'hd851;
        src184 <= 16'heb64;
        exp <= 24'h5cf736;
        #1
        src0 <= 16'haf49;
        src1 <= 16'h1df;
        src2 <= 16'ha190;
        src3 <= 16'h7a90;
        src4 <= 16'hcc38;
        src5 <= 16'h98d6;
        src6 <= 16'ha981;
        src7 <= 16'hcf11;
        src8 <= 16'hced1;
        src9 <= 16'hb006;
        src10 <= 16'h7e70;
        src11 <= 16'hcb8;
        src12 <= 16'h5c42;
        src13 <= 16'h9df5;
        src14 <= 16'h932d;
        src15 <= 16'h6de3;
        src16 <= 16'hc54d;
        src17 <= 16'h8531;
        src18 <= 16'hf832;
        src19 <= 16'hbe71;
        src20 <= 16'h6cb8;
        src21 <= 16'hdfd6;
        src22 <= 16'h45cf;
        src23 <= 16'h23dd;
        src24 <= 16'h2d5;
        src25 <= 16'h8363;
        src26 <= 16'h1524;
        src27 <= 16'hf685;
        src28 <= 16'hdac;
        src29 <= 16'h8113;
        src30 <= 16'hdf2b;
        src31 <= 16'h17de;
        src32 <= 16'hd16f;
        src33 <= 16'hbe0c;
        src34 <= 16'hcc93;
        src35 <= 16'h8bd0;
        src36 <= 16'he954;
        src37 <= 16'h3caf;
        src38 <= 16'h2d57;
        src39 <= 16'h12be;
        src40 <= 16'h7f38;
        src41 <= 16'hddf9;
        src42 <= 16'h6a30;
        src43 <= 16'h1743;
        src44 <= 16'hbd3c;
        src45 <= 16'h20cc;
        src46 <= 16'hc0b4;
        src47 <= 16'hf459;
        src48 <= 16'h7ae6;
        src49 <= 16'h21c4;
        src50 <= 16'h714d;
        src51 <= 16'h75d5;
        src52 <= 16'h9d80;
        src53 <= 16'h3665;
        src54 <= 16'h51d0;
        src55 <= 16'hffc7;
        src56 <= 16'h50db;
        src57 <= 16'h7cf9;
        src58 <= 16'h347d;
        src59 <= 16'h3b5d;
        src60 <= 16'hd556;
        src61 <= 16'heb02;
        src62 <= 16'h1532;
        src63 <= 16'hea66;
        src64 <= 16'he466;
        src65 <= 16'he656;
        src66 <= 16'hb6b9;
        src67 <= 16'h2cf;
        src68 <= 16'h4c34;
        src69 <= 16'h10c2;
        src70 <= 16'hf500;
        src71 <= 16'he354;
        src72 <= 16'hf7fd;
        src73 <= 16'ha66d;
        src74 <= 16'h2d2c;
        src75 <= 16'hb2ba;
        src76 <= 16'hccdf;
        src77 <= 16'h3fc0;
        src78 <= 16'h8233;
        src79 <= 16'h3c6d;
        src80 <= 16'h3fc;
        src81 <= 16'h3a8b;
        src82 <= 16'hdf4e;
        src83 <= 16'hdb39;
        src84 <= 16'h3f7f;
        src85 <= 16'hc49d;
        src86 <= 16'hab96;
        src87 <= 16'hef2f;
        src88 <= 16'h5a3c;
        src89 <= 16'h6730;
        src90 <= 16'h4e8a;
        src91 <= 16'he8ef;
        src92 <= 16'h5d5;
        src93 <= 16'ha99b;
        src94 <= 16'h5a9b;
        src95 <= 16'h1e14;
        src96 <= 16'hb793;
        src97 <= 16'he7e5;
        src98 <= 16'h7a0;
        src99 <= 16'h735f;
        src100 <= 16'hd55d;
        src101 <= 16'h6671;
        src102 <= 16'hb301;
        src103 <= 16'h8774;
        src104 <= 16'h9935;
        src105 <= 16'h184;
        src106 <= 16'hc6a1;
        src107 <= 16'hf905;
        src108 <= 16'hbc4d;
        src109 <= 16'h9f28;
        src110 <= 16'hc60b;
        src111 <= 16'h43a6;
        src112 <= 16'he85f;
        src113 <= 16'hc054;
        src114 <= 16'h124a;
        src115 <= 16'h1c22;
        src116 <= 16'h521e;
        src117 <= 16'h4deb;
        src118 <= 16'h1f10;
        src119 <= 16'h1006;
        src120 <= 16'hd230;
        src121 <= 16'haacf;
        src122 <= 16'h9469;
        src123 <= 16'h622c;
        src124 <= 16'h8f1b;
        src125 <= 16'h9107;
        src126 <= 16'h4f39;
        src127 <= 16'h24a8;
        src128 <= 16'h5e76;
        src129 <= 16'h5f32;
        src130 <= 16'h13b9;
        src131 <= 16'ha0ac;
        src132 <= 16'hbcc7;
        src133 <= 16'ha61c;
        src134 <= 16'h1e84;
        src135 <= 16'heb5d;
        src136 <= 16'h6ea;
        src137 <= 16'hf8f8;
        src138 <= 16'h5862;
        src139 <= 16'hd6b;
        src140 <= 16'h7990;
        src141 <= 16'he826;
        src142 <= 16'h86db;
        src143 <= 16'h6176;
        src144 <= 16'h4f98;
        src145 <= 16'h620e;
        src146 <= 16'hbc5d;
        src147 <= 16'h66dc;
        src148 <= 16'h66d9;
        src149 <= 16'hd7;
        src150 <= 16'h89c5;
        src151 <= 16'hbdf1;
        src152 <= 16'hbc1b;
        src153 <= 16'he6f2;
        src154 <= 16'heb44;
        src155 <= 16'hcfe9;
        src156 <= 16'h940d;
        src157 <= 16'he25d;
        src158 <= 16'h4d00;
        src159 <= 16'h4304;
        src160 <= 16'hc015;
        src161 <= 16'he40d;
        src162 <= 16'h523;
        src163 <= 16'hc12a;
        src164 <= 16'h32a;
        src165 <= 16'h6df6;
        src166 <= 16'hb19;
        src167 <= 16'hee4f;
        src168 <= 16'h110f;
        src169 <= 16'h9de0;
        src170 <= 16'hfbf0;
        src171 <= 16'hf36;
        src172 <= 16'h9b05;
        src173 <= 16'hcba7;
        src174 <= 16'h76b5;
        src175 <= 16'h58df;
        src176 <= 16'hd977;
        src177 <= 16'he0b2;
        src178 <= 16'h265;
        src179 <= 16'he0b6;
        src180 <= 16'h79b9;
        src181 <= 16'hb699;
        src182 <= 16'hebb4;
        src183 <= 16'h2200;
        src184 <= 16'h11ca;
        exp <= 24'h5ec9bf;
        #1
        src0 <= 16'h140c;
        src1 <= 16'hd213;
        src2 <= 16'h9d60;
        src3 <= 16'h4fd1;
        src4 <= 16'h294b;
        src5 <= 16'h726c;
        src6 <= 16'h767e;
        src7 <= 16'hffbf;
        src8 <= 16'hd439;
        src9 <= 16'he67;
        src10 <= 16'ha767;
        src11 <= 16'h4dcb;
        src12 <= 16'hf8ea;
        src13 <= 16'h1fe8;
        src14 <= 16'h3e21;
        src15 <= 16'h9181;
        src16 <= 16'he6b8;
        src17 <= 16'h46c9;
        src18 <= 16'h729e;
        src19 <= 16'h95b6;
        src20 <= 16'ha7c2;
        src21 <= 16'h1c66;
        src22 <= 16'heb81;
        src23 <= 16'he9f4;
        src24 <= 16'h740e;
        src25 <= 16'hec9e;
        src26 <= 16'hbcbf;
        src27 <= 16'h237b;
        src28 <= 16'h7260;
        src29 <= 16'h6d85;
        src30 <= 16'he193;
        src31 <= 16'he11;
        src32 <= 16'h8825;
        src33 <= 16'haba6;
        src34 <= 16'h6649;
        src35 <= 16'h90e8;
        src36 <= 16'hbccf;
        src37 <= 16'hbc8;
        src38 <= 16'hcb0d;
        src39 <= 16'hb047;
        src40 <= 16'hbf48;
        src41 <= 16'h66bc;
        src42 <= 16'hed4c;
        src43 <= 16'hebd0;
        src44 <= 16'heb8f;
        src45 <= 16'h5a15;
        src46 <= 16'h1c8f;
        src47 <= 16'ha940;
        src48 <= 16'hf5da;
        src49 <= 16'ha2a2;
        src50 <= 16'h4362;
        src51 <= 16'had47;
        src52 <= 16'h1352;
        src53 <= 16'hf0dd;
        src54 <= 16'hd894;
        src55 <= 16'h210a;
        src56 <= 16'h5edc;
        src57 <= 16'h3879;
        src58 <= 16'h457;
        src59 <= 16'h2f7f;
        src60 <= 16'h1262;
        src61 <= 16'h5994;
        src62 <= 16'hc671;
        src63 <= 16'h539e;
        src64 <= 16'h3075;
        src65 <= 16'hba9c;
        src66 <= 16'hef8f;
        src67 <= 16'h536b;
        src68 <= 16'he8c5;
        src69 <= 16'h1396;
        src70 <= 16'h6f6a;
        src71 <= 16'hb087;
        src72 <= 16'hb157;
        src73 <= 16'h4be9;
        src74 <= 16'h3d3a;
        src75 <= 16'h35a3;
        src76 <= 16'hda57;
        src77 <= 16'h978d;
        src78 <= 16'h4aff;
        src79 <= 16'hb041;
        src80 <= 16'h5dea;
        src81 <= 16'hed2e;
        src82 <= 16'hcea6;
        src83 <= 16'h4528;
        src84 <= 16'hf404;
        src85 <= 16'h567a;
        src86 <= 16'hcf1e;
        src87 <= 16'h57ed;
        src88 <= 16'hc2d;
        src89 <= 16'hba7;
        src90 <= 16'h8940;
        src91 <= 16'h8be8;
        src92 <= 16'hf193;
        src93 <= 16'h3074;
        src94 <= 16'h257;
        src95 <= 16'h9864;
        src96 <= 16'hbea;
        src97 <= 16'h91ec;
        src98 <= 16'ha2f8;
        src99 <= 16'h8085;
        src100 <= 16'h217c;
        src101 <= 16'had44;
        src102 <= 16'h9db4;
        src103 <= 16'hc669;
        src104 <= 16'h1bac;
        src105 <= 16'h1b64;
        src106 <= 16'h96dd;
        src107 <= 16'h5d93;
        src108 <= 16'h688a;
        src109 <= 16'hf20c;
        src110 <= 16'h507;
        src111 <= 16'hfc47;
        src112 <= 16'h5312;
        src113 <= 16'h58df;
        src114 <= 16'h8f84;
        src115 <= 16'h288d;
        src116 <= 16'hbce5;
        src117 <= 16'h631c;
        src118 <= 16'hb352;
        src119 <= 16'hc91b;
        src120 <= 16'he27;
        src121 <= 16'hb399;
        src122 <= 16'ha8ea;
        src123 <= 16'h7716;
        src124 <= 16'h424;
        src125 <= 16'h91ee;
        src126 <= 16'h6f27;
        src127 <= 16'hbef7;
        src128 <= 16'he905;
        src129 <= 16'h8b72;
        src130 <= 16'ha9e7;
        src131 <= 16'hf7af;
        src132 <= 16'h5ce8;
        src133 <= 16'ha034;
        src134 <= 16'h924a;
        src135 <= 16'hf1c8;
        src136 <= 16'hed1;
        src137 <= 16'hfd40;
        src138 <= 16'h3c49;
        src139 <= 16'h54af;
        src140 <= 16'hd21;
        src141 <= 16'h332c;
        src142 <= 16'h69c4;
        src143 <= 16'ha28b;
        src144 <= 16'h8aa2;
        src145 <= 16'h62ac;
        src146 <= 16'hc650;
        src147 <= 16'h5be8;
        src148 <= 16'h12c7;
        src149 <= 16'h286;
        src150 <= 16'hfeb1;
        src151 <= 16'h723;
        src152 <= 16'h5369;
        src153 <= 16'hefa8;
        src154 <= 16'he97a;
        src155 <= 16'hac1e;
        src156 <= 16'he725;
        src157 <= 16'h95ea;
        src158 <= 16'hc6f8;
        src159 <= 16'h4318;
        src160 <= 16'hf126;
        src161 <= 16'h2130;
        src162 <= 16'h8455;
        src163 <= 16'h54fe;
        src164 <= 16'h4f52;
        src165 <= 16'h7abd;
        src166 <= 16'h7cf3;
        src167 <= 16'hc124;
        src168 <= 16'h1260;
        src169 <= 16'h9702;
        src170 <= 16'h8620;
        src171 <= 16'h801b;
        src172 <= 16'h5683;
        src173 <= 16'h545f;
        src174 <= 16'h837a;
        src175 <= 16'h7acc;
        src176 <= 16'he18f;
        src177 <= 16'h171d;
        src178 <= 16'h2dc4;
        src179 <= 16'hd66d;
        src180 <= 16'h21c0;
        src181 <= 16'hb629;
        src182 <= 16'h189f;
        src183 <= 16'h20df;
        src184 <= 16'h8455;
        exp <= 24'h5bc53c;
        #1
        src0 <= 16'h8b0f;
        src1 <= 16'ha693;
        src2 <= 16'h6daa;
        src3 <= 16'hb1ad;
        src4 <= 16'h4c65;
        src5 <= 16'hf118;
        src6 <= 16'h12dc;
        src7 <= 16'h4c20;
        src8 <= 16'hdba4;
        src9 <= 16'hf304;
        src10 <= 16'ha118;
        src11 <= 16'h8248;
        src12 <= 16'hf713;
        src13 <= 16'h5710;
        src14 <= 16'h6307;
        src15 <= 16'h490e;
        src16 <= 16'h45a0;
        src17 <= 16'haec;
        src18 <= 16'h6496;
        src19 <= 16'hf018;
        src20 <= 16'h92b3;
        src21 <= 16'h19d6;
        src22 <= 16'hc199;
        src23 <= 16'h4fca;
        src24 <= 16'h900a;
        src25 <= 16'hc880;
        src26 <= 16'h6bbd;
        src27 <= 16'h8cf3;
        src28 <= 16'he945;
        src29 <= 16'he207;
        src30 <= 16'h189c;
        src31 <= 16'h5021;
        src32 <= 16'hdd4d;
        src33 <= 16'ha7bd;
        src34 <= 16'h849d;
        src35 <= 16'h73d4;
        src36 <= 16'hbc08;
        src37 <= 16'hd81e;
        src38 <= 16'h82b7;
        src39 <= 16'hdcb3;
        src40 <= 16'h2e93;
        src41 <= 16'h1949;
        src42 <= 16'hab06;
        src43 <= 16'h88a6;
        src44 <= 16'hc0b5;
        src45 <= 16'h5e56;
        src46 <= 16'hd73a;
        src47 <= 16'ha683;
        src48 <= 16'h9975;
        src49 <= 16'h8c5e;
        src50 <= 16'h8e45;
        src51 <= 16'h8c76;
        src52 <= 16'h40e4;
        src53 <= 16'h9f08;
        src54 <= 16'ha5ea;
        src55 <= 16'hbcb9;
        src56 <= 16'hb629;
        src57 <= 16'h15f2;
        src58 <= 16'h384b;
        src59 <= 16'h60c5;
        src60 <= 16'hab68;
        src61 <= 16'he5c4;
        src62 <= 16'h2152;
        src63 <= 16'h515d;
        src64 <= 16'h80d0;
        src65 <= 16'h2514;
        src66 <= 16'h39f3;
        src67 <= 16'h81ae;
        src68 <= 16'h58b8;
        src69 <= 16'hdd95;
        src70 <= 16'h64c7;
        src71 <= 16'h382d;
        src72 <= 16'hcb3c;
        src73 <= 16'hc2b7;
        src74 <= 16'hcb54;
        src75 <= 16'h5fb4;
        src76 <= 16'hd68d;
        src77 <= 16'h4f6;
        src78 <= 16'h31a2;
        src79 <= 16'h65f8;
        src80 <= 16'he32d;
        src81 <= 16'hcf2f;
        src82 <= 16'h47f5;
        src83 <= 16'h78f6;
        src84 <= 16'h4372;
        src85 <= 16'h54d3;
        src86 <= 16'h5c7f;
        src87 <= 16'h97e0;
        src88 <= 16'ha830;
        src89 <= 16'h9b7f;
        src90 <= 16'hc00c;
        src91 <= 16'h58e5;
        src92 <= 16'hacac;
        src93 <= 16'hf0bd;
        src94 <= 16'h2967;
        src95 <= 16'heecb;
        src96 <= 16'hee1;
        src97 <= 16'h705c;
        src98 <= 16'h3d92;
        src99 <= 16'hd726;
        src100 <= 16'ha374;
        src101 <= 16'h5b53;
        src102 <= 16'h73f5;
        src103 <= 16'h2200;
        src104 <= 16'h28b4;
        src105 <= 16'hfeea;
        src106 <= 16'h435;
        src107 <= 16'hbff8;
        src108 <= 16'hd5c7;
        src109 <= 16'h3b23;
        src110 <= 16'hc3ff;
        src111 <= 16'h4c63;
        src112 <= 16'h8cb;
        src113 <= 16'h6460;
        src114 <= 16'h7a50;
        src115 <= 16'hdccd;
        src116 <= 16'h9ee0;
        src117 <= 16'h8ca;
        src118 <= 16'h9236;
        src119 <= 16'h6b07;
        src120 <= 16'h7606;
        src121 <= 16'h7a7d;
        src122 <= 16'hab86;
        src123 <= 16'h6c31;
        src124 <= 16'hd580;
        src125 <= 16'h8a2;
        src126 <= 16'hce61;
        src127 <= 16'h6fb2;
        src128 <= 16'h5966;
        src129 <= 16'h3508;
        src130 <= 16'h608f;
        src131 <= 16'h7218;
        src132 <= 16'h6f95;
        src133 <= 16'hca8f;
        src134 <= 16'h162d;
        src135 <= 16'h262e;
        src136 <= 16'h9399;
        src137 <= 16'h5e9f;
        src138 <= 16'h268c;
        src139 <= 16'ha286;
        src140 <= 16'hded9;
        src141 <= 16'h101d;
        src142 <= 16'h85fe;
        src143 <= 16'h8d43;
        src144 <= 16'hae28;
        src145 <= 16'hdfcc;
        src146 <= 16'h3c16;
        src147 <= 16'hf99;
        src148 <= 16'he110;
        src149 <= 16'h8b18;
        src150 <= 16'h24d7;
        src151 <= 16'h4cf7;
        src152 <= 16'hb615;
        src153 <= 16'h581e;
        src154 <= 16'h3d6b;
        src155 <= 16'hb586;
        src156 <= 16'he3a;
        src157 <= 16'hfd90;
        src158 <= 16'h8923;
        src159 <= 16'h1e9c;
        src160 <= 16'hbf57;
        src161 <= 16'hf15b;
        src162 <= 16'hee7e;
        src163 <= 16'h8e6b;
        src164 <= 16'hc1be;
        src165 <= 16'h4e7d;
        src166 <= 16'h4104;
        src167 <= 16'hfceb;
        src168 <= 16'h2ec;
        src169 <= 16'h7ab4;
        src170 <= 16'h2720;
        src171 <= 16'hcd0d;
        src172 <= 16'h8b23;
        src173 <= 16'h9461;
        src174 <= 16'h6b9a;
        src175 <= 16'h7369;
        src176 <= 16'h9114;
        src177 <= 16'h9f68;
        src178 <= 16'h716a;
        src179 <= 16'hc062;
        src180 <= 16'ha8fa;
        src181 <= 16'h841d;
        src182 <= 16'hf5a9;
        src183 <= 16'h951e;
        src184 <= 16'h16c2;
        exp <= 24'h5d8c5f;
        #1
        src0 <= 16'h87a8;
        src1 <= 16'h35e2;
        src2 <= 16'hc226;
        src3 <= 16'he921;
        src4 <= 16'hd1c8;
        src5 <= 16'h2f7e;
        src6 <= 16'h478a;
        src7 <= 16'hc7d;
        src8 <= 16'hb5e7;
        src9 <= 16'h4c04;
        src10 <= 16'h59;
        src11 <= 16'h10e6;
        src12 <= 16'h617d;
        src13 <= 16'h8233;
        src14 <= 16'h601f;
        src15 <= 16'h15fb;
        src16 <= 16'h7d92;
        src17 <= 16'hd752;
        src18 <= 16'hc4fc;
        src19 <= 16'h31e4;
        src20 <= 16'h7938;
        src21 <= 16'h262;
        src22 <= 16'h62ef;
        src23 <= 16'h4a84;
        src24 <= 16'h914e;
        src25 <= 16'hbf84;
        src26 <= 16'h4fe0;
        src27 <= 16'h9786;
        src28 <= 16'h5adc;
        src29 <= 16'h8722;
        src30 <= 16'h982d;
        src31 <= 16'hc82c;
        src32 <= 16'h7b9;
        src33 <= 16'h919b;
        src34 <= 16'h6cb5;
        src35 <= 16'hdcaf;
        src36 <= 16'hc7ae;
        src37 <= 16'hf5f9;
        src38 <= 16'h5289;
        src39 <= 16'hed6a;
        src40 <= 16'h14b5;
        src41 <= 16'h72da;
        src42 <= 16'hfea9;
        src43 <= 16'h513a;
        src44 <= 16'hc143;
        src45 <= 16'h9c0e;
        src46 <= 16'h4f69;
        src47 <= 16'h593;
        src48 <= 16'ha496;
        src49 <= 16'h6167;
        src50 <= 16'h1192;
        src51 <= 16'hc16f;
        src52 <= 16'hefc7;
        src53 <= 16'h6ac3;
        src54 <= 16'hf856;
        src55 <= 16'h736e;
        src56 <= 16'hf411;
        src57 <= 16'h8f0;
        src58 <= 16'hce07;
        src59 <= 16'hd6d1;
        src60 <= 16'hc077;
        src61 <= 16'h2379;
        src62 <= 16'h5542;
        src63 <= 16'hb67b;
        src64 <= 16'hc199;
        src65 <= 16'hc17f;
        src66 <= 16'hf43;
        src67 <= 16'hbbbf;
        src68 <= 16'h156c;
        src69 <= 16'hcee8;
        src70 <= 16'h6777;
        src71 <= 16'hedf9;
        src72 <= 16'h7e54;
        src73 <= 16'h75fb;
        src74 <= 16'h9b8;
        src75 <= 16'had;
        src76 <= 16'haa2f;
        src77 <= 16'h5a54;
        src78 <= 16'h5c3d;
        src79 <= 16'h88c0;
        src80 <= 16'h12e3;
        src81 <= 16'h9f30;
        src82 <= 16'h9d2f;
        src83 <= 16'h72ea;
        src84 <= 16'h3db9;
        src85 <= 16'he89c;
        src86 <= 16'h267;
        src87 <= 16'h7f55;
        src88 <= 16'h17a7;
        src89 <= 16'ha374;
        src90 <= 16'h346a;
        src91 <= 16'he535;
        src92 <= 16'h5496;
        src93 <= 16'h349c;
        src94 <= 16'hbb49;
        src95 <= 16'h6d43;
        src96 <= 16'h700f;
        src97 <= 16'h506f;
        src98 <= 16'hb8a6;
        src99 <= 16'ha913;
        src100 <= 16'h196a;
        src101 <= 16'h83ba;
        src102 <= 16'hf17c;
        src103 <= 16'h1b47;
        src104 <= 16'h4e41;
        src105 <= 16'hbc7;
        src106 <= 16'hf058;
        src107 <= 16'ha1f1;
        src108 <= 16'h78af;
        src109 <= 16'h49ca;
        src110 <= 16'h1a05;
        src111 <= 16'he884;
        src112 <= 16'h7b0a;
        src113 <= 16'h1e01;
        src114 <= 16'hc3be;
        src115 <= 16'he91d;
        src116 <= 16'h4e8e;
        src117 <= 16'haee7;
        src118 <= 16'hf6f8;
        src119 <= 16'h61ad;
        src120 <= 16'h1b56;
        src121 <= 16'h5793;
        src122 <= 16'hf6db;
        src123 <= 16'h46a5;
        src124 <= 16'ha8c2;
        src125 <= 16'ha1f9;
        src126 <= 16'h5518;
        src127 <= 16'hb6f8;
        src128 <= 16'h9df6;
        src129 <= 16'h32a8;
        src130 <= 16'h456;
        src131 <= 16'hcdba;
        src132 <= 16'h23b4;
        src133 <= 16'hcfb0;
        src134 <= 16'h44aa;
        src135 <= 16'h86d8;
        src136 <= 16'hc9af;
        src137 <= 16'hda6b;
        src138 <= 16'hb674;
        src139 <= 16'hf4b2;
        src140 <= 16'h3f8b;
        src141 <= 16'hfa77;
        src142 <= 16'habac;
        src143 <= 16'hd01e;
        src144 <= 16'hb7da;
        src145 <= 16'ha1cc;
        src146 <= 16'h41a7;
        src147 <= 16'h9825;
        src148 <= 16'h558f;
        src149 <= 16'h3931;
        src150 <= 16'h8e81;
        src151 <= 16'h54c8;
        src152 <= 16'h16f6;
        src153 <= 16'hed4;
        src154 <= 16'h4d44;
        src155 <= 16'h77c5;
        src156 <= 16'h4754;
        src157 <= 16'h6e7f;
        src158 <= 16'h11c0;
        src159 <= 16'hd215;
        src160 <= 16'h7e80;
        src161 <= 16'hd53c;
        src162 <= 16'h7315;
        src163 <= 16'h7ff7;
        src164 <= 16'h40c0;
        src165 <= 16'hc117;
        src166 <= 16'h96b4;
        src167 <= 16'h9375;
        src168 <= 16'h5e51;
        src169 <= 16'h37a;
        src170 <= 16'h4833;
        src171 <= 16'h91fb;
        src172 <= 16'h5e92;
        src173 <= 16'h61b5;
        src174 <= 16'hc590;
        src175 <= 16'h2e3f;
        src176 <= 16'h7d77;
        src177 <= 16'h4b32;
        src178 <= 16'h5148;
        src179 <= 16'hc092;
        src180 <= 16'hc87;
        src181 <= 16'h3b8a;
        src182 <= 16'h15b;
        src183 <= 16'h8c19;
        src184 <= 16'h172a;
        exp <= 24'h57f160;
        #1
        src0 <= 16'h565;
        src1 <= 16'h1e71;
        src2 <= 16'h23ae;
        src3 <= 16'hf1e7;
        src4 <= 16'hc09f;
        src5 <= 16'h49c0;
        src6 <= 16'h571e;
        src7 <= 16'hbac2;
        src8 <= 16'hdc3e;
        src9 <= 16'h912a;
        src10 <= 16'h718c;
        src11 <= 16'hc88;
        src12 <= 16'hfe6b;
        src13 <= 16'ha8fd;
        src14 <= 16'hfd6;
        src15 <= 16'h18eb;
        src16 <= 16'h671b;
        src17 <= 16'he58e;
        src18 <= 16'haabf;
        src19 <= 16'h990f;
        src20 <= 16'h3190;
        src21 <= 16'hb57f;
        src22 <= 16'h6e6f;
        src23 <= 16'h555e;
        src24 <= 16'ha3d4;
        src25 <= 16'ha903;
        src26 <= 16'hefac;
        src27 <= 16'h5125;
        src28 <= 16'hc63c;
        src29 <= 16'ha323;
        src30 <= 16'h592c;
        src31 <= 16'h75fe;
        src32 <= 16'h6a3d;
        src33 <= 16'hcc03;
        src34 <= 16'h7e58;
        src35 <= 16'h6949;
        src36 <= 16'h77fc;
        src37 <= 16'h5c4d;
        src38 <= 16'hbb13;
        src39 <= 16'h3e61;
        src40 <= 16'h125e;
        src41 <= 16'he000;
        src42 <= 16'ha312;
        src43 <= 16'h1e54;
        src44 <= 16'h3e6;
        src45 <= 16'hb5ae;
        src46 <= 16'h1749;
        src47 <= 16'hd287;
        src48 <= 16'hb439;
        src49 <= 16'hf1d3;
        src50 <= 16'hc98e;
        src51 <= 16'hddbc;
        src52 <= 16'h3b6b;
        src53 <= 16'he211;
        src54 <= 16'h270d;
        src55 <= 16'hb0ff;
        src56 <= 16'h1aab;
        src57 <= 16'hb48d;
        src58 <= 16'hae1a;
        src59 <= 16'hab0c;
        src60 <= 16'hb426;
        src61 <= 16'h6ef2;
        src62 <= 16'h6d85;
        src63 <= 16'hab2e;
        src64 <= 16'h5c5e;
        src65 <= 16'hc99d;
        src66 <= 16'h1285;
        src67 <= 16'hbf7;
        src68 <= 16'h7bb1;
        src69 <= 16'h17b9;
        src70 <= 16'hd33b;
        src71 <= 16'h976b;
        src72 <= 16'h2557;
        src73 <= 16'he13e;
        src74 <= 16'h8de3;
        src75 <= 16'h65bf;
        src76 <= 16'h407c;
        src77 <= 16'h4ed9;
        src78 <= 16'h40c7;
        src79 <= 16'h271a;
        src80 <= 16'h5e0f;
        src81 <= 16'h9c63;
        src82 <= 16'he3c3;
        src83 <= 16'h1152;
        src84 <= 16'h5812;
        src85 <= 16'haf9d;
        src86 <= 16'hb94f;
        src87 <= 16'h9118;
        src88 <= 16'hc527;
        src89 <= 16'h8fdc;
        src90 <= 16'haf16;
        src91 <= 16'hdd4e;
        src92 <= 16'h5f31;
        src93 <= 16'h61b3;
        src94 <= 16'h78c3;
        src95 <= 16'he2;
        src96 <= 16'hfc6a;
        src97 <= 16'h16dd;
        src98 <= 16'h6c5c;
        src99 <= 16'h5be;
        src100 <= 16'h8b05;
        src101 <= 16'hc235;
        src102 <= 16'hde32;
        src103 <= 16'h7bc2;
        src104 <= 16'ha239;
        src105 <= 16'hadbb;
        src106 <= 16'h972a;
        src107 <= 16'h4c67;
        src108 <= 16'hd762;
        src109 <= 16'he827;
        src110 <= 16'h72cc;
        src111 <= 16'h28f2;
        src112 <= 16'h661d;
        src113 <= 16'hf5ac;
        src114 <= 16'h6f27;
        src115 <= 16'hb45d;
        src116 <= 16'he720;
        src117 <= 16'h6cf9;
        src118 <= 16'h9921;
        src119 <= 16'h65ca;
        src120 <= 16'h3acc;
        src121 <= 16'hcb06;
        src122 <= 16'h9b0f;
        src123 <= 16'h70a6;
        src124 <= 16'h342;
        src125 <= 16'h6ab1;
        src126 <= 16'hd13a;
        src127 <= 16'hf2cd;
        src128 <= 16'h5b56;
        src129 <= 16'h81f1;
        src130 <= 16'h45a4;
        src131 <= 16'h42ae;
        src132 <= 16'h567b;
        src133 <= 16'h4f2b;
        src134 <= 16'hd21f;
        src135 <= 16'hb302;
        src136 <= 16'h1354;
        src137 <= 16'h9894;
        src138 <= 16'hb6be;
        src139 <= 16'h6de8;
        src140 <= 16'h1012;
        src141 <= 16'h31ab;
        src142 <= 16'hd4db;
        src143 <= 16'h9ece;
        src144 <= 16'h763;
        src145 <= 16'h1e81;
        src146 <= 16'hf241;
        src147 <= 16'h5dc4;
        src148 <= 16'h9984;
        src149 <= 16'h1e3c;
        src150 <= 16'h228a;
        src151 <= 16'h3641;
        src152 <= 16'hbff3;
        src153 <= 16'h4da9;
        src154 <= 16'hc095;
        src155 <= 16'h8f1a;
        src156 <= 16'h12a5;
        src157 <= 16'h2beb;
        src158 <= 16'h605a;
        src159 <= 16'h15bc;
        src160 <= 16'h353;
        src161 <= 16'h271c;
        src162 <= 16'hbf18;
        src163 <= 16'ha50b;
        src164 <= 16'h5e2d;
        src165 <= 16'hdb59;
        src166 <= 16'h4b70;
        src167 <= 16'hf8dc;
        src168 <= 16'hc0a0;
        src169 <= 16'hb573;
        src170 <= 16'hc1f4;
        src171 <= 16'ha056;
        src172 <= 16'h999b;
        src173 <= 16'h26f8;
        src174 <= 16'h3505;
        src175 <= 16'hee96;
        src176 <= 16'ha0dd;
        src177 <= 16'hca5d;
        src178 <= 16'hb636;
        src179 <= 16'h6b0b;
        src180 <= 16'h92;
        src181 <= 16'had68;
        src182 <= 16'h1735;
        src183 <= 16'h87e8;
        src184 <= 16'h84dd;
        exp <= 24'h5b3565;
        #1
        src0 <= 16'hbbfb;
        src1 <= 16'h8f4f;
        src2 <= 16'h14db;
        src3 <= 16'h6cba;
        src4 <= 16'hc7f7;
        src5 <= 16'hb082;
        src6 <= 16'h55be;
        src7 <= 16'h9f94;
        src8 <= 16'h3334;
        src9 <= 16'h21c7;
        src10 <= 16'h73d1;
        src11 <= 16'h9db0;
        src12 <= 16'h6258;
        src13 <= 16'hddd2;
        src14 <= 16'h34c2;
        src15 <= 16'hc842;
        src16 <= 16'h1b27;
        src17 <= 16'h33fc;
        src18 <= 16'h12ea;
        src19 <= 16'h3ded;
        src20 <= 16'h8ccd;
        src21 <= 16'h43c7;
        src22 <= 16'hd322;
        src23 <= 16'h8243;
        src24 <= 16'h55bb;
        src25 <= 16'he421;
        src26 <= 16'h4500;
        src27 <= 16'h582b;
        src28 <= 16'h8e6f;
        src29 <= 16'h5156;
        src30 <= 16'hd4c4;
        src31 <= 16'h7320;
        src32 <= 16'h446c;
        src33 <= 16'h3047;
        src34 <= 16'h5cba;
        src35 <= 16'h5aa3;
        src36 <= 16'h723;
        src37 <= 16'h1081;
        src38 <= 16'h8a5a;
        src39 <= 16'hab07;
        src40 <= 16'hddcf;
        src41 <= 16'hcea3;
        src42 <= 16'hd00a;
        src43 <= 16'hdd7b;
        src44 <= 16'ha2ff;
        src45 <= 16'he347;
        src46 <= 16'h6e67;
        src47 <= 16'h5b23;
        src48 <= 16'h803;
        src49 <= 16'h62e4;
        src50 <= 16'h732e;
        src51 <= 16'h2a5d;
        src52 <= 16'he488;
        src53 <= 16'hb1d3;
        src54 <= 16'h53c3;
        src55 <= 16'hd8b0;
        src56 <= 16'h2f6a;
        src57 <= 16'hde70;
        src58 <= 16'h793a;
        src59 <= 16'hf980;
        src60 <= 16'h9da5;
        src61 <= 16'h3aed;
        src62 <= 16'h4ac0;
        src63 <= 16'hd6c5;
        src64 <= 16'h88de;
        src65 <= 16'h58a7;
        src66 <= 16'h5adb;
        src67 <= 16'heb58;
        src68 <= 16'h3fbc;
        src69 <= 16'h3e50;
        src70 <= 16'hdc7f;
        src71 <= 16'hb809;
        src72 <= 16'hcc92;
        src73 <= 16'hfe99;
        src74 <= 16'h2b4a;
        src75 <= 16'h3f6d;
        src76 <= 16'he134;
        src77 <= 16'hf5ab;
        src78 <= 16'h25b2;
        src79 <= 16'h9f2e;
        src80 <= 16'h1f0;
        src81 <= 16'h4b0e;
        src82 <= 16'h95ce;
        src83 <= 16'h51b6;
        src84 <= 16'hac7d;
        src85 <= 16'h1f20;
        src86 <= 16'h1f99;
        src87 <= 16'hf94a;
        src88 <= 16'hf7aa;
        src89 <= 16'h941c;
        src90 <= 16'hb9b3;
        src91 <= 16'h8388;
        src92 <= 16'h3d;
        src93 <= 16'ha73d;
        src94 <= 16'h6fed;
        src95 <= 16'h8248;
        src96 <= 16'h6cea;
        src97 <= 16'h5368;
        src98 <= 16'h5b47;
        src99 <= 16'h603;
        src100 <= 16'h9cfb;
        src101 <= 16'h64;
        src102 <= 16'h793;
        src103 <= 16'h63db;
        src104 <= 16'h181c;
        src105 <= 16'h571c;
        src106 <= 16'h37ed;
        src107 <= 16'h310d;
        src108 <= 16'hfbc2;
        src109 <= 16'hb5d3;
        src110 <= 16'he482;
        src111 <= 16'h9fcb;
        src112 <= 16'h3d0d;
        src113 <= 16'h5891;
        src114 <= 16'h957f;
        src115 <= 16'h4501;
        src116 <= 16'hf129;
        src117 <= 16'h13a1;
        src118 <= 16'ha968;
        src119 <= 16'h74ad;
        src120 <= 16'h9245;
        src121 <= 16'hfb09;
        src122 <= 16'hf6ee;
        src123 <= 16'hff42;
        src124 <= 16'h41a0;
        src125 <= 16'h1b0;
        src126 <= 16'hdb43;
        src127 <= 16'hfc2b;
        src128 <= 16'h1457;
        src129 <= 16'h4b53;
        src130 <= 16'h8290;
        src131 <= 16'h3560;
        src132 <= 16'h8173;
        src133 <= 16'h2731;
        src134 <= 16'hec5f;
        src135 <= 16'hcb90;
        src136 <= 16'h1d2a;
        src137 <= 16'h47cc;
        src138 <= 16'h1b71;
        src139 <= 16'h5aa2;
        src140 <= 16'haea7;
        src141 <= 16'he509;
        src142 <= 16'he4af;
        src143 <= 16'head6;
        src144 <= 16'h4a18;
        src145 <= 16'ha96;
        src146 <= 16'haf5f;
        src147 <= 16'h11d0;
        src148 <= 16'h46bc;
        src149 <= 16'h73f4;
        src150 <= 16'ha310;
        src151 <= 16'h1d27;
        src152 <= 16'h36f4;
        src153 <= 16'hccd7;
        src154 <= 16'h1d68;
        src155 <= 16'h9588;
        src156 <= 16'hb2d8;
        src157 <= 16'ha18e;
        src158 <= 16'hbff7;
        src159 <= 16'h5311;
        src160 <= 16'h6414;
        src161 <= 16'h8691;
        src162 <= 16'hc452;
        src163 <= 16'h5861;
        src164 <= 16'h7933;
        src165 <= 16'ha78b;
        src166 <= 16'hcf92;
        src167 <= 16'hd69b;
        src168 <= 16'h7099;
        src169 <= 16'ha8ea;
        src170 <= 16'h8684;
        src171 <= 16'h596;
        src172 <= 16'h1cbd;
        src173 <= 16'hd6fe;
        src174 <= 16'hdbaa;
        src175 <= 16'h7e9;
        src176 <= 16'h8f61;
        src177 <= 16'h6d9f;
        src178 <= 16'he195;
        src179 <= 16'h29a;
        src180 <= 16'h1c55;
        src181 <= 16'hb223;
        src182 <= 16'he2f0;
        src183 <= 16'h471f;
        src184 <= 16'hf7fd;
        exp <= 24'h5a7f4c;
        #1
        src0 <= 16'h6b41;
        src1 <= 16'ha867;
        src2 <= 16'hb612;
        src3 <= 16'h50e4;
        src4 <= 16'h7f0c;
        src5 <= 16'ha0cb;
        src6 <= 16'h8799;
        src7 <= 16'h170e;
        src8 <= 16'h9292;
        src9 <= 16'h6098;
        src10 <= 16'h2c66;
        src11 <= 16'h6534;
        src12 <= 16'hfe05;
        src13 <= 16'ha1bf;
        src14 <= 16'h76ef;
        src15 <= 16'h6feb;
        src16 <= 16'h41df;
        src17 <= 16'h2ecd;
        src18 <= 16'h8924;
        src19 <= 16'h901f;
        src20 <= 16'h1fe9;
        src21 <= 16'h4de2;
        src22 <= 16'ha7b2;
        src23 <= 16'h7062;
        src24 <= 16'h1d05;
        src25 <= 16'h20c6;
        src26 <= 16'h5698;
        src27 <= 16'hf592;
        src28 <= 16'h7174;
        src29 <= 16'h7d3;
        src30 <= 16'hcebc;
        src31 <= 16'h775d;
        src32 <= 16'h198c;
        src33 <= 16'he1d7;
        src34 <= 16'h8191;
        src35 <= 16'h4d97;
        src36 <= 16'h6491;
        src37 <= 16'h483c;
        src38 <= 16'hb479;
        src39 <= 16'h9896;
        src40 <= 16'h1ffc;
        src41 <= 16'h6778;
        src42 <= 16'h85cb;
        src43 <= 16'hdfaf;
        src44 <= 16'h7f96;
        src45 <= 16'h613e;
        src46 <= 16'he334;
        src47 <= 16'hf389;
        src48 <= 16'h4a60;
        src49 <= 16'h7f65;
        src50 <= 16'h8c75;
        src51 <= 16'hd8a2;
        src52 <= 16'h17d7;
        src53 <= 16'hddc1;
        src54 <= 16'h8bfd;
        src55 <= 16'h72a3;
        src56 <= 16'h78ac;
        src57 <= 16'h22a6;
        src58 <= 16'hb458;
        src59 <= 16'h2630;
        src60 <= 16'h1995;
        src61 <= 16'h5bd8;
        src62 <= 16'ha3e5;
        src63 <= 16'h3782;
        src64 <= 16'ha9a6;
        src65 <= 16'h96f2;
        src66 <= 16'h6f18;
        src67 <= 16'hd112;
        src68 <= 16'hb9c2;
        src69 <= 16'hbd57;
        src70 <= 16'he708;
        src71 <= 16'h692f;
        src72 <= 16'h6e39;
        src73 <= 16'h9b62;
        src74 <= 16'h383d;
        src75 <= 16'h29df;
        src76 <= 16'he3cb;
        src77 <= 16'h43bd;
        src78 <= 16'hd09;
        src79 <= 16'h2dbc;
        src80 <= 16'h491d;
        src81 <= 16'h6580;
        src82 <= 16'hff23;
        src83 <= 16'hbeb8;
        src84 <= 16'h6f85;
        src85 <= 16'h60d;
        src86 <= 16'hce5b;
        src87 <= 16'he33e;
        src88 <= 16'he6b7;
        src89 <= 16'h16c3;
        src90 <= 16'hcc14;
        src91 <= 16'h57e7;
        src92 <= 16'h6ced;
        src93 <= 16'hc92d;
        src94 <= 16'h35c;
        src95 <= 16'h826;
        src96 <= 16'hd868;
        src97 <= 16'h4246;
        src98 <= 16'hda0f;
        src99 <= 16'h2a0d;
        src100 <= 16'h2a89;
        src101 <= 16'h5501;
        src102 <= 16'hfcb2;
        src103 <= 16'h5909;
        src104 <= 16'hfca1;
        src105 <= 16'he40;
        src106 <= 16'hb244;
        src107 <= 16'h8a7e;
        src108 <= 16'h9597;
        src109 <= 16'hcd4c;
        src110 <= 16'h4b08;
        src111 <= 16'hf67f;
        src112 <= 16'h1ccf;
        src113 <= 16'h4a0b;
        src114 <= 16'h11dd;
        src115 <= 16'h92ce;
        src116 <= 16'h6b14;
        src117 <= 16'h1be9;
        src118 <= 16'hef78;
        src119 <= 16'h1c6c;
        src120 <= 16'hea19;
        src121 <= 16'h642c;
        src122 <= 16'h8b63;
        src123 <= 16'hf5eb;
        src124 <= 16'h22be;
        src125 <= 16'hf663;
        src126 <= 16'h1893;
        src127 <= 16'hfa5b;
        src128 <= 16'h65ae;
        src129 <= 16'h3852;
        src130 <= 16'h12aa;
        src131 <= 16'h8f54;
        src132 <= 16'hd3f8;
        src133 <= 16'h5deb;
        src134 <= 16'h74dc;
        src135 <= 16'h4d34;
        src136 <= 16'hfecc;
        src137 <= 16'hff68;
        src138 <= 16'h12f6;
        src139 <= 16'hd7;
        src140 <= 16'h3ae0;
        src141 <= 16'h526f;
        src142 <= 16'ha118;
        src143 <= 16'h2ed9;
        src144 <= 16'he9aa;
        src145 <= 16'hf8ee;
        src146 <= 16'h5335;
        src147 <= 16'hc2f8;
        src148 <= 16'hd2b5;
        src149 <= 16'ha937;
        src150 <= 16'h5ab0;
        src151 <= 16'hd0aa;
        src152 <= 16'h5da4;
        src153 <= 16'h82ad;
        src154 <= 16'h24b2;
        src155 <= 16'h3765;
        src156 <= 16'hf41d;
        src157 <= 16'haf0a;
        src158 <= 16'hca55;
        src159 <= 16'h8435;
        src160 <= 16'h4241;
        src161 <= 16'h8151;
        src162 <= 16'h3d45;
        src163 <= 16'hd050;
        src164 <= 16'ha947;
        src165 <= 16'h94f4;
        src166 <= 16'hb90d;
        src167 <= 16'hc7ab;
        src168 <= 16'hd7fb;
        src169 <= 16'hdc2d;
        src170 <= 16'h31a6;
        src171 <= 16'h8f10;
        src172 <= 16'h4b2e;
        src173 <= 16'ha0a3;
        src174 <= 16'hf06f;
        src175 <= 16'h6315;
        src176 <= 16'h6d90;
        src177 <= 16'h8b7a;
        src178 <= 16'h26a2;
        src179 <= 16'h18aa;
        src180 <= 16'hfd7b;
        src181 <= 16'ha1e3;
        src182 <= 16'h9ffc;
        src183 <= 16'h4ba4;
        src184 <= 16'h3b01;
        exp <= 24'h5bcb2f;
        #1
        src0 <= 16'h6b9b;
        src1 <= 16'h3f38;
        src2 <= 16'h28f7;
        src3 <= 16'h6326;
        src4 <= 16'h9955;
        src5 <= 16'hd733;
        src6 <= 16'hc5c8;
        src7 <= 16'h2087;
        src8 <= 16'h39e5;
        src9 <= 16'h3f08;
        src10 <= 16'h48b5;
        src11 <= 16'h138f;
        src12 <= 16'h4251;
        src13 <= 16'hdee7;
        src14 <= 16'he305;
        src15 <= 16'h1e24;
        src16 <= 16'h4b9;
        src17 <= 16'hff92;
        src18 <= 16'h4154;
        src19 <= 16'hc97f;
        src20 <= 16'hbf6b;
        src21 <= 16'h8676;
        src22 <= 16'h1fa1;
        src23 <= 16'hb886;
        src24 <= 16'h920d;
        src25 <= 16'hec2e;
        src26 <= 16'hb610;
        src27 <= 16'hc6db;
        src28 <= 16'h2903;
        src29 <= 16'hb014;
        src30 <= 16'hcfaf;
        src31 <= 16'ha114;
        src32 <= 16'hb209;
        src33 <= 16'h3fe1;
        src34 <= 16'h8858;
        src35 <= 16'hd34e;
        src36 <= 16'hbac8;
        src37 <= 16'hc4eb;
        src38 <= 16'h8578;
        src39 <= 16'h840a;
        src40 <= 16'hbb6f;
        src41 <= 16'hc7c7;
        src42 <= 16'h4164;
        src43 <= 16'h8b25;
        src44 <= 16'h2d5e;
        src45 <= 16'h44c8;
        src46 <= 16'hbf37;
        src47 <= 16'hf432;
        src48 <= 16'hd9a9;
        src49 <= 16'h4920;
        src50 <= 16'h4162;
        src51 <= 16'h8606;
        src52 <= 16'hcb16;
        src53 <= 16'hec49;
        src54 <= 16'hf53e;
        src55 <= 16'h6317;
        src56 <= 16'h53b;
        src57 <= 16'h6493;
        src58 <= 16'hbdbb;
        src59 <= 16'hc76b;
        src60 <= 16'he42a;
        src61 <= 16'h5e34;
        src62 <= 16'h9f49;
        src63 <= 16'hb8ec;
        src64 <= 16'h644b;
        src65 <= 16'h97e2;
        src66 <= 16'hfc03;
        src67 <= 16'h2eee;
        src68 <= 16'h2265;
        src69 <= 16'hf32e;
        src70 <= 16'hc826;
        src71 <= 16'hebc5;
        src72 <= 16'ha22;
        src73 <= 16'h6e97;
        src74 <= 16'h1a94;
        src75 <= 16'h3805;
        src76 <= 16'h8aee;
        src77 <= 16'h7d64;
        src78 <= 16'habb5;
        src79 <= 16'hb8fb;
        src80 <= 16'h2e4;
        src81 <= 16'h5ceb;
        src82 <= 16'h3c1d;
        src83 <= 16'hce06;
        src84 <= 16'hc467;
        src85 <= 16'hf93e;
        src86 <= 16'h3e08;
        src87 <= 16'h2e7e;
        src88 <= 16'h3233;
        src89 <= 16'h4103;
        src90 <= 16'he48b;
        src91 <= 16'h61ae;
        src92 <= 16'h951e;
        src93 <= 16'h62f1;
        src94 <= 16'h511e;
        src95 <= 16'hfc24;
        src96 <= 16'hf35e;
        src97 <= 16'h82fa;
        src98 <= 16'h8589;
        src99 <= 16'h63a3;
        src100 <= 16'h5fbc;
        src101 <= 16'hc15c;
        src102 <= 16'h781a;
        src103 <= 16'h11b6;
        src104 <= 16'hcdfb;
        src105 <= 16'h6ce0;
        src106 <= 16'h2c52;
        src107 <= 16'h89c1;
        src108 <= 16'h1ba8;
        src109 <= 16'ha20d;
        src110 <= 16'h44c9;
        src111 <= 16'h58bf;
        src112 <= 16'h673;
        src113 <= 16'h1e21;
        src114 <= 16'h27b3;
        src115 <= 16'h604c;
        src116 <= 16'hdd8a;
        src117 <= 16'h6387;
        src118 <= 16'h992d;
        src119 <= 16'h46a6;
        src120 <= 16'hc98;
        src121 <= 16'hcc3a;
        src122 <= 16'h37d0;
        src123 <= 16'h11b;
        src124 <= 16'h5026;
        src125 <= 16'h1a19;
        src126 <= 16'h7d81;
        src127 <= 16'h3af9;
        src128 <= 16'hf8d3;
        src129 <= 16'ha73f;
        src130 <= 16'h870;
        src131 <= 16'hb3cb;
        src132 <= 16'hb62a;
        src133 <= 16'hbb4d;
        src134 <= 16'h5452;
        src135 <= 16'h7032;
        src136 <= 16'h53a2;
        src137 <= 16'h3873;
        src138 <= 16'h522e;
        src139 <= 16'h8793;
        src140 <= 16'h6f5f;
        src141 <= 16'hc608;
        src142 <= 16'hccfd;
        src143 <= 16'h7ea8;
        src144 <= 16'h1ba9;
        src145 <= 16'h50b7;
        src146 <= 16'h8084;
        src147 <= 16'hcdc8;
        src148 <= 16'ha90c;
        src149 <= 16'h5d3a;
        src150 <= 16'h48e7;
        src151 <= 16'h7f11;
        src152 <= 16'h1790;
        src153 <= 16'h7c3c;
        src154 <= 16'h7074;
        src155 <= 16'hac74;
        src156 <= 16'h9b4e;
        src157 <= 16'h553a;
        src158 <= 16'h9208;
        src159 <= 16'hfc3c;
        src160 <= 16'hec18;
        src161 <= 16'hb9bb;
        src162 <= 16'hcc5c;
        src163 <= 16'habf5;
        src164 <= 16'h5f66;
        src165 <= 16'h9e46;
        src166 <= 16'h14c4;
        src167 <= 16'h8e66;
        src168 <= 16'h4e47;
        src169 <= 16'h8c26;
        src170 <= 16'h672a;
        src171 <= 16'h45c8;
        src172 <= 16'h79f;
        src173 <= 16'h6dc2;
        src174 <= 16'hf08c;
        src175 <= 16'hd80e;
        src176 <= 16'h5d3c;
        src177 <= 16'h44b8;
        src178 <= 16'h7b3a;
        src179 <= 16'h75ef;
        src180 <= 16'h4b96;
        src181 <= 16'h591f;
        src182 <= 16'h85ad;
        src183 <= 16'h9d92;
        src184 <= 16'h1338;
        exp <= 24'h5aff80;
        #1
        src0 <= 16'h73c6;
        src1 <= 16'h3a2;
        src2 <= 16'h7a69;
        src3 <= 16'h5e83;
        src4 <= 16'hf526;
        src5 <= 16'hd008;
        src6 <= 16'h7a37;
        src7 <= 16'hf2c2;
        src8 <= 16'hde3b;
        src9 <= 16'hb8ea;
        src10 <= 16'h273e;
        src11 <= 16'h3782;
        src12 <= 16'h14de;
        src13 <= 16'hbf8e;
        src14 <= 16'h77a0;
        src15 <= 16'h81a6;
        src16 <= 16'hfc41;
        src17 <= 16'h5da8;
        src18 <= 16'hc367;
        src19 <= 16'hf128;
        src20 <= 16'h5d6;
        src21 <= 16'h7285;
        src22 <= 16'h6b01;
        src23 <= 16'h1d09;
        src24 <= 16'hb3fd;
        src25 <= 16'h491b;
        src26 <= 16'ha264;
        src27 <= 16'he2d4;
        src28 <= 16'h4f7f;
        src29 <= 16'hf4ec;
        src30 <= 16'haa82;
        src31 <= 16'h9430;
        src32 <= 16'hf445;
        src33 <= 16'h5498;
        src34 <= 16'h5cd5;
        src35 <= 16'hb381;
        src36 <= 16'hbd44;
        src37 <= 16'h3b20;
        src38 <= 16'h78a4;
        src39 <= 16'h57ca;
        src40 <= 16'hb773;
        src41 <= 16'ha463;
        src42 <= 16'h6e77;
        src43 <= 16'hcb35;
        src44 <= 16'h85f7;
        src45 <= 16'h383;
        src46 <= 16'hba67;
        src47 <= 16'hde8c;
        src48 <= 16'hd9cd;
        src49 <= 16'hbf56;
        src50 <= 16'hd3b;
        src51 <= 16'h96d3;
        src52 <= 16'h62c1;
        src53 <= 16'h53;
        src54 <= 16'h9fb6;
        src55 <= 16'hc390;
        src56 <= 16'hbdf6;
        src57 <= 16'hd722;
        src58 <= 16'h6448;
        src59 <= 16'hfa90;
        src60 <= 16'h86a1;
        src61 <= 16'haf17;
        src62 <= 16'h6210;
        src63 <= 16'hf388;
        src64 <= 16'h2513;
        src65 <= 16'he151;
        src66 <= 16'h8551;
        src67 <= 16'hfa0c;
        src68 <= 16'h5318;
        src69 <= 16'h2993;
        src70 <= 16'hfb81;
        src71 <= 16'hb45a;
        src72 <= 16'hbae5;
        src73 <= 16'h3e76;
        src74 <= 16'he565;
        src75 <= 16'h2295;
        src76 <= 16'h8fa9;
        src77 <= 16'hd587;
        src78 <= 16'haaaf;
        src79 <= 16'h5e93;
        src80 <= 16'h73d9;
        src81 <= 16'h9084;
        src82 <= 16'he3ec;
        src83 <= 16'h322;
        src84 <= 16'he46f;
        src85 <= 16'hf59;
        src86 <= 16'hc04c;
        src87 <= 16'h3ef4;
        src88 <= 16'hb564;
        src89 <= 16'h1c3f;
        src90 <= 16'h70aa;
        src91 <= 16'hdca;
        src92 <= 16'h7df1;
        src93 <= 16'h8600;
        src94 <= 16'ha955;
        src95 <= 16'hdd84;
        src96 <= 16'hec5e;
        src97 <= 16'hc792;
        src98 <= 16'hb4db;
        src99 <= 16'h1c08;
        src100 <= 16'hb133;
        src101 <= 16'ha77c;
        src102 <= 16'h4a26;
        src103 <= 16'hb9ce;
        src104 <= 16'ha823;
        src105 <= 16'ha2b4;
        src106 <= 16'hba9d;
        src107 <= 16'h393c;
        src108 <= 16'hd408;
        src109 <= 16'hed04;
        src110 <= 16'hc594;
        src111 <= 16'h6;
        src112 <= 16'hc483;
        src113 <= 16'hba80;
        src114 <= 16'h18b0;
        src115 <= 16'h8d77;
        src116 <= 16'hdadc;
        src117 <= 16'h4c27;
        src118 <= 16'hebdf;
        src119 <= 16'h4e51;
        src120 <= 16'hf507;
        src121 <= 16'h4b24;
        src122 <= 16'h51a6;
        src123 <= 16'h4d6c;
        src124 <= 16'h2272;
        src125 <= 16'hd626;
        src126 <= 16'h4bc6;
        src127 <= 16'h9fb0;
        src128 <= 16'hae9c;
        src129 <= 16'h5e1d;
        src130 <= 16'h1f89;
        src131 <= 16'h2896;
        src132 <= 16'hd56c;
        src133 <= 16'h6279;
        src134 <= 16'haf98;
        src135 <= 16'h2c;
        src136 <= 16'had46;
        src137 <= 16'hd456;
        src138 <= 16'h697;
        src139 <= 16'h61b7;
        src140 <= 16'hc6b2;
        src141 <= 16'hcd6d;
        src142 <= 16'h72bb;
        src143 <= 16'hf364;
        src144 <= 16'h38f5;
        src145 <= 16'h67e3;
        src146 <= 16'ha6c7;
        src147 <= 16'h4b32;
        src148 <= 16'h1c78;
        src149 <= 16'h1d32;
        src150 <= 16'h38e0;
        src151 <= 16'h7aba;
        src152 <= 16'ha99a;
        src153 <= 16'h3fed;
        src154 <= 16'hda1a;
        src155 <= 16'h3651;
        src156 <= 16'h32d0;
        src157 <= 16'h21d6;
        src158 <= 16'h66d;
        src159 <= 16'h0;
        src160 <= 16'h4476;
        src161 <= 16'h2e9e;
        src162 <= 16'h80c8;
        src163 <= 16'hf9c5;
        src164 <= 16'h272d;
        src165 <= 16'h466c;
        src166 <= 16'h9363;
        src167 <= 16'h779b;
        src168 <= 16'ha0c3;
        src169 <= 16'h2500;
        src170 <= 16'h535d;
        src171 <= 16'h1a73;
        src172 <= 16'h333;
        src173 <= 16'h94d6;
        src174 <= 16'hdd87;
        src175 <= 16'he0a9;
        src176 <= 16'hf32d;
        src177 <= 16'hb61e;
        src178 <= 16'h627f;
        src179 <= 16'hcb01;
        src180 <= 16'ha70e;
        src181 <= 16'h4cc0;
        src182 <= 16'h310e;
        src183 <= 16'hab7d;
        src184 <= 16'hc748;
        exp <= 24'h5fd724;
        #1
        src0 <= 16'h4639;
        src1 <= 16'h957b;
        src2 <= 16'hdb6c;
        src3 <= 16'hbd18;
        src4 <= 16'h2988;
        src5 <= 16'h69e8;
        src6 <= 16'h63b7;
        src7 <= 16'h283d;
        src8 <= 16'h6d02;
        src9 <= 16'he9b9;
        src10 <= 16'he7c1;
        src11 <= 16'hc942;
        src12 <= 16'h9a48;
        src13 <= 16'h2828;
        src14 <= 16'haaa9;
        src15 <= 16'hfbda;
        src16 <= 16'hf60f;
        src17 <= 16'hadab;
        src18 <= 16'h98f9;
        src19 <= 16'ha70d;
        src20 <= 16'hbb1d;
        src21 <= 16'h783f;
        src22 <= 16'h3f87;
        src23 <= 16'hcf98;
        src24 <= 16'h597b;
        src25 <= 16'h1a5d;
        src26 <= 16'h6488;
        src27 <= 16'h1efc;
        src28 <= 16'h606a;
        src29 <= 16'h7771;
        src30 <= 16'hc44;
        src31 <= 16'h5d6;
        src32 <= 16'hf20d;
        src33 <= 16'h5c9e;
        src34 <= 16'hf82d;
        src35 <= 16'h74c2;
        src36 <= 16'hed54;
        src37 <= 16'hd228;
        src38 <= 16'h7ec4;
        src39 <= 16'h34e7;
        src40 <= 16'hec8e;
        src41 <= 16'hcfe5;
        src42 <= 16'h34ff;
        src43 <= 16'ha258;
        src44 <= 16'hfc46;
        src45 <= 16'hb491;
        src46 <= 16'h80c1;
        src47 <= 16'h68d5;
        src48 <= 16'hbbdc;
        src49 <= 16'h4742;
        src50 <= 16'hbfa1;
        src51 <= 16'ha0d9;
        src52 <= 16'h676a;
        src53 <= 16'h4b99;
        src54 <= 16'h66c4;
        src55 <= 16'h2a6c;
        src56 <= 16'he978;
        src57 <= 16'h59a7;
        src58 <= 16'hd85b;
        src59 <= 16'hecf5;
        src60 <= 16'hd9e0;
        src61 <= 16'h7150;
        src62 <= 16'heb17;
        src63 <= 16'hef1b;
        src64 <= 16'hdda1;
        src65 <= 16'h6f96;
        src66 <= 16'h796e;
        src67 <= 16'hc8a;
        src68 <= 16'hd8ac;
        src69 <= 16'h5b7b;
        src70 <= 16'hd409;
        src71 <= 16'h2b3b;
        src72 <= 16'h67c;
        src73 <= 16'h9690;
        src74 <= 16'h86fe;
        src75 <= 16'hd753;
        src76 <= 16'h1a4;
        src77 <= 16'h79e5;
        src78 <= 16'h4eab;
        src79 <= 16'h53c0;
        src80 <= 16'h291b;
        src81 <= 16'h22b5;
        src82 <= 16'h4c7f;
        src83 <= 16'h9c3c;
        src84 <= 16'h59dd;
        src85 <= 16'h8ff7;
        src86 <= 16'h1ea9;
        src87 <= 16'hc1a5;
        src88 <= 16'h64c2;
        src89 <= 16'h62c1;
        src90 <= 16'h1019;
        src91 <= 16'h9d47;
        src92 <= 16'hd985;
        src93 <= 16'ha2a7;
        src94 <= 16'h9309;
        src95 <= 16'he996;
        src96 <= 16'h483f;
        src97 <= 16'h750b;
        src98 <= 16'hb925;
        src99 <= 16'hec62;
        src100 <= 16'h3807;
        src101 <= 16'h52c3;
        src102 <= 16'h8ed3;
        src103 <= 16'h3a35;
        src104 <= 16'hc9e1;
        src105 <= 16'h6a51;
        src106 <= 16'h4402;
        src107 <= 16'h42b;
        src108 <= 16'h4d88;
        src109 <= 16'hdf05;
        src110 <= 16'h2eab;
        src111 <= 16'hbbd7;
        src112 <= 16'ha722;
        src113 <= 16'h5d82;
        src114 <= 16'h21cd;
        src115 <= 16'hf367;
        src116 <= 16'h4a9;
        src117 <= 16'h780c;
        src118 <= 16'h335c;
        src119 <= 16'h67e3;
        src120 <= 16'he862;
        src121 <= 16'h1e59;
        src122 <= 16'hd42c;
        src123 <= 16'hd619;
        src124 <= 16'hc31a;
        src125 <= 16'h3dee;
        src126 <= 16'h17b4;
        src127 <= 16'h3dbc;
        src128 <= 16'h9aba;
        src129 <= 16'h59ff;
        src130 <= 16'hec85;
        src131 <= 16'h7235;
        src132 <= 16'h9516;
        src133 <= 16'hbc1e;
        src134 <= 16'h71fc;
        src135 <= 16'hd583;
        src136 <= 16'h8ef3;
        src137 <= 16'h4df1;
        src138 <= 16'h8346;
        src139 <= 16'hf984;
        src140 <= 16'h2ad1;
        src141 <= 16'h502a;
        src142 <= 16'hd5a0;
        src143 <= 16'h27ab;
        src144 <= 16'h815b;
        src145 <= 16'h58e3;
        src146 <= 16'hee1c;
        src147 <= 16'hd17b;
        src148 <= 16'h2b00;
        src149 <= 16'hf935;
        src150 <= 16'h3c0b;
        src151 <= 16'hf7f3;
        src152 <= 16'h71f8;
        src153 <= 16'hdf30;
        src154 <= 16'h7fbe;
        src155 <= 16'h75e7;
        src156 <= 16'h8593;
        src157 <= 16'h279d;
        src158 <= 16'h7e01;
        src159 <= 16'h984d;
        src160 <= 16'h2f0e;
        src161 <= 16'hc013;
        src162 <= 16'h21f8;
        src163 <= 16'h275;
        src164 <= 16'hf739;
        src165 <= 16'h3a5e;
        src166 <= 16'h657d;
        src167 <= 16'h46;
        src168 <= 16'hfa97;
        src169 <= 16'hc1f2;
        src170 <= 16'h2e84;
        src171 <= 16'had1b;
        src172 <= 16'h57e8;
        src173 <= 16'h483b;
        src174 <= 16'h5c9c;
        src175 <= 16'h3760;
        src176 <= 16'h4af0;
        src177 <= 16'h9ade;
        src178 <= 16'hfe7c;
        src179 <= 16'hed62;
        src180 <= 16'h19e2;
        src181 <= 16'hbfd2;
        src182 <= 16'he23a;
        src183 <= 16'h259;
        src184 <= 16'h3432;
        exp <= 24'h5e43c9;
        #1
        src0 <= 16'hf66;
        src1 <= 16'h270b;
        src2 <= 16'h5e64;
        src3 <= 16'h335e;
        src4 <= 16'h6036;
        src5 <= 16'h45ed;
        src6 <= 16'hd7b0;
        src7 <= 16'h823c;
        src8 <= 16'h4a90;
        src9 <= 16'h6700;
        src10 <= 16'hc6a0;
        src11 <= 16'he4;
        src12 <= 16'h2ce4;
        src13 <= 16'h9933;
        src14 <= 16'hb5b0;
        src15 <= 16'he4a5;
        src16 <= 16'heef7;
        src17 <= 16'he425;
        src18 <= 16'h71ad;
        src19 <= 16'hf24;
        src20 <= 16'h6250;
        src21 <= 16'h12b2;
        src22 <= 16'h6f68;
        src23 <= 16'hf2ae;
        src24 <= 16'h4257;
        src25 <= 16'hdb1c;
        src26 <= 16'h5a98;
        src27 <= 16'hbb26;
        src28 <= 16'h50e4;
        src29 <= 16'h888d;
        src30 <= 16'h7496;
        src31 <= 16'hd621;
        src32 <= 16'hcf92;
        src33 <= 16'hd8c1;
        src34 <= 16'h2c2b;
        src35 <= 16'hc98f;
        src36 <= 16'h6833;
        src37 <= 16'h60f1;
        src38 <= 16'hbd15;
        src39 <= 16'h55bc;
        src40 <= 16'h52fe;
        src41 <= 16'hde;
        src42 <= 16'ha743;
        src43 <= 16'h97f5;
        src44 <= 16'h1289;
        src45 <= 16'h5fa;
        src46 <= 16'h7085;
        src47 <= 16'h3fb2;
        src48 <= 16'h8081;
        src49 <= 16'h3e74;
        src50 <= 16'ha46;
        src51 <= 16'he6fc;
        src52 <= 16'h9fc9;
        src53 <= 16'hfb80;
        src54 <= 16'hb640;
        src55 <= 16'ha1ea;
        src56 <= 16'h33e;
        src57 <= 16'h7269;
        src58 <= 16'h9df3;
        src59 <= 16'h67b3;
        src60 <= 16'hc9b;
        src61 <= 16'h593a;
        src62 <= 16'h9b60;
        src63 <= 16'hbc9b;
        src64 <= 16'h4bbc;
        src65 <= 16'h4edb;
        src66 <= 16'h7232;
        src67 <= 16'hbe4b;
        src68 <= 16'h154;
        src69 <= 16'h2d51;
        src70 <= 16'hc741;
        src71 <= 16'h443e;
        src72 <= 16'h9bf8;
        src73 <= 16'hcaec;
        src74 <= 16'h62b0;
        src75 <= 16'h4056;
        src76 <= 16'hc209;
        src77 <= 16'hddf7;
        src78 <= 16'hab53;
        src79 <= 16'h8deb;
        src80 <= 16'hfe14;
        src81 <= 16'h1c6f;
        src82 <= 16'haf98;
        src83 <= 16'h745c;
        src84 <= 16'h5ca4;
        src85 <= 16'h87af;
        src86 <= 16'h1268;
        src87 <= 16'he566;
        src88 <= 16'ha7d6;
        src89 <= 16'hc14b;
        src90 <= 16'h1584;
        src91 <= 16'h5586;
        src92 <= 16'h1870;
        src93 <= 16'hbe82;
        src94 <= 16'h9627;
        src95 <= 16'h6a77;
        src96 <= 16'h8eda;
        src97 <= 16'hfd7b;
        src98 <= 16'hcf5d;
        src99 <= 16'hca29;
        src100 <= 16'h7af3;
        src101 <= 16'h5c8;
        src102 <= 16'hce3c;
        src103 <= 16'h96c3;
        src104 <= 16'hd8ec;
        src105 <= 16'h7412;
        src106 <= 16'h5e78;
        src107 <= 16'h92bd;
        src108 <= 16'h1949;
        src109 <= 16'hefe8;
        src110 <= 16'hcef9;
        src111 <= 16'he8d9;
        src112 <= 16'h1df5;
        src113 <= 16'h38f4;
        src114 <= 16'ha967;
        src115 <= 16'h68a;
        src116 <= 16'h6443;
        src117 <= 16'h4f2f;
        src118 <= 16'hee0c;
        src119 <= 16'h6edd;
        src120 <= 16'hccee;
        src121 <= 16'h91d4;
        src122 <= 16'h937;
        src123 <= 16'h930e;
        src124 <= 16'hd605;
        src125 <= 16'he917;
        src126 <= 16'h3b0f;
        src127 <= 16'hd5fa;
        src128 <= 16'hfa93;
        src129 <= 16'h8df9;
        src130 <= 16'h9ae7;
        src131 <= 16'h7087;
        src132 <= 16'ha266;
        src133 <= 16'h1092;
        src134 <= 16'h826a;
        src135 <= 16'hbd27;
        src136 <= 16'ha477;
        src137 <= 16'h21a4;
        src138 <= 16'h877e;
        src139 <= 16'h4263;
        src140 <= 16'h4;
        src141 <= 16'hc0c1;
        src142 <= 16'h9826;
        src143 <= 16'h4d90;
        src144 <= 16'ha5b8;
        src145 <= 16'ha85;
        src146 <= 16'h92bf;
        src147 <= 16'h9068;
        src148 <= 16'h2ab0;
        src149 <= 16'h1428;
        src150 <= 16'hb353;
        src151 <= 16'hc259;
        src152 <= 16'h5a32;
        src153 <= 16'h5918;
        src154 <= 16'ha5d8;
        src155 <= 16'h1cf6;
        src156 <= 16'ha728;
        src157 <= 16'hb4ad;
        src158 <= 16'h5b22;
        src159 <= 16'hffa9;
        src160 <= 16'ha747;
        src161 <= 16'hc4cf;
        src162 <= 16'h6e70;
        src163 <= 16'hbcbc;
        src164 <= 16'h7fa6;
        src165 <= 16'hbf40;
        src166 <= 16'h444a;
        src167 <= 16'ha594;
        src168 <= 16'h7a45;
        src169 <= 16'h6d33;
        src170 <= 16'h3442;
        src171 <= 16'h48fb;
        src172 <= 16'h530;
        src173 <= 16'hae66;
        src174 <= 16'h493a;
        src175 <= 16'h7f15;
        src176 <= 16'h7923;
        src177 <= 16'h3651;
        src178 <= 16'h11d;
        src179 <= 16'h75d8;
        src180 <= 16'h8384;
        src181 <= 16'h60fa;
        src182 <= 16'h7514;
        src183 <= 16'h866d;
        src184 <= 16'h79d6;
        exp <= 24'h5a050e;
        #1
        src0 <= 16'h3ef6;
        src1 <= 16'hf1be;
        src2 <= 16'hd751;
        src3 <= 16'h22d6;
        src4 <= 16'h4eff;
        src5 <= 16'haef7;
        src6 <= 16'h11f6;
        src7 <= 16'h207c;
        src8 <= 16'hf46e;
        src9 <= 16'hfb6c;
        src10 <= 16'hb6c9;
        src11 <= 16'h9a46;
        src12 <= 16'hc26;
        src13 <= 16'h721a;
        src14 <= 16'he2df;
        src15 <= 16'h82f6;
        src16 <= 16'h75cb;
        src17 <= 16'hf8a0;
        src18 <= 16'h257b;
        src19 <= 16'he69f;
        src20 <= 16'ha1a2;
        src21 <= 16'h790c;
        src22 <= 16'h7cb2;
        src23 <= 16'h9242;
        src24 <= 16'hf99d;
        src25 <= 16'ha596;
        src26 <= 16'hb069;
        src27 <= 16'h1aef;
        src28 <= 16'hb074;
        src29 <= 16'h9429;
        src30 <= 16'hd945;
        src31 <= 16'hbc36;
        src32 <= 16'hfc23;
        src33 <= 16'hf760;
        src34 <= 16'h820b;
        src35 <= 16'h5de6;
        src36 <= 16'h5dfc;
        src37 <= 16'h236c;
        src38 <= 16'h6ac2;
        src39 <= 16'h5959;
        src40 <= 16'h219;
        src41 <= 16'h64d5;
        src42 <= 16'h5da;
        src43 <= 16'h1845;
        src44 <= 16'hb381;
        src45 <= 16'hdd1f;
        src46 <= 16'hc31;
        src47 <= 16'h7bbe;
        src48 <= 16'hd0ad;
        src49 <= 16'hd427;
        src50 <= 16'h3325;
        src51 <= 16'hafe5;
        src52 <= 16'ha449;
        src53 <= 16'hd727;
        src54 <= 16'hdc20;
        src55 <= 16'h2d95;
        src56 <= 16'hed9;
        src57 <= 16'h6403;
        src58 <= 16'hd4b3;
        src59 <= 16'hf742;
        src60 <= 16'hde1e;
        src61 <= 16'h74f8;
        src62 <= 16'h4859;
        src63 <= 16'h7e53;
        src64 <= 16'h6b70;
        src65 <= 16'hc70c;
        src66 <= 16'hafc9;
        src67 <= 16'h2296;
        src68 <= 16'hea5e;
        src69 <= 16'h1d20;
        src70 <= 16'h3693;
        src71 <= 16'h4f5c;
        src72 <= 16'ha8d3;
        src73 <= 16'hf027;
        src74 <= 16'hebdf;
        src75 <= 16'hfe82;
        src76 <= 16'h712b;
        src77 <= 16'h5841;
        src78 <= 16'h6d9b;
        src79 <= 16'hcc72;
        src80 <= 16'h172d;
        src81 <= 16'hcdf4;
        src82 <= 16'h6b34;
        src83 <= 16'h42d5;
        src84 <= 16'hfccb;
        src85 <= 16'h41bd;
        src86 <= 16'hf032;
        src87 <= 16'h98c3;
        src88 <= 16'ha58f;
        src89 <= 16'hd25d;
        src90 <= 16'hfb6;
        src91 <= 16'h7d13;
        src92 <= 16'h16ab;
        src93 <= 16'h1c7f;
        src94 <= 16'hfd7;
        src95 <= 16'h865a;
        src96 <= 16'h74ef;
        src97 <= 16'haff4;
        src98 <= 16'h33ed;
        src99 <= 16'h5270;
        src100 <= 16'had33;
        src101 <= 16'h8bf4;
        src102 <= 16'hf5b9;
        src103 <= 16'h7ffb;
        src104 <= 16'h34ab;
        src105 <= 16'hfa2d;
        src106 <= 16'hca54;
        src107 <= 16'h6e41;
        src108 <= 16'hce08;
        src109 <= 16'h33cd;
        src110 <= 16'hb7eb;
        src111 <= 16'h69f0;
        src112 <= 16'h1f5;
        src113 <= 16'ha7f1;
        src114 <= 16'hfefc;
        src115 <= 16'h52d3;
        src116 <= 16'h885c;
        src117 <= 16'h181;
        src118 <= 16'h9d76;
        src119 <= 16'hb263;
        src120 <= 16'hb90a;
        src121 <= 16'h61d7;
        src122 <= 16'h2f9b;
        src123 <= 16'h6488;
        src124 <= 16'hd820;
        src125 <= 16'hfab8;
        src126 <= 16'h4e37;
        src127 <= 16'h6cb1;
        src128 <= 16'h1aaf;
        src129 <= 16'h36e7;
        src130 <= 16'h4f93;
        src131 <= 16'h923d;
        src132 <= 16'h4b24;
        src133 <= 16'hefab;
        src134 <= 16'h160c;
        src135 <= 16'h4b6e;
        src136 <= 16'h14fb;
        src137 <= 16'h587c;
        src138 <= 16'hb0a9;
        src139 <= 16'hf90b;
        src140 <= 16'h2893;
        src141 <= 16'ha67c;
        src142 <= 16'h52b5;
        src143 <= 16'h74c;
        src144 <= 16'hbda3;
        src145 <= 16'hea63;
        src146 <= 16'h11d7;
        src147 <= 16'hc77f;
        src148 <= 16'hf1a;
        src149 <= 16'h93e8;
        src150 <= 16'h9a76;
        src151 <= 16'h8fd1;
        src152 <= 16'hec7c;
        src153 <= 16'h7130;
        src154 <= 16'he582;
        src155 <= 16'hb146;
        src156 <= 16'hdaac;
        src157 <= 16'hdddf;
        src158 <= 16'h2235;
        src159 <= 16'he9ac;
        src160 <= 16'h407f;
        src161 <= 16'h7eb;
        src162 <= 16'h7386;
        src163 <= 16'hd7c6;
        src164 <= 16'h35ea;
        src165 <= 16'hf30b;
        src166 <= 16'h37b4;
        src167 <= 16'hf077;
        src168 <= 16'h779;
        src169 <= 16'h23f3;
        src170 <= 16'h39a8;
        src171 <= 16'hd05a;
        src172 <= 16'h2eb7;
        src173 <= 16'h8773;
        src174 <= 16'ha626;
        src175 <= 16'h72f9;
        src176 <= 16'hcd48;
        src177 <= 16'h21d2;
        src178 <= 16'h2f39;
        src179 <= 16'h29f2;
        src180 <= 16'h3cb;
        src181 <= 16'hc461;
        src182 <= 16'h5bd1;
        src183 <= 16'h575c;
        src184 <= 16'h455f;
        exp <= 24'h5dc867;
        #1
        src0 <= 16'h1615;
        src1 <= 16'h5ffb;
        src2 <= 16'ha1e;
        src3 <= 16'haa75;
        src4 <= 16'h8d8c;
        src5 <= 16'h936a;
        src6 <= 16'h7de7;
        src7 <= 16'h1059;
        src8 <= 16'hd8a6;
        src9 <= 16'h1001;
        src10 <= 16'h4d4e;
        src11 <= 16'hc5c2;
        src12 <= 16'h6396;
        src13 <= 16'h4d75;
        src14 <= 16'h7e4e;
        src15 <= 16'hd0eb;
        src16 <= 16'h38b6;
        src17 <= 16'h2276;
        src18 <= 16'h895c;
        src19 <= 16'hb43e;
        src20 <= 16'hbbaa;
        src21 <= 16'h27f0;
        src22 <= 16'h9734;
        src23 <= 16'hfb77;
        src24 <= 16'h9a9f;
        src25 <= 16'h5560;
        src26 <= 16'hd2e9;
        src27 <= 16'h7878;
        src28 <= 16'h8fbe;
        src29 <= 16'hfcb7;
        src30 <= 16'h7e89;
        src31 <= 16'h3731;
        src32 <= 16'h72b9;
        src33 <= 16'h8207;
        src34 <= 16'h4745;
        src35 <= 16'he4f5;
        src36 <= 16'h3560;
        src37 <= 16'h63bf;
        src38 <= 16'h9b9c;
        src39 <= 16'hb71c;
        src40 <= 16'hfe3;
        src41 <= 16'h939f;
        src42 <= 16'h95a7;
        src43 <= 16'h8e4f;
        src44 <= 16'h8545;
        src45 <= 16'h1a12;
        src46 <= 16'h332f;
        src47 <= 16'h6ac5;
        src48 <= 16'he767;
        src49 <= 16'he317;
        src50 <= 16'h4698;
        src51 <= 16'hde81;
        src52 <= 16'h671b;
        src53 <= 16'h699f;
        src54 <= 16'ha2bd;
        src55 <= 16'h724d;
        src56 <= 16'ha32f;
        src57 <= 16'h1be9;
        src58 <= 16'hed5d;
        src59 <= 16'hae0d;
        src60 <= 16'hbf00;
        src61 <= 16'h53ed;
        src62 <= 16'hcdbb;
        src63 <= 16'hfcf;
        src64 <= 16'he795;
        src65 <= 16'h8572;
        src66 <= 16'hdf20;
        src67 <= 16'ha07a;
        src68 <= 16'h1068;
        src69 <= 16'h4c13;
        src70 <= 16'ha1d3;
        src71 <= 16'h7bd4;
        src72 <= 16'h6a30;
        src73 <= 16'h1f7b;
        src74 <= 16'h20fd;
        src75 <= 16'h2646;
        src76 <= 16'h5640;
        src77 <= 16'h7b1;
        src78 <= 16'h3b3d;
        src79 <= 16'hc8bc;
        src80 <= 16'h920a;
        src81 <= 16'h8ecf;
        src82 <= 16'h890a;
        src83 <= 16'hb8c;
        src84 <= 16'h1637;
        src85 <= 16'hfad7;
        src86 <= 16'hd0e7;
        src87 <= 16'ha0f9;
        src88 <= 16'he63d;
        src89 <= 16'hb56f;
        src90 <= 16'h8da3;
        src91 <= 16'h9362;
        src92 <= 16'h8540;
        src93 <= 16'ha39e;
        src94 <= 16'hadb8;
        src95 <= 16'hc73d;
        src96 <= 16'h32a0;
        src97 <= 16'hf2cc;
        src98 <= 16'h500a;
        src99 <= 16'h68b3;
        src100 <= 16'hf21e;
        src101 <= 16'h724f;
        src102 <= 16'hdf8e;
        src103 <= 16'h20a5;
        src104 <= 16'hd163;
        src105 <= 16'hbb41;
        src106 <= 16'h1d8b;
        src107 <= 16'h79c5;
        src108 <= 16'h6170;
        src109 <= 16'hd8c9;
        src110 <= 16'h4fd0;
        src111 <= 16'h4696;
        src112 <= 16'h43e9;
        src113 <= 16'h6834;
        src114 <= 16'h7735;
        src115 <= 16'h559f;
        src116 <= 16'h90aa;
        src117 <= 16'hc21;
        src118 <= 16'h789f;
        src119 <= 16'hacf4;
        src120 <= 16'hc8a7;
        src121 <= 16'hfa9;
        src122 <= 16'h624d;
        src123 <= 16'h2d77;
        src124 <= 16'hcb5d;
        src125 <= 16'h7706;
        src126 <= 16'he3fb;
        src127 <= 16'h5c6d;
        src128 <= 16'hf273;
        src129 <= 16'h5ee4;
        src130 <= 16'hd379;
        src131 <= 16'h5bbe;
        src132 <= 16'h3603;
        src133 <= 16'h662b;
        src134 <= 16'hcf5e;
        src135 <= 16'h6acb;
        src136 <= 16'h9ed0;
        src137 <= 16'h3baf;
        src138 <= 16'h7c1b;
        src139 <= 16'h1e81;
        src140 <= 16'hc231;
        src141 <= 16'hc680;
        src142 <= 16'h847c;
        src143 <= 16'h238f;
        src144 <= 16'h4875;
        src145 <= 16'h16b3;
        src146 <= 16'hc857;
        src147 <= 16'hb21d;
        src148 <= 16'ha718;
        src149 <= 16'h7c46;
        src150 <= 16'h6d3b;
        src151 <= 16'h8658;
        src152 <= 16'h73a3;
        src153 <= 16'h7e6c;
        src154 <= 16'h466d;
        src155 <= 16'hc546;
        src156 <= 16'h57fe;
        src157 <= 16'h5c63;
        src158 <= 16'he6fa;
        src159 <= 16'h5fcb;
        src160 <= 16'hc8fe;
        src161 <= 16'h52b3;
        src162 <= 16'h97f;
        src163 <= 16'hff35;
        src164 <= 16'h2b23;
        src165 <= 16'h8546;
        src166 <= 16'h222a;
        src167 <= 16'h1aff;
        src168 <= 16'haeb9;
        src169 <= 16'he21;
        src170 <= 16'h2a25;
        src171 <= 16'h62b7;
        src172 <= 16'hb74c;
        src173 <= 16'h129f;
        src174 <= 16'h41c0;
        src175 <= 16'hb139;
        src176 <= 16'h6cdd;
        src177 <= 16'h9016;
        src178 <= 16'h8ca2;
        src179 <= 16'h522d;
        src180 <= 16'h4a1e;
        src181 <= 16'hf52f;
        src182 <= 16'haaef;
        src183 <= 16'h246b;
        src184 <= 16'had29;
        exp <= 24'h59b4b0;
        #1
        src0 <= 16'h7495;
        src1 <= 16'hb50a;
        src2 <= 16'hb94a;
        src3 <= 16'he59f;
        src4 <= 16'h1e76;
        src5 <= 16'h440a;
        src6 <= 16'h577c;
        src7 <= 16'h41a3;
        src8 <= 16'hbe72;
        src9 <= 16'hf42d;
        src10 <= 16'h4419;
        src11 <= 16'hc82;
        src12 <= 16'hd17e;
        src13 <= 16'h1c2d;
        src14 <= 16'h6111;
        src15 <= 16'h4e0b;
        src16 <= 16'h634;
        src17 <= 16'hd451;
        src18 <= 16'h850a;
        src19 <= 16'h25fb;
        src20 <= 16'hb6ea;
        src21 <= 16'hdf5c;
        src22 <= 16'h56f2;
        src23 <= 16'ha978;
        src24 <= 16'h5c36;
        src25 <= 16'hc924;
        src26 <= 16'hfeae;
        src27 <= 16'h175;
        src28 <= 16'hcd38;
        src29 <= 16'h606d;
        src30 <= 16'h7f52;
        src31 <= 16'h5691;
        src32 <= 16'he55b;
        src33 <= 16'h4e9;
        src34 <= 16'hf43b;
        src35 <= 16'h6318;
        src36 <= 16'h28ae;
        src37 <= 16'hd8b9;
        src38 <= 16'h46e1;
        src39 <= 16'h5e03;
        src40 <= 16'h4c65;
        src41 <= 16'hc93f;
        src42 <= 16'h1eac;
        src43 <= 16'h2006;
        src44 <= 16'ha129;
        src45 <= 16'ha5de;
        src46 <= 16'h1f30;
        src47 <= 16'h694e;
        src48 <= 16'h2021;
        src49 <= 16'h61;
        src50 <= 16'he991;
        src51 <= 16'hb8e2;
        src52 <= 16'ha09c;
        src53 <= 16'h60ad;
        src54 <= 16'h6aa7;
        src55 <= 16'h6f02;
        src56 <= 16'h6015;
        src57 <= 16'h3a5c;
        src58 <= 16'h2c4a;
        src59 <= 16'h2a04;
        src60 <= 16'hcc67;
        src61 <= 16'hce71;
        src62 <= 16'hea09;
        src63 <= 16'he60b;
        src64 <= 16'hab2e;
        src65 <= 16'h7ba3;
        src66 <= 16'h517e;
        src67 <= 16'h2d14;
        src68 <= 16'h56a6;
        src69 <= 16'h517e;
        src70 <= 16'hbb50;
        src71 <= 16'hb9c;
        src72 <= 16'hf57e;
        src73 <= 16'h9c63;
        src74 <= 16'hb8a5;
        src75 <= 16'h5c44;
        src76 <= 16'h5f61;
        src77 <= 16'h5fb3;
        src78 <= 16'h291f;
        src79 <= 16'hf539;
        src80 <= 16'haac;
        src81 <= 16'h2c4a;
        src82 <= 16'hc2b;
        src83 <= 16'h800c;
        src84 <= 16'hdf92;
        src85 <= 16'hbe63;
        src86 <= 16'he051;
        src87 <= 16'h8991;
        src88 <= 16'h1479;
        src89 <= 16'hf907;
        src90 <= 16'h4c90;
        src91 <= 16'h99ae;
        src92 <= 16'h9701;
        src93 <= 16'h30a5;
        src94 <= 16'h5ea9;
        src95 <= 16'hfcc6;
        src96 <= 16'h5094;
        src97 <= 16'h9dcf;
        src98 <= 16'h3aea;
        src99 <= 16'h2e09;
        src100 <= 16'hf66e;
        src101 <= 16'h9295;
        src102 <= 16'h42a7;
        src103 <= 16'hae0f;
        src104 <= 16'hb7d;
        src105 <= 16'h4ea1;
        src106 <= 16'h6087;
        src107 <= 16'ha345;
        src108 <= 16'h9ba8;
        src109 <= 16'h9957;
        src110 <= 16'h2b1f;
        src111 <= 16'hef2c;
        src112 <= 16'h2782;
        src113 <= 16'hd684;
        src114 <= 16'hec7c;
        src115 <= 16'h4e75;
        src116 <= 16'h568a;
        src117 <= 16'h84d6;
        src118 <= 16'h2426;
        src119 <= 16'h855c;
        src120 <= 16'he7d4;
        src121 <= 16'h15ad;
        src122 <= 16'he983;
        src123 <= 16'h17bf;
        src124 <= 16'h2a7c;
        src125 <= 16'h4e8f;
        src126 <= 16'hf142;
        src127 <= 16'h7ae3;
        src128 <= 16'h49f1;
        src129 <= 16'h4a73;
        src130 <= 16'h20da;
        src131 <= 16'hc7df;
        src132 <= 16'h7d55;
        src133 <= 16'h42da;
        src134 <= 16'he3d3;
        src135 <= 16'h1ea3;
        src136 <= 16'h349b;
        src137 <= 16'h42a;
        src138 <= 16'h999a;
        src139 <= 16'hc0;
        src140 <= 16'h8b56;
        src141 <= 16'hdc17;
        src142 <= 16'hd296;
        src143 <= 16'h97d4;
        src144 <= 16'hc482;
        src145 <= 16'had8f;
        src146 <= 16'h6bf2;
        src147 <= 16'hf8d;
        src148 <= 16'h88e;
        src149 <= 16'hd3d6;
        src150 <= 16'hb9a5;
        src151 <= 16'h43dc;
        src152 <= 16'h946d;
        src153 <= 16'h5d1a;
        src154 <= 16'h5b9e;
        src155 <= 16'h8628;
        src156 <= 16'h99ea;
        src157 <= 16'h22f7;
        src158 <= 16'h822a;
        src159 <= 16'ha746;
        src160 <= 16'h486d;
        src161 <= 16'h2c8d;
        src162 <= 16'h44dd;
        src163 <= 16'h11dc;
        src164 <= 16'h5e54;
        src165 <= 16'h5061;
        src166 <= 16'h4408;
        src167 <= 16'h746e;
        src168 <= 16'h95d6;
        src169 <= 16'h4077;
        src170 <= 16'h33fc;
        src171 <= 16'h2a06;
        src172 <= 16'h8c4e;
        src173 <= 16'haf3a;
        src174 <= 16'h343;
        src175 <= 16'hf1e2;
        src176 <= 16'h5105;
        src177 <= 16'h6a8e;
        src178 <= 16'h2898;
        src179 <= 16'hb46a;
        src180 <= 16'h17a1;
        src181 <= 16'hc690;
        src182 <= 16'h9e87;
        src183 <= 16'hf798;
        src184 <= 16'h811;
        exp <= 24'h555be0;
        #1
        src0 <= 16'hcb8e;
        src1 <= 16'head;
        src2 <= 16'hb35f;
        src3 <= 16'h6899;
        src4 <= 16'h1b8b;
        src5 <= 16'hd919;
        src6 <= 16'h3d52;
        src7 <= 16'hf69b;
        src8 <= 16'h4181;
        src9 <= 16'h5fa4;
        src10 <= 16'he192;
        src11 <= 16'h4738;
        src12 <= 16'h4dd0;
        src13 <= 16'h890b;
        src14 <= 16'h1534;
        src15 <= 16'hc287;
        src16 <= 16'hc3a1;
        src17 <= 16'h3996;
        src18 <= 16'hc728;
        src19 <= 16'h614c;
        src20 <= 16'h5a5a;
        src21 <= 16'he65d;
        src22 <= 16'h3540;
        src23 <= 16'hbc36;
        src24 <= 16'h4328;
        src25 <= 16'hcf35;
        src26 <= 16'h60b5;
        src27 <= 16'h6afb;
        src28 <= 16'hca15;
        src29 <= 16'h9a2b;
        src30 <= 16'h426f;
        src31 <= 16'hb79a;
        src32 <= 16'he460;
        src33 <= 16'hbf81;
        src34 <= 16'hec21;
        src35 <= 16'hb13c;
        src36 <= 16'heab0;
        src37 <= 16'hbbd6;
        src38 <= 16'hb3bd;
        src39 <= 16'h77e1;
        src40 <= 16'haf81;
        src41 <= 16'h213a;
        src42 <= 16'h37ca;
        src43 <= 16'ha55a;
        src44 <= 16'h1469;
        src45 <= 16'h5241;
        src46 <= 16'h76ed;
        src47 <= 16'hcdc4;
        src48 <= 16'h9002;
        src49 <= 16'hf808;
        src50 <= 16'h3684;
        src51 <= 16'h1524;
        src52 <= 16'he372;
        src53 <= 16'h551d;
        src54 <= 16'h1673;
        src55 <= 16'h7812;
        src56 <= 16'he02b;
        src57 <= 16'hd874;
        src58 <= 16'h575c;
        src59 <= 16'hbc82;
        src60 <= 16'h3b5e;
        src61 <= 16'hb0;
        src62 <= 16'h7280;
        src63 <= 16'h4d9e;
        src64 <= 16'h23de;
        src65 <= 16'h28d5;
        src66 <= 16'hab6c;
        src67 <= 16'hfd9;
        src68 <= 16'hfcb4;
        src69 <= 16'h221;
        src70 <= 16'hb1b7;
        src71 <= 16'h376a;
        src72 <= 16'ha17f;
        src73 <= 16'h2983;
        src74 <= 16'hbbc;
        src75 <= 16'hc55;
        src76 <= 16'hb13d;
        src77 <= 16'ha98f;
        src78 <= 16'h32cc;
        src79 <= 16'hab72;
        src80 <= 16'ha167;
        src81 <= 16'h3ba;
        src82 <= 16'h39f5;
        src83 <= 16'hc8b9;
        src84 <= 16'h219d;
        src85 <= 16'h99ff;
        src86 <= 16'h87bf;
        src87 <= 16'h80b6;
        src88 <= 16'h52e8;
        src89 <= 16'h5736;
        src90 <= 16'hcbd5;
        src91 <= 16'h2660;
        src92 <= 16'hf824;
        src93 <= 16'h1038;
        src94 <= 16'hac7e;
        src95 <= 16'hd2e7;
        src96 <= 16'hff88;
        src97 <= 16'h800c;
        src98 <= 16'h931b;
        src99 <= 16'h2645;
        src100 <= 16'h6044;
        src101 <= 16'h8881;
        src102 <= 16'h7d35;
        src103 <= 16'haa8d;
        src104 <= 16'h2c1b;
        src105 <= 16'h471c;
        src106 <= 16'h125c;
        src107 <= 16'heacb;
        src108 <= 16'h71d0;
        src109 <= 16'h76a7;
        src110 <= 16'h9f94;
        src111 <= 16'h76b2;
        src112 <= 16'hdc1b;
        src113 <= 16'he761;
        src114 <= 16'h646;
        src115 <= 16'hfba5;
        src116 <= 16'h30d5;
        src117 <= 16'haba0;
        src118 <= 16'h9895;
        src119 <= 16'h2999;
        src120 <= 16'hb796;
        src121 <= 16'h28b;
        src122 <= 16'h6e96;
        src123 <= 16'h8e3a;
        src124 <= 16'h56e;
        src125 <= 16'hd7a4;
        src126 <= 16'h2096;
        src127 <= 16'h4b32;
        src128 <= 16'he4f7;
        src129 <= 16'h6026;
        src130 <= 16'ha80c;
        src131 <= 16'hd40d;
        src132 <= 16'hfc71;
        src133 <= 16'ha1a;
        src134 <= 16'h7e46;
        src135 <= 16'hd90b;
        src136 <= 16'h8b72;
        src137 <= 16'h83ec;
        src138 <= 16'he0e4;
        src139 <= 16'h62c6;
        src140 <= 16'hb935;
        src141 <= 16'h2ee5;
        src142 <= 16'hf309;
        src143 <= 16'hf86;
        src144 <= 16'h724c;
        src145 <= 16'h2176;
        src146 <= 16'h7e8e;
        src147 <= 16'h8487;
        src148 <= 16'h8662;
        src149 <= 16'h5047;
        src150 <= 16'h47c1;
        src151 <= 16'h79fa;
        src152 <= 16'h7256;
        src153 <= 16'heea4;
        src154 <= 16'h196e;
        src155 <= 16'hd2ac;
        src156 <= 16'h30b8;
        src157 <= 16'h2471;
        src158 <= 16'h235d;
        src159 <= 16'h5e4b;
        src160 <= 16'h38b6;
        src161 <= 16'h9f66;
        src162 <= 16'h476a;
        src163 <= 16'he605;
        src164 <= 16'haa0d;
        src165 <= 16'hf5dd;
        src166 <= 16'h8a58;
        src167 <= 16'h32c7;
        src168 <= 16'h7ad8;
        src169 <= 16'hc1e3;
        src170 <= 16'h2f30;
        src171 <= 16'hf6b4;
        src172 <= 16'h2678;
        src173 <= 16'h2da6;
        src174 <= 16'h7fda;
        src175 <= 16'h8ba8;
        src176 <= 16'h51f9;
        src177 <= 16'he218;
        src178 <= 16'hd24e;
        src179 <= 16'hc337;
        src180 <= 16'h75a;
        src181 <= 16'ha175;
        src182 <= 16'hc4a4;
        src183 <= 16'hb021;
        src184 <= 16'h2838;
        exp <= 24'h5a9804;
        #1
        src0 <= 16'h471e;
        src1 <= 16'h89dc;
        src2 <= 16'h2224;
        src3 <= 16'hba37;
        src4 <= 16'h38c4;
        src5 <= 16'h7a2f;
        src6 <= 16'h897f;
        src7 <= 16'haa13;
        src8 <= 16'h28c0;
        src9 <= 16'h25fb;
        src10 <= 16'h1424;
        src11 <= 16'h5a58;
        src12 <= 16'h6260;
        src13 <= 16'he924;
        src14 <= 16'h2cc9;
        src15 <= 16'hef4b;
        src16 <= 16'h245a;
        src17 <= 16'he4;
        src18 <= 16'h9079;
        src19 <= 16'hd09;
        src20 <= 16'h51a1;
        src21 <= 16'h72d7;
        src22 <= 16'h17bd;
        src23 <= 16'hf680;
        src24 <= 16'h9513;
        src25 <= 16'hc3ab;
        src26 <= 16'hcd98;
        src27 <= 16'ha160;
        src28 <= 16'hefc1;
        src29 <= 16'hee1f;
        src30 <= 16'h7;
        src31 <= 16'h215f;
        src32 <= 16'h3044;
        src33 <= 16'he495;
        src34 <= 16'h1b3f;
        src35 <= 16'ha7e2;
        src36 <= 16'hea02;
        src37 <= 16'hd0ac;
        src38 <= 16'hfdb9;
        src39 <= 16'hec5e;
        src40 <= 16'h11e6;
        src41 <= 16'h433f;
        src42 <= 16'hc651;
        src43 <= 16'hc108;
        src44 <= 16'h4d7f;
        src45 <= 16'h4938;
        src46 <= 16'h8f77;
        src47 <= 16'h801b;
        src48 <= 16'h8deb;
        src49 <= 16'hb09b;
        src50 <= 16'hcda9;
        src51 <= 16'h4966;
        src52 <= 16'ha89f;
        src53 <= 16'h32c8;
        src54 <= 16'h7588;
        src55 <= 16'heaba;
        src56 <= 16'h949f;
        src57 <= 16'he196;
        src58 <= 16'h2eca;
        src59 <= 16'hceb6;
        src60 <= 16'h6a9a;
        src61 <= 16'hf8f9;
        src62 <= 16'ha9b5;
        src63 <= 16'h6fbf;
        src64 <= 16'hc98c;
        src65 <= 16'h31e1;
        src66 <= 16'hf18f;
        src67 <= 16'ha279;
        src68 <= 16'h8ff1;
        src69 <= 16'h3485;
        src70 <= 16'hf63f;
        src71 <= 16'h26ca;
        src72 <= 16'he152;
        src73 <= 16'h16ed;
        src74 <= 16'ha58a;
        src75 <= 16'hee31;
        src76 <= 16'hdbf9;
        src77 <= 16'hd1d;
        src78 <= 16'h9322;
        src79 <= 16'he313;
        src80 <= 16'h538b;
        src81 <= 16'h677e;
        src82 <= 16'h26a9;
        src83 <= 16'hf7fb;
        src84 <= 16'hae0d;
        src85 <= 16'h47ea;
        src86 <= 16'h3083;
        src87 <= 16'hb9a8;
        src88 <= 16'h24a1;
        src89 <= 16'h85a4;
        src90 <= 16'hc549;
        src91 <= 16'h4222;
        src92 <= 16'h61dd;
        src93 <= 16'h5b53;
        src94 <= 16'h4625;
        src95 <= 16'h5ed8;
        src96 <= 16'h7abd;
        src97 <= 16'h53f7;
        src98 <= 16'h498;
        src99 <= 16'h5f41;
        src100 <= 16'hbb;
        src101 <= 16'h4386;
        src102 <= 16'h796e;
        src103 <= 16'h78f8;
        src104 <= 16'h19f2;
        src105 <= 16'hcfe1;
        src106 <= 16'hf68c;
        src107 <= 16'hfe84;
        src108 <= 16'h6089;
        src109 <= 16'h70b0;
        src110 <= 16'h28ee;
        src111 <= 16'hdc25;
        src112 <= 16'h2f92;
        src113 <= 16'h89ac;
        src114 <= 16'h664b;
        src115 <= 16'h5e76;
        src116 <= 16'h6e4;
        src117 <= 16'h19eb;
        src118 <= 16'ha1c7;
        src119 <= 16'hbc90;
        src120 <= 16'h66f7;
        src121 <= 16'hf347;
        src122 <= 16'h73ca;
        src123 <= 16'h3ac1;
        src124 <= 16'h60fa;
        src125 <= 16'h60d6;
        src126 <= 16'h79d0;
        src127 <= 16'h7df2;
        src128 <= 16'h1f0f;
        src129 <= 16'h927a;
        src130 <= 16'h367e;
        src131 <= 16'h3b1a;
        src132 <= 16'h53ec;
        src133 <= 16'hfc1f;
        src134 <= 16'ha4c8;
        src135 <= 16'h690f;
        src136 <= 16'h925c;
        src137 <= 16'h5eab;
        src138 <= 16'ha37f;
        src139 <= 16'h867b;
        src140 <= 16'hafea;
        src141 <= 16'hc3d2;
        src142 <= 16'h211f;
        src143 <= 16'h6ba5;
        src144 <= 16'hd935;
        src145 <= 16'h62da;
        src146 <= 16'h9b7a;
        src147 <= 16'he61b;
        src148 <= 16'ha68c;
        src149 <= 16'h9a42;
        src150 <= 16'hba13;
        src151 <= 16'h686a;
        src152 <= 16'ha275;
        src153 <= 16'h3a04;
        src154 <= 16'hfc36;
        src155 <= 16'hf30f;
        src156 <= 16'h27f8;
        src157 <= 16'h43af;
        src158 <= 16'h39e6;
        src159 <= 16'hd383;
        src160 <= 16'hfef8;
        src161 <= 16'hc5e2;
        src162 <= 16'h6b43;
        src163 <= 16'hdf1a;
        src164 <= 16'h4038;
        src165 <= 16'h798b;
        src166 <= 16'h7ac1;
        src167 <= 16'hcaee;
        src168 <= 16'h550f;
        src169 <= 16'h43ab;
        src170 <= 16'hdcda;
        src171 <= 16'h2f5b;
        src172 <= 16'h7003;
        src173 <= 16'hdabb;
        src174 <= 16'h1410;
        src175 <= 16'h3969;
        src176 <= 16'ha46a;
        src177 <= 16'h85c9;
        src178 <= 16'h184b;
        src179 <= 16'ha772;
        src180 <= 16'h8a75;
        src181 <= 16'h94bc;
        src182 <= 16'ha5b;
        src183 <= 16'hcdb6;
        src184 <= 16'ha564;
        exp <= 24'h5c7308;
        #1
        src0 <= 16'h551b;
        src1 <= 16'hc7fc;
        src2 <= 16'h446;
        src3 <= 16'h99c4;
        src4 <= 16'h8675;
        src5 <= 16'hdefc;
        src6 <= 16'h987d;
        src7 <= 16'h81ea;
        src8 <= 16'ha7ac;
        src9 <= 16'hdbc3;
        src10 <= 16'h14bc;
        src11 <= 16'ha88b;
        src12 <= 16'h8dd0;
        src13 <= 16'h4a3b;
        src14 <= 16'hf323;
        src15 <= 16'hb93a;
        src16 <= 16'hc36b;
        src17 <= 16'h82ee;
        src18 <= 16'hc9df;
        src19 <= 16'h3bf9;
        src20 <= 16'h326b;
        src21 <= 16'hcb1a;
        src22 <= 16'h98b7;
        src23 <= 16'h1fbe;
        src24 <= 16'ha733;
        src25 <= 16'h7517;
        src26 <= 16'hfb79;
        src27 <= 16'hc214;
        src28 <= 16'h8a80;
        src29 <= 16'h4fee;
        src30 <= 16'hdb8c;
        src31 <= 16'h3efc;
        src32 <= 16'h66fd;
        src33 <= 16'h8503;
        src34 <= 16'hcbe;
        src35 <= 16'h1a19;
        src36 <= 16'h71be;
        src37 <= 16'h8dd6;
        src38 <= 16'h6175;
        src39 <= 16'h5822;
        src40 <= 16'h979;
        src41 <= 16'hdc91;
        src42 <= 16'h4d11;
        src43 <= 16'h26e8;
        src44 <= 16'h3727;
        src45 <= 16'hb2d6;
        src46 <= 16'h6584;
        src47 <= 16'hc1a4;
        src48 <= 16'ha704;
        src49 <= 16'ha382;
        src50 <= 16'hb36e;
        src51 <= 16'hf378;
        src52 <= 16'h867e;
        src53 <= 16'hdb5a;
        src54 <= 16'hef1;
        src55 <= 16'h4938;
        src56 <= 16'hbb9c;
        src57 <= 16'h9553;
        src58 <= 16'h21da;
        src59 <= 16'h79df;
        src60 <= 16'hb84;
        src61 <= 16'h7b80;
        src62 <= 16'he3a1;
        src63 <= 16'hccd8;
        src64 <= 16'hebd6;
        src65 <= 16'h6392;
        src66 <= 16'h2ca;
        src67 <= 16'h35ca;
        src68 <= 16'hc75e;
        src69 <= 16'h43c9;
        src70 <= 16'hcf9a;
        src71 <= 16'h9c86;
        src72 <= 16'h2c11;
        src73 <= 16'habc6;
        src74 <= 16'h5531;
        src75 <= 16'h7d52;
        src76 <= 16'hc0be;
        src77 <= 16'h3305;
        src78 <= 16'ha211;
        src79 <= 16'hf81c;
        src80 <= 16'h43a1;
        src81 <= 16'h2a80;
        src82 <= 16'h4fee;
        src83 <= 16'h7d9a;
        src84 <= 16'h126f;
        src85 <= 16'h4dd7;
        src86 <= 16'h16cd;
        src87 <= 16'h3a5;
        src88 <= 16'ha76d;
        src89 <= 16'h26cd;
        src90 <= 16'hb3e;
        src91 <= 16'h48b8;
        src92 <= 16'h1222;
        src93 <= 16'h46d2;
        src94 <= 16'hdad8;
        src95 <= 16'h80f5;
        src96 <= 16'h5bb9;
        src97 <= 16'h5d80;
        src98 <= 16'hee04;
        src99 <= 16'hab05;
        src100 <= 16'h55d8;
        src101 <= 16'h6e43;
        src102 <= 16'he1f1;
        src103 <= 16'h3657;
        src104 <= 16'hb7c2;
        src105 <= 16'haf5d;
        src106 <= 16'h858f;
        src107 <= 16'hac2a;
        src108 <= 16'h19c0;
        src109 <= 16'h9b;
        src110 <= 16'hfb90;
        src111 <= 16'h1b3f;
        src112 <= 16'h9d2e;
        src113 <= 16'haeb;
        src114 <= 16'hd9db;
        src115 <= 16'h4242;
        src116 <= 16'h19ea;
        src117 <= 16'h4b24;
        src118 <= 16'h75b2;
        src119 <= 16'h1918;
        src120 <= 16'hb93f;
        src121 <= 16'h4923;
        src122 <= 16'h55bf;
        src123 <= 16'hc1aa;
        src124 <= 16'h7cd2;
        src125 <= 16'hb0f5;
        src126 <= 16'h42a8;
        src127 <= 16'h207e;
        src128 <= 16'h29dd;
        src129 <= 16'hd40b;
        src130 <= 16'h6733;
        src131 <= 16'h97c6;
        src132 <= 16'h8304;
        src133 <= 16'he7b7;
        src134 <= 16'h73cb;
        src135 <= 16'h694;
        src136 <= 16'hb83d;
        src137 <= 16'hf3ad;
        src138 <= 16'h33b6;
        src139 <= 16'hf025;
        src140 <= 16'hd046;
        src141 <= 16'ha608;
        src142 <= 16'h363;
        src143 <= 16'h5745;
        src144 <= 16'h5505;
        src145 <= 16'hf004;
        src146 <= 16'h4a1c;
        src147 <= 16'he7ca;
        src148 <= 16'h2d18;
        src149 <= 16'h7552;
        src150 <= 16'h3c5c;
        src151 <= 16'h500b;
        src152 <= 16'h423e;
        src153 <= 16'haa28;
        src154 <= 16'h2f50;
        src155 <= 16'he448;
        src156 <= 16'hbfe3;
        src157 <= 16'h1b03;
        src158 <= 16'hcff3;
        src159 <= 16'hc39b;
        src160 <= 16'h9e;
        src161 <= 16'hdc0;
        src162 <= 16'hadad;
        src163 <= 16'hab1a;
        src164 <= 16'hb365;
        src165 <= 16'h2a47;
        src166 <= 16'hbb43;
        src167 <= 16'hbda5;
        src168 <= 16'h2cdc;
        src169 <= 16'h3efd;
        src170 <= 16'hc9c3;
        src171 <= 16'hc84f;
        src172 <= 16'h465b;
        src173 <= 16'h14be;
        src174 <= 16'hdb79;
        src175 <= 16'hacd7;
        src176 <= 16'ha8ae;
        src177 <= 16'hf6bc;
        src178 <= 16'h2ead;
        src179 <= 16'ha3e7;
        src180 <= 16'h89bd;
        src181 <= 16'h9f7a;
        src182 <= 16'h906e;
        src183 <= 16'h9f3e;
        src184 <= 16'h761d;
        exp <= 24'h596f0a;
        #1
        $finish;
    end
endmodule

