module testbench();
    reg [27:0] src0;
    reg [27:0] src1;
    reg [27:0] src2;
    reg [27:0] src3;
    reg [27:0] src4;
    reg [27:0] src5;
    reg [27:0] src6;
    reg [27:0] src7;
    reg [27:0] src8;
    reg [27:0] src9;
    reg [27:0] src10;
    reg [27:0] src11;
    reg [27:0] src12;
    reg [27:0] src13;
    reg [27:0] src14;
    reg [27:0] src15;
    reg [27:0] src16;
    reg [27:0] src17;
    reg [27:0] src18;
    reg [27:0] src19;
    reg [27:0] src20;
    reg [27:0] src21;
    reg [27:0] src22;
    reg [27:0] src23;
    reg [27:0] src24;
    reg [27:0] src25;
    reg [27:0] src26;
    reg [27:0] src27;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [32:0] srcsum;
    wire [32:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76d29cbd10031bcc9abe4be96784e9bda6360ded141f05b799d61b5dd029aff8bcdc7e76cf9102b57b84350a253b41d34b0a3addd7ed43d424315851311172282ee8a9616d0d0de0992018ee49cfef0cdd0fd487a0705f92e22fb6ae7dc29f947463;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40f48b407246e2f3993e488afa19887f8266067a6af6e8b564dca9f2d28104b91a3f6db48754c9526b2f7afe9d39221f6c330a4d3ba3e7352189fe4a40c55ea0ae7d8f698fbffd1779e1003f677e117ff52ca6fbe5cb8cbc9579d844ad0c7853f111;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81808dd542f3b15f44c92270e2aa78a250fd87d5794a2fdf2bb031876dfecfc6c8c89648fc88e7dfd4af9cc9af7cf8c18dd704268489b6fd70391b7d9c486aeb9bc72e11031023f8bdab13ca9448abdd26d2aaa76472d9a0ef9952966faece7e3d5f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d1e8dcf03db0b7866574cddb8cfffc7f8a08f5cf04604deb6b1ffba66cf1a7ac858a1a8fb20c9c98bca1b76d2458dd509b3fb12a2938dfc943a3dd40955b0021dbdb8e1a43d69f7bf8d58a8664a7d476d6dc487df0c4e6e3a77730d842f9a152514;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7601efe20de3960c49397ec81a7787fd5d1d3c82d67862d950970b5fd093537f0c15fd309ca84004f2cd43e98a1613a6cef54dfb742d70d8f7073f1658b54d3bfdcccc96b88ac56626260954d4412dea1ec17c068b2fbd472510e73734205d5582f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5654b2ce253d6cea74ccb604196e202b6d678cb04472af3525c2ff08d5f71a32e18675c20389509d1bc7912d9956ba3da2732c42d0fa84834278a7d931c2aa02289d528bbdad338cec55ba9bc34281b968ddd7896ca5385a89afab6d8e6b86f7032;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h213ee4908a6af38f405cde705155899d6bb02f8a031f8c4d6ea6141b21c2e6b82f7b593bc4ed76625fb8784fad436ac91922cc97fcdf0ab2f2f5f14cefe44fd374e83317090e44b48692664587d6615abc9321c7b90880ef67180f06e1ee45e59d5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef41493b83c79800889a4164701efec8bfed3b49927b9980d0d0ca3c9eee4233b7fc9af754764310f521c6a2a48e36a90ac148ea581338c1262a56bf1e91e32fee9e66f093650fac4ce2a9304c62ec29c23c746ae0c06f4cdf98fe7735bb1bba6853;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfee6ca99bab35053219e59f4a6ac189cd9d97271d091a6b108778a4e6542d7ee11e8a6dc81c130422004e305fbfc3701293e72fbacae5e9a2c2a75588739cffa15fa1aa86d3f11eadac21b0032caea984ace8e009474b8f0130542b7a5b1b5e9fed4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb731bcec5b02c1394ddbd314a4a8c36244d7a17a7668db8d46200d02e469bead5b8911db3e273c8ccab91a4f69b25e0f3f5cde4db9c53031d061a95ff8840328005032d5f5188cdd6c2903594013b5cc3e7d5d72666619c8661f87c269850af2916d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77b32d75044bda23936d77803738de127f6fff787e7b36176537952c71d17a3a3ac24cb7917949f05361e0c09beca14caf07e3aa192223aa8a4b36c14ad0c6a5e5bca4e11db2adce409e8f6f66cb44b6565927403916cd514a8f1b4193a05400d192;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c91dc52719b77febf0a81c6240b49e558adbf890dc1913ef1e18e6be5889552bbf3996bf8dfd91b3de16a1e31c0deb11ed608e9a5d5639d42035900a78a8b9d3933c3a7f9d34fe83c12d19cd305027b6a00390235f46873b1f86abcdcccd6be1b71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fc15b55da1ea10a9ab17bf9034a2bef3377a2757dcbe1be903e1dfcca301eb42b369b3ce49d874941cdd8dec64cb79a75aaeed6cf5800e9b84060674e21ffccb294ad0f208fba60c82db2a4608305a85dfe2b3cd886f5ee2dceab9ed3d224d72697;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6edc0748496795ea8ff1404d5a0ab025868258c3d2954d8ff0623f645b65434ba72a1955d85d1199d6a26ddf997738472cd75b0e7883f63dec356c577232146ca21b65f9b3e7c2f115e6a68525597b8b35c48cd04bf7c98990bf96a1a506ec6d45b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13208050429befcda521acbc81e8940e8158c5aa7aaa4ba8225e7bfb79a9978a40a9cee2882812ce1e6303533b6374969a9a5e66f339261968f46e9790249b777e70bbb56ed4d61d8c196c1d59b682d6503997988b041b1eef8aeb9a6eaa305ea3ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7f7b37672d2a79a43d873171035fcef29e24b9ebb3b74a86f7860356fa191a486e06b2f9a680b285fbb0ea779d6399f861354fcd6af9de460f2b9ba90472bddf829a1ebcead0ac76ca084d55a1251959164b2cbbeb95431ad2ef9a59a7a1e6685f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7f453137e0a71a7349f9d9e0347c42ed54b6bece83dee2470d45c51aad58f1f1278efc01eb80139acdb5366770ccef0f7d04bead75cbc22b7ef35b8114117b070a91a8b0ba6c8997eda36d806c639e41880478d4454a264621f8f9c0f74826bddd6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b1c9d6682c162aefed0abdba6e8b0c3214dd81907f8c073088babb8a7cf3aaf9dc46e82af50dbeddb7d1c14c4c48d0697cf8ff20f221d48b4888221edca4be8364d591d80d1b41cee2b3f11284329f722a8872e25f1a06f86a60120e07698b24af9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2668012b6695a3d47a938fec5333c470f30038a1beb3c5bfbfff361605a44b319c7c3d798a5835012c0e5410ddefefc5e2414a84cd0ec13afc9d1e94f2d4f97803a89b802c66479eb7b57c8e2caf9570e2611b286530f14574f1b739887a6be2a67d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cedd7d9685c43f8abe9b733a00dc44d3c77022a1c19845f0e7d4523475760c489a1c30c337573e982e431928b6f46f58f862138f91c7698e748c0f9e2878c2bb3e3583d9f89e59d3960115abb15c64424d69f6d85b6747b8a15fab7521f2615a362;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4e9a30aba72b55b48319ccace524e406d8fa73ebe4b80bec4d240e5b225c53972759cdafc5de8df7ffcafbb2f8d144b38a075d646a8dc6db174d15ac31d984e164e9b4d6e8e09397d27683f6a6f8ea6af0dd0cc07a21bea8d55e2a3d13256a075a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0a3302ba87dc1ff691ab457a12966b6f5d58659d6309ae467acb15c339869ba13309e7d78e7de9b0ac7cacfbbf62d615d0d13b9de62e5afabc21e559045a47be51476f386a117ea9e274366e3339c8e24dff58791cfb0d1dfbbac2f1e172b44035b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24be3cb94bd14d7e3d9db86afeaec7aaf3387cd10b741ba687f9690ebcbc7fd1365f1e1066a43b258c8e8af347d9daee966b79118a917f8a41e38053bfc363eaa71025598f6fee1cd41919daa78f028b380a47e8eb417ae652587c70c00d4fe2dea3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d8e9d37c405abac8af7aed38d733483ad73e932965225419c27e8139d9999bfaf8097a6239fafcb40d36f60b856c5a72ebe41aeef83fd0f56536cc1c31d47ad60cf0d621834ff0f097a7f59c9bad2749e32163bc4513fd22e3f527cc947148ba9cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa2354ecc38818d8a8bcdd1a9980a68f4a252724b3b84c5b9ac454dfe795bc3c0f35f772e1d81d1a020930824f2dc402c299311ff86895842e51c335ad461689ba2e75730c3c9c14974e8eafb9fcece63aaac87845620dd5e95767f8deb81bd234c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe4bba5d76d1c44989aa0e59714e9ad7c1583ac5e2876a0f5e7ac6ade3ece431f5180381110aac7880d90089b8bc18f307227b5bdef19ff7c7673f4f8e41cac7928e008d072fa2ef065bfb2be3f344aa09ce61b7c5c101236dcf8a8370c1e941ee69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8fd719cc343d4e42bf58f13b1793c8f59ef4c943da2d060817bce803acffb1743cb51f6f76eb3f704f1a3fc3229a67996b54a81fe902a4e4d9b2e0ec0696bfcf982fb3376adcb276c62d1423236e98a577073d7c3028837b5b970516272271bef68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haad6422ac1245c3c727b670e9c6fa08271708677d503948b66bd792a26811798094cd55ec5e51815f652f67c4ce528e76f7f1b150a4fa6a67e09fd5d774237652f2e319ec0da51226c3e8b80ecfc58c6ee076c1a9aaeb70125627e04fee366773db2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f8da360d91c79e362b807038d7d517f073915dd345ae2553618d49cd91574cc81f7006c6dc68d3bb5e96a5d5d89f8a67713e027942274440c138ee2c47eb1ecb15d085afb29b9e8e53b0d3c4fb1a7e2eb4c80193543098eb17d33e47bfeb44a97a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebf8f58f56411ec95990ffa575708823830b157bdf7dfbab43b9069dccc09e316f035d10838a287de059a911bc29603639b0a18a000cf1bcc9c13a03fad2713b954e79d210fca7f6872b390cf72ce30012ee76e2e256c6dceb504576240ac0f3bf96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe38fe9c16194eca927dad8894a2a7e0f6a14ef3a02f388a3458d9887b01514a2c73aba3a10f67595c0f96acfde543e1f0b9359366799a2ecbf42b911d9ad40c925ca041fe1c454019d613154f531de33603e749cc2f99dafade000228a6d7e1cddc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h737b148e47abd1193fe3e608f7ae20684b3ef2aecf7e4be2a127283b68ef3662b80583b90fb38a6ac3ba393df1796a79abcedc1e1fb969d0a6e93c490fe9b17d953da9b65b990c011db35943ea7f527b04926f77fbcaec1ab69e4b31125e8ec09902;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf91bb7be1b529b8bf026a3e1a8e393dfc7e22a26d66a3a98aa186aea7ba354e0b64c0e81689c2a8b17f3aa2df69a3b4e96bbad49bf4ca552bbe16b15ab95da57754da826557a55debe1495fc64f9e76a5bda5791cf74704772101480d6e6c0fbde6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb3e55dc325e6b83d8db072d9fe59892eba86e75c88a6daebaef85294ebe566a26a5f75d2ce751bd6ecda359204b421add060652ca58b84569c91a794dde544e50c535907c7a47a1db783519288bd65e71192b489dee8fc7d8738faba6de71dad46c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67802f640e732ba9edada3db6680db4fa019b833c181b70fe7a152a4c06f71d9436af995ccf9f1c9bb619a312b0ed8af8e95a25ad1a2345ea43350faac191d3ecd31233850a8efedd628093820dfc740c6718202a2ceb326a3094da82b9de7e6fbce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb65e1faba1b11c838f7a403e96b19fa9506ac8b982ecfd4682e82ffe192ff13f5a01285edd90f262bc27a2c3742ff69274bec14e99e0feac4288b0060e76f1c1bdb2b238b503eb3b8e6d34ff537d770ac300a9269f3ee9f6cdfdc7fb24aec454f9b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcc67a57366fee5c975bcf38cb860bb89323f527bbf7c26ef3478aa93541d112851f50100442c4628a2077938d83b0798b28dad5d0b3bd6b5eca9de3b23dc1cc3bf09cf1e6a601e9e1813a2aa057d1f1d074d7c00b12d14f275fd069adfd69870ddb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6082ef5b97715ecb434eb57a7e1afe04552c28567eb72d05894a7baa862daa57b6dd78d971031ed72d35d8283991dab164fa684996de0a17e26798cd7cdb3bc58476a2a0025a1b03aac82a0056f2c3956779eea032abab144fed3611c40b1e0e53eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb27cb803f41d70ee465dd226f7bec2f3463d2f1c7b0db0807886ce1e227328e1eb123f613352c37e47d8c24fe730d6bbef8a50ac0971dfa59ab7de76ec3d4e9221987e9e04e0a1abbfb7bed5ab244d7676675689adf6d10442b4febcfc666890c2d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8e7be49c87b0a1939284b1e6f9ff39523d14dfa5b467af23ffca5dd0933fd2428e21149ab46d5bd3262d1c5cdda21b6501f3dca3ef118893828da9a3f203e52b3480cdec0ba2e88ed200ce7070589d2e45e645041162b213456f7e2ef3fd37019c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85cbebd0545d430fd05aa3c5bce711bd3d2fda9ef3881dc77116574db8dcf36c8b2a9bb9c0739c4181cda34e17cce4310e20ac86e5fde1db39307eeb9fa516accff997eb60155ccfa6685ca3be955a101c0021eb11ee84f1ac387acf6002d168ea4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91e8a8f8c448b06aa971286707e41b3e40aa9c74903a2f165928cdf3140978cbe04649ae4381931997897cccda85be18ec81747fef199e156d6282e6da8525f3ae0b9485af6c3371a86643262685f650a83619f40fb9e32b88df22455e089aa79d4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19fd4493512b22eb93774ad857d062129f81b50b58e274b73e5b2f73f607230732f261942e40579e805ade472f4b8c61bd7df71e8d4e724a197a00df48264af154cee55059cb20ca83732b2aa80a38bfe17e081714c171a2239d199c4ef1054f9849;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf3686a8d1b53d5d2b887deed4ad8c49399d7c2c71150bf2d5ac7f69669da0740e4cfe450fff5670585c4b2e8e9ce05e69b0be8583de79b668fabc8640a6ccb3f7138669e3f2663be9359528283b1ecae583a15d2caa7d2e022d0fadbfedb659f84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2b1e84f43d92ca47d0b07f9b9ad7174310c130f7622c80e2ca50fea8dc7688aa45b5d6a47b41f59a6505f6a1b2b9a3d6b603a5846ce26f37624ce448331ea487b6735cc8913c089eba84142b8345b1ed51b247c70db111646576a8b35bd8a688e6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8062c5382d831d791d2194f0484a40f3df48f4406abb33ec397a768212edf110235dbf36c76a5302f71ffdee212b4fc01ad5acb662dad3ee553a86fb3873e22e1c6e244b205be3ea3f7444ace36d36fe302e1863d1267368567356e2e07a6b46bcaf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha01e11a1826d2bffc211f87484083b8799aa57932faf9749667f3f62a0514637c81c1a3e5c37470b76a81251ae15075b541398080353116e1d0b05ce4c78b885033d634cc1823b3e313c06b9b76f141596c22f60c885c5765e634f1f739d22864832;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h821b842ffdf5e1442bbf80c13fc56d9d6f3b35414a308670e04a2b815f0aae7c96da86cbb7c29292504ff94687dfbada8c177cb5b17d7f71a8715dca4677064e9740e23b3ad4d7407777bc47d92f3202915c41244dd7e06847d91a955b51c634d1cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had5c89685937e90e7833a5efd46e199c8833b5aaac56c9c07f8b0f0c835a12766145d172e110caaad10ed5079b2253958f598606b20a753a83b63eae491b09e862db897c65c868acc9f36e7346c8eafc77e0694a567233a7d745410752714be04937;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fcd81d45321600681f12969a728faceb76b83510302e6246eaf14a94715f73ca8c545eb956114b496e6d7ac72209bbd397eaca10dcc9f45da8fb56c8b1438d5c807e899d27f06bf06f0e45a692b2ea24af7da42fe7ff5108a339473f78543f8fd6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab77b987db6e6a26a575dac919ecb6002c05f65b8fcaa0e28dd1b6e82b39ec4899179cd5d53efcafa85b8c192d660ccf3ed6eb9b1bfa5685bd84eb910929964645f414c48ed33b5acdbd1c534d048120ad31abb6918429b484e30c05cf4e95bdb843;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h342e35c43414dad27cb5c9531521335478244792a82446ae3164508119bb8d48ba62bbff1f593b5614af74d91570d0868443fb588dd10a39001f9b25aad337f2deac15df1d558c8d45bf9e8eecb3b977e203347b14a91c5c2f98b2ab83a2f7594c26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92bef4a4e2d2106633faa41e40664766b9607c4e2b10c018135fdf3acc491551dfd69c686b409e5dae53733f6a482626f0d17b7ceecce2f9712ecfb32e8db0b92dc1118c37d52db4dcc8674961f5eabf614db3a63db56afa413f7806e97a4c527c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe3b1846472230e85846de7889b6acdb82c1311c961cc03d4c3e764b16c041807137bb4de2bef1b8752346cf74368288ad3dee49d22456f9a78950b001d59c17f0b7c0f388a7c74bd86de5d15b2aab345d0ce94634b677db627b88d08e9bb77476a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0a36d7e1e5381a19ffa945a6c7b87e94ca9e935a3cc5dbd4d5e72a0aae08f8e801e05c8a8436267e5329c0984da49279239fc4f9607ef2728f165c8dce1b95140f12e9e2b84ccaedc0f19333ac5a1f461d7f361e4675888d9e68c4735b957fec375;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a306112a6c6792e262031093c9ced44bf09e72c11bb02869abe946b769e1cf615bae484611070501cc3a8bbac519b2cdc06c7c679b556a7e045580313b87f5d01d986ffa345550097299f63674f49d46c7cf52f1c554a10ba772443e497241d0a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c4c909670361254fdacce85deeffb5082bd672bba2b666f772031453a6e20c8de7397b68786cbd3334f781c4a1b55731053076fe065d66ec5f076d85d901c101b6ca0f0b62d6ac4bc1f6731e0bd0d14cb630b3119ed9fa0d5f07496daacc86e50e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52f526cd08aaecfb7da53599bcfd21f6a62a263b69c2c7f26a7f3eab77befd7897e90ea950e5009dda835a7d5a639362eac8a3e5d5eb8f695a659c74a3254a042cca148ca948cf89e6c25a0b8cbfdf12f30c922b02c7befa1d13c2fc4faefdfb8ea3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h407af2f7e1181f6ca857629ffce70e8e02b59c743c8f88ae3332958ccc5eab41e1c4e42f435b4fd3749e16c10459acca44f7e961ed2d9a1bb7fd191e75ba2586dd5b354cc2b6a62d238a36afcb974cfbc48d48529f9c00bae20eaff572c8d8d0a7e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38214b83c07b8a5983b4431de3fe0220ba9a4014bc000c377c9dd41fbd41f9a850fa8d57c726c872a95d9462fa17788adbbd0c503a25cf63d6d2a81f1b233ddc24ad704a2cc4c2718f2c6801c8353e0036975314615248621e3c96feb20b09b0f755;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha18215afb2efc192b9485e523b7c9c540702c661d79b2c01e8929b87fd3e894cad976959d8d78524812903abd4b4df3678bc71f1230f2d99421d1c547748b58084af3620c027d42b45d89572d6e042ad6c6385636b23c798a75f6d02dfaa84f00924;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98b66c38d287c46989555c6f1087644d3c3568c6d03af9b206aa08a34e1038ad2a5f55ae196c4d9708770df9b9257da146c69bed5c8c6ca56bb7c70928733457b4e0c3fb1459b0b1ea22fa35fea4fe2fb388c31fecb40fe902de53191c1e68cecaf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h801af1f58ae2d88e8438777e412432160b28705befa3dd6fa03045f28db66c69feb75eb57ee6a3de575be55ebbf2047d9441f325f0ec1031e72573f79f87b6a45837d08269442d028c75da70cb705130dc0cceac93fa65f84391cc5b53d7f290df3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f19117e78aaddeaa863d2076239fa750d060fbb36cb7d4563e4790af0237092bde32312cbdea8bc65c6c3f7fedd2bfc5239fd7bdaa0182bef7433f5f911451be49c6511fd3ccf77a7f45d46d9bb336cd965ec640b3213bcdf5823ca7c1acacef5af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd63fd4db001736341acc8ade766a9dd93356d26bfafc24b2f960e5d7777593edbec91b00601cc94b5865fcd7764d92aef02f1226c0d5904b2de44747a7773867cc8b5f1efeed2c01d14389fb49b907368f6fa470ed9597b2b42789bd0155b2c8e98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27b89c5627b5d33c12b1e6c56f42dfd0f3eda169b34aa4fad122e66e9e527043daa7bf5469c681d8d335255ffe5dd800ba3633a7f464306c8fe0522c21f880f3b4f696fd8f11788ec66e1fa839a1ac43823fcf18fdff94c9a5563919619a0120e538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15f0618278b0ed93be678121a61a164cdf2239b51541490fbf0c4656647ff58fb4294b1279b611bbcde2f1f74c35ae7a0ee6654826283fcb6041350765f4c3b8023b6d498dc72d7fd54c6ba81e1492939c9f1c3b7e301e6cbcfe590b5cd0d6585a79;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53461255ca5ef79205ae019f3d4c10609dc0037903c70c9d9b60d81b8099a045996f4a52cb4f9880a6c955629802c70fe96582f782b35c18c5f97bffac66b896e39214b99d8850b6419357672d34219b9476ad9bdc9c18df2b029455201fc389d1ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a92fc792a0a477d44c6b0a18eda367db131b84de3eb7538c010ae4404577ccb265d468631123eb81f2d4a613cf5289b60938120f0c9737736537fd585b3661a1b44ddd7667991e1fe739037b5abb169231d322c9c421da06c5fa626b6c8ee35af7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40346bd31a048749e464e8a3d48d61dea15755ac8964a7973b1f200742ab407de46bc10048bfb7b02e4a0ecf5af1e2b9c88419e6dc9b9e733101986b5f3da6a0fd7498e414094ff1053f93bdaac5a8878b41e77ccdcfe0a847ec63b31ed35e795d53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5a705220f5c9d28ea782361b7d91f6111c5bc0953a8ec694a4f89114c25b5fa37b0d8056cc182ac9240cb853cd30cddb06601dff0119c886affab09fe60f45c0093ffac75b5e1eec3da651256043368f8fef3d781cef9de1c830d8ee3746365f868;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a37152d1925c0db26bdecfc853d011eb8f27d6e012cd140dad8f9ee9b345b8b5e38baa3ee15f896b01a5ca1b26fd8e9482398928e00db752b010cd28af12bc2ba34f218c63b0c3bbeed70f22084b900b11f4b197e0cec6db73a3cf7d34f215f97a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1f03f6dfa133aae38349f29a7403b5687857e9ca5ba745dd6b216542974d18f30d59e2cf4d3c4bd0828ac0e109b429f7a67e8335b19559fd800eea8312180d1e64f84a655e894aeb502c84b9aee3b3c1c3f565a4cc9c488cf49d2a133b764f4b7b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b3adb8ef6137b77a4b2b8c1eb3422368447d60a47003931124e88edf48e39ce979e841f00a1f7614fd679b5c4be26a8f0a183b9efd3493c6fb99f1a90e9f09373890d8aa44e3c244498b8285e8ce3ed44738a832112bf391b207712824f46be7ccc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hede63bc24c3ef2f307cc0b007b72b03028c0c5381322e018f21482942b588376e60cd75d8e5cbecd34b8146b3e685b9f43e1ec26e209510a1c71424e2bfe20f07aa771859f3a8b568f4d2601fc4085794e7b22cbbd82c263d87dc67293343d99891a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a21285e3f2e9afbac6c494053edcb569dff2e184ebedce49d0212015c2ed5b09fe17c999e81042bb82aab4730fb080d2d88180046b3dd3c08d83e41922e8b3820151763911c63d3a88b938310a8cd83e297d7b7cf154dcef0e93f457c5bba6c9de6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he88d98efdd475e0197adc5d3bddb585dfd50f0a9bc93ad66d1adf0f8ed83140b4e01699c74ca9e9f468d576cfc03a839849eabbd7cc670311f590b1903a805e2b23a0654377248ff65f7e5025f2901b1b5537bb135e93c47e49d7da520ba58482cc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69484975a75b5b4fc3bda9a38edc716384c4e4a4e4c3b765dc05c8a60366173e33b2d5755da671fd5b49ced7c867f96902e6cc2049884f2823a6d0a6895f298e0953e5b54883ac5d6f3c7f546725077b499a8de7b109a24990511b0ed4ef4acd5d72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h679a713df8bcb4f4a5bf9e91337fe6cb4d2cc1232aa07c2a8d959fd96774d04da94328aff33b5618b669232632e56c0b41cdd0b362ed03c120de613a1122e2c58d1194c4f6fed450a84f0852e38c9a55a728f42b4638018d16d1600585f9d3e2f587;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10e96315cb77322634b85a17b2761d49015cc31463b8d710dcf1cf82001347f06e4126fc2c4daa5732a55d0f8328014caa302ad6b3523b807337f0f534e7164b058c2f49905cec66fa070c8284fbdd392ecd34f003e2949cd519274e4eb60010ac53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8e637ed7bdca52f36a338ce18b56c51c566da3b3f633a12370a5623e4515982d1f763d0d60d91c4142a785d53dab7863bfe1b03d1a8384a5675bcb81ff0ce7ac2fabc171e28474c353e0dbd3e3846da5188b657b29027425c87aec9c1c27bc9595e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87b80865e9a58c81d1d610cae5992b1fe57f6a0d82991d4a129e9bc2b9ece7c7857d2dbb53cdd072364ff2ef0eb9bc3e19685716c2289e2b81cad10d5f444ee30fa6b94033e33a31bf19c23ff6f447f58d8872ca7367aef20d633b8e329d320be93f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb731905f33923de622c14ca319140bc3c65d141d6c0aafbaab73f0c70e32e60f5b867f4bf24d0df46da9b0c8f2fb75861c33c68e6482f700d1891952ad4047bb740290d462c5cad8a7769a79ba30e7878c62c9fcbf32efdcd5956c370c11f754f15e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd399d5688fb9f2b90f344213e6d705a6f71760a40896c6d1b2953434fa91e9b029caedef3162f1cd52091aba43b257e11b97fd4d533a816212a8cb48712c1bf42446fdb7010c05cdc2afc7ef512079c99115894542abe50ed5b5feae6e27fc588c63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ba26217c0d16babb890040bcc66bd3d0fb6fee01513e7dd2933c74c8921312450e5cd596e7ac8e4fa21ceb3587855bea86df524e037f13e0bfc9abedf805bb1e713dbb0304a3a066d78c814de13fd51f4f727a489ff1eefe033c61082390c1b9d74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h156ff9fd8fa3c3741afca76e9c4e8bfb942b5776cf5fd7c7e6f60c7da221626c4874abb4eaf5681a3e6a47633246eb74dfa0d30df83c645618e492b19539f34f437990d419782218c29f1fb658b9b04537ae58eae6968c2aec168a693138322a915b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd26846fbd944821398659881248aac56db0efe319ac1bf010fff0aaada1c87daff78a55f968b846519e8335d9477a517c92102e8b7ff3959063cc6b0874186998951378c597c9f1ca14deaff0ff8a0c7eba64c89e1551730487da482cdb96c7987c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8ee9796a6f02833abf525ae9019e9162b1b943d2b1ad1356e0d33872613dacb7311e79483cdfeab6acda5371a5b05088df723d2a416bf8c4fe9778e1f251af156fd26b3e586096b4596924ab314079db12f74313655ae7f0f0087371e05e1b6c2eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fb2b5820b342432aabcf63f0efe660c29f519eaf77fa2feca726ef8be127c843aeb1a936d4684cf1c0b9db5d3c9b5acba685826489bb16d56a72f067ae88ad6fce2722ae04f4dc1306cf2b8de78a292340d9b58e7d69d28a1eee8e2ce1e29b72a82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37c8440534342399e86f3a860b3a4fd34601acf5c38036a7158d54053962d09ffc7d4bb4a096ea84bee8b6dd5c7518b1047be5bbb422a2a9e590816070990d992e6d4ccdf8a21e3c897e151d581448ffee5d2e4d8b718853c62fbfa4d8f904cbf5be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h587dd6be0ccf051bd1d30b2e1d6650da26235e2d81735859f97e97ef4520e06ea8c4672117d911e4cd05a21b68fd065b7b64475e7179d7b0e32d382bdcad90768b5aa49523cb92ab7013fcd9c9dcee8608bd45aad5b0ed60736ce5e33995ed445724;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b9b5d38d4db5a59eba238f2b961fce0df9d81147b699ca7817a265934cbbfcc7dabfc8992ab0eea0fdccfaf6ebdd0f59cb5e34d445baed3ecb4b4d19fa586482e13fc4742aba8981423569091038d39fbf3ad5cc7c63f733b9ea7019a3c6759d6f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heac791f2e6464dc6b5078f80da634a314f83e584175d552e412d33408219ad1042624674b8c2c6bb43ce20471b4d21f2b42e8ce556c0585a671e0988a92bec4811089d97fd0baa2ecb47e8407e6a19782b2c797105e53379c1450a50eb5399d5e94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc01f5d6ff9c4d665a373b18ac2ce50080d579060b1615f18b9357094678a09940077f252d4af26e4754f6a30d92f411b53cc6a94a1055844a0f85dcd6e012c7cbe0083cda0f1246b3f3c94b0765fea7e9635da13046c51b973882405d79781db08fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb23dba5a37cb818487c7770b64879a0c2d22f7d983b0018b4b359fc325977afd103b8d2cf45e7c26301aeaf4c26f2bfd2fb62773997efbc441c96f2b97092f8305e1d63c3612836e485559b8345db77f8a9d5e3298b7b41b209455b36e2b94327bc5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a06568408d44f551f3f923753c2aa96414b67784e78f376e2b94d93a3787435a80996c0cd56cd449c8fe7faa2e0c9979569742f6f703ee2cb71033d9b03e9e35364a424b8f9c3b44d6fe862291306cc584d67e30cc62ea36999788198ac6341b274;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf06904ae94ee322c615a2916870e4898018b3c543240f158b7be3f97301d7bfe0810c373f115f6f06e51c2ae99bb3cf104e76fc77a8e8e3e0420f42141c08636882b1ffde761972cba8d342687ed0cf6525eced1169eb7c570386589abf0508aa8d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfba878f159554b069ead30f2a1e366aa47a90e107b90a4b61a6e2c5c0c25431e323a4ce08cb072eab4a3f375adb10ef4a34c5ecebc62718594e9f9ba7fb85d9edaa5c961a0148fbddb13665077987ab35db0b87fbcf8606fe9428c2c952eec77eb0c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fb09635713f932c1921f97c7d083f46cfee729b5cd6401e6e5800d9340c8021f7b8269e01493bae8aa0e76929224199374e85bba2c3fffe786c38947961be44713888d578440f0bb5e71a2c08bfb4761348500be5fde4bc189ec2125639830fb9fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28feae072f7b0a47eead05e6ae41566079627aa6fee8ac4cc7a7ee4e0a24245b23051463fed7690b109ef41e3772374c7244d73c18ddefe4a51876ec165b3a24ddad30dd338812aa0d1adcfad884cda64e42f402df03be419661bf02ab7b9c09c300;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11e96b1ec6d1f181e4a5bb437f23e3bba1d9628d2947a5fbde0332d08ba55ee8eb7a955b7f6e288bc980224b716cadd322f7d42c5c60ca2172b60a6481e88c13e3d27dfe0a4f384b4f96f92b816d6dd22134beaed31f758704fb267b19f5a89a1046;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h634a0d1b26c0cea09a8ef2ea49e3b89052960fa96244d26b5ecec0d66f3a862ee59cf4710beb498da8e978d45b4e41ff8cca6f6780523fb41342b4a45f5df33c7f7acd6be6d29b3f26a8b50cc94d9d9fb12a9664c7010b0b86a250100e8cc10a63f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98d0e5c474828a72f8e93599ab4312e356600d357621687bf235dcc97d9e415bd7e1eecf0954ae95b3f13050fe3281e1e28b786b59dd02f7f7f2cc801968462a5c8df2cbca13c5bcf0f110df3ad5d5bf85b85175b8924e008409011825a15f174c5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h430e5e876890e93e4ef787fbd377abef86146789a4c96839121244820b67e43523182b496a94a72d7694a731456e5ac3c0a5ceffcfba29d3544f309f3cc6f9dabd265e271c2fedf46acbf9f85bd5d5479e18a897504ceeed320e637d76676fc7bd23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h122236c829da1f6bd253e2b7cc50a330de9a71db927ff8e7185b55d3dec67e9bdcdf99898fd0f5927cc3983c62aa28e13177ac2ebea0e4c3354ca069ab006382f74103a02da6ce9ab1da587cbe040568f57e17d95b9700821574a59a462bd8c7f851;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6056864b41de10831dcdeedf7ded100c92cde4c53dbaf66aef9106ca109e02d731917904356f753c8d4baf18651a841fb408c1d84129ff7d9f7ee02869b2380ded11cfb0b845476da02c96126e1083ce0085019cf778f873747c2cdffcd3d8ebce48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9539e0a53fcd210d80e871e17fed636d9ff9d3d94539855b5fa36e152f943bb6ce736bfa441a31e6d642b2631d9b627a9f102b520e6a0c76abb6c1e1ab74b9dfb22110f24a79c6857dd753328185615abd2ec2bc873ee48248e34dfb3422c19fb8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab635927c7553ae478478a0a5f2fed9f9e01ae80695ca91a33904c85cef409f76660c25d453ea0d8eecf03a01ff2fa87aa25b3b847611cf70a0a149fc0c5b6fe165158db1dba5c1204c08b3204242646f257c62dc2c1b31c8be38e09f736a7c2f3d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5717adddd5143cda430b91cf846ee5e3230fba7b3a506810da8e18ce7e3ee09d5431c3df38ed29b68b08a0a2e20b2bec737bfa3af44b64478d7782b82c491d8b3dc6a3ef774f2b85c38b379f4da4f96681dfcb57e14b37546b3b18577a541be7a05c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45dc19be3a15871c520c9f712019746ae8cf018bae36b5e88e45c709220c41a56f4785b6bcd48965a50c4f2a849c79898cacf8b736cc0694ad27bbf17211345b8f41582922212cf2945621447d8d9dece0510c9387edb8852f0394db9cb3de457e4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee3e202b1a965763c80e888ca8707ee8b088475f2498424cecfe87486a24f33b7b17c7430f5df04762f2fb605a42182689999f44c6bfa4d78ec8be3e7b9edb4bf36f1b7972730d5fadbbad95f83adb107add457142d8aebd600d81a20abbf8d78e9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcddc3c02e818a04986772a137e0757c3cd778b960f2a802045c88abe1db9730b6764e99b3047a8ada400ed35273a2d609c259fca29442541dc3fdfda5f8f6ce2a53fde8e7bc93a945d72ff1584d8e194f7b3010aac6838414b8f4db5bd242c01807d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ed703e8bcf47756c956b0a63932b2a05d84d0379ea7791927bfab986ddef670a95e1000d46b3c944ad531fe1685cf5acb0e45bbb45346525a3d305d96f5d47beb033d346512039db33d4eb84790d6ad4149a4bfbf65d542cda8283574762c5f6e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h715c74eb4f7ff95c8d8346519bf3934df89868313b31afd941d25ba22c3469095dace6bccbc8e29f7aa3f71fc55350a0ca39e54cf8e17ffe4966dad4568062c41d5f1013306747a82ba591b1a2659cf018d05adf8d1dc6630d1d5208e6c5897a057;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61496ce6d0b424ed6787ba5d9b617257084bfa701b3796c01a081514265f67447639a75f5d7db40078301a016b8cfa4237ed4c9f8a0b4045436b8b07db951704c0bc9d76dce5602ce2725f2846cca1efe233d05bf1e171f605d7349a98e5f2e77c27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fbf2cbc20a2d21bb3e2d02fdab092f352ae3dfe47a615a44d7167c3cb3eff53dd1fa095d6efeb0cb96da5b1328f7f831d18053211a2a7aa752614907021648f538b473a42b39b157cbd407f4ef4ec6cb1c73a911271721348a48b8f04f48f2d935d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf33ba3d04bd90d129eded2b1f517d369bc5fcec34a782a4de437841e9fc6a1f73b41259ca04dc86ad98ff2e7b077f5130c3cf901b188dd63edfd86a7a34b4b36b350adc00666a195029a69f3ecd60f78c1622c1261a1975b1e87ac7c9b529514450;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39a530d8f2a607c443e989259b69c1964dcb302002be22b1864caa59082b25319c061c231f3eeb5b5be993acb234c25640c40f82337601d572b1930aabb4ca34595d7d3fc27afd85c43ca3c552ebcc180945e19e9fcbfce50c320bd8c132ac4c0868;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6c0371b6af87c7b7e6b567186918d646ef253740abba329f23751732ac61bf50e28c2610b27a981263411f1abd66b5393a3c08f4c6cdfe14dfe81d2206b0ad1fcfc431b962353cfdb87b0ee13c052cd90eedad32eaec962b405da345b4750f21ba3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf28eaa7336d0cb8df11764fea1aad468a875a2ea5b8deb0b92b9f3e84752a2e3737c97944d5a7ff4d2e8f5f61c96636b2e53216c3a19f8bce7d37716eb9b8b7028e0474ef678b1f6b51f1b48bf33b8630bcdec64a74c1c3060853614493790aca64e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habed57b491c0170b4bbad023a7ed158a39f7b7a9a5bf879a6231e1b046a2c29c9a0608298842dcef42961bd9c44347f1347924a8e8329d015eac7526d3e75b1bdcde5d23a4624d34d9b793753ac877f6818a9ea189c34a350ef7f6c0d261f91b73b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7358452d25bc0a45b5608174a2f6ef40c2cc9d036c256450c83b8e032a88869ffa67fa9b57c5de56dcad04d89f2b20dc189076bfa03a41f41a9c9521a7817e8103981c6fc7c491942fb58cfc9d0e06aefd42522c0d4618563b882e59c2c01eb82f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefea3dac01694b04dc08890db5e7111e3392100531f17eb693cd345dc1d07e20c2dec00177f381fd6a3272a0b41fbb921b3b59b7487a783b6d8867ed489331fbcd389fb8294188a8422f659d97dcdafb3ea040589385393f18828ed5b55c802ab42d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf547e4995b145acbb7d804275ea8646c33e9fcb64608f0ab6c6833dc91dc3d6e46a9bbb3c177a0e72ee2af621d15e68ef6a57856ce900411e6b24545eb025624a9b252bebd8c712674d58772e82b60ae1364924784aea90299ec268e8b8bd171e001;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4618f6c8a11af7206acd74e76088faa46999f0d8514f8c7be5bb68d75bc40177e8d156112557662c032d6e617e47c0ceef2cef8e05026d652d52168a25d145601a126ecb1f5004cdac2a4930bd8f1c2647ef96d5d0063e658f57c1673e53a080615c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba1593e41eec32468c243b24dc86d048d0a5cef443fb0b75e70054120183ae0c8353216ef5c740167fd87a651c391e02c545f16b23bf88bf6ca4a5ee9fdb98b7af1fa0d4cbe6fe36cefef6c94d9f148b7ea630fe3becc372fed070ca3678d6c732a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d2a3cf8c8333c861f35c74623b00cb8c5d93ebd4c8c0d15dfa5820dc4cfbc7f339ac7bdad34663d8c3cf68be9332ac23277cc9c3e1e7fdf041ac0beafc073db29e46d5e7fd9878275a292e896edfc94bf155779d89ce89abd7076e0540950dde5fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71e956c0ded7d01794bf383b40d97a9c3cb40c2f326ecae6d8a9dc3c86d4ca97b6b7ed897df58013dfbe249f9cc8e3f09ff13e44713c5dad11fb6ca18203d6b3f983ffec16809e39fd1d78680a2455e04c0ee835d5b1117c3b088345b28175ce422e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec5f1516f569fab22297ef36b79c8ff76031a75e841515efc5f9861bc67ac7781cac4ac6b51a7e60f1fde3d7e1ac1433a271a346afa77821603019129a62f88f733511679d5692be69d07c0dbc42635a83f4bab8fff209c57a2f841f50d9b3dbf060;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeca215cd3e497c3f324e732d57acddf6f60f18953473e458ddd955025abc17fdfbcc6418ca81028eff93886ff259225ef9c87a701e29d8a441d8b3cc2935bb3a493c7e610b1efcbf640f65a49925666f122feaa8615e53ed514405bc4ed0900c262;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h718f85f6973fe5613b0937506362b13d376ad8c3aa17d43c9a42c0cc4f00dec4cd8b9c3b9297094b15d268dcea27046d00fe9961611c0a6be7acd5de5bed9c17a6778ee7ada4ee0f4290309745481d161d71576322a8c8c8e379828150b66be8c581;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1ec0dd85318fd3fe9a14740dcf2367c213a102aa19f315f4785cada84b6287760de521d89419732872e3bdd571ca1b7eedf532dd58b17743ca708fd8e331049d8324e156ea07ba0df30d94978ca237f0767ae5cdbab3383d0cc1f113f395d14b9a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44e50e3f0bff152fa3fe1c314771105bdf5f139832cb6472352774120966fcf3ca03078e81941395387d1a1cf3df569496e1cf84229c5414978f885c93f4a4d8f48b262732ebd7055f19410ea1b826cbc1df6bffe8f4e820d7347b3af1b5c3fc819c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb59934390e376129116b5682b953ab1c90bf3f5001ed1e8661daf91880d3ce4239a6b83d04ca90822940b7321661b8d89a9f28061172552a1f06877cf810bb20102864aded6bd2a8c92c5f10bb82f2373094c1815ab19a227462cf8573064fbdff2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ac4be1680934cef624c5f5398aea56aad3fc8ac1342a1626209fb6289252f238059162c9e83a023075c8ee55d7973f43cb28dc78309e7fdf31bd48428d674920241c5386ba7d64c58a02b4c747a7ea87900e47fd44cee55c27ae2479f6df6b6b58b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd36f246c65cb13fa692dfc86fbe47e86e374e807b2f448a84b49aded79e4c5ced8afb9074dde7375b53ae025dfe7f83955149304b0a27cd3ae58fb40f8617bbb9016a77e77ff0fbb17c1c036865baa68b24dcc473254304308208f0c774249d964e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6de31b7d7f5c088a916bfb2ed84d8b2c06c5075bf81595b1d5a295a1a6843af01752199d94df437b7dccb2d8295d49ecf5b4eb3b18c575d7ca6c8dc8b0b917bcee2b08ce0461fdace6072edebdfde39535c420ecbaf2f7017210ad408e02ff7f2cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3eb90fdfd9ee75b4cca290e3efc2c3d117cb0a1edf0b14e5664b02bba2ac50c5831f363bc2a9df9d329f9b82c2e7123da7dfb70b43361c8b7f11f0fcaebbfb3828ba513aa9dc68aaf6e461d26320e0e38dc38f8e8d7acbcb0c2f2ae283cb6b89dc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h732d499b31eb88ad4f02a0b4b4dd437007f123548df1a5fc5e5e54fcdbe500a697dc5ae69b65693ab731805fe62b07f589fd3a03cc188bb1cec3501df2a5069e2786b31f4ece1ecc13c4a1daf974d961def9182198cfe93ac60fec7a357840c4419d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d83187047d19f62776e4e008d4c76dee584d401ee246d2f41372850ff33e8e28c5a7798754d3b5e00056b6243f79659a0a95bccc9c6adacb35958892a85ceb4761d4fb5b95cbefc2da5c3fbc09dc42076f18801dc42539df5b7d29824fd469c2d24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f96f244c8f0eddb752fdea161dd356afe52f9ad96a0439ca8b1e720e87588d8044e000732d7f88bf785226e5eaa66851393748d4ea9f0f1930a5ce7693702e068c09ea4a21cbcbb8eb29efbf3bae9ee0f8f7ce48b8a3ecec63e4f299e50cf6853ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a268bb9c9e788e17aae4a6e496af82ea1959aadc49dec13ab37b342ac4e169ecf6611085a8b116ca1e3439080bd6598eab83e2f5a276d8e342685f5f61235111c17389c17172b539a16ca43a5db3c726b341ae0f013a405dc24049b33826ee27ad8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9efb2fe6717feed72a0dcfcd23cd8d16e0f1eacc5b57daeaa3c639c9ecd4c1c3162a52de5b0df64840dadb46d62fbade0fb7004d76d1eeea1a551ea76aee2d1ff1c76b15cd9a2401922f6666f7442cf498eaf307f4e27268a78960b8126a4fbc7e15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2032d886889c4121ff03a32b171027ee54396c82c0167bffb78fc7004ee1618812906830cd6a5690353a8a9142f24e7a3714fe1df7156134476dd91b2c57060043a7d0ae034e0f3ea22617082c523fd62f00d08d727d4e0211967a9a6d354287e3fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88aecda2d66c9963ef4f25cb174fc7168ecd1f40c26f47296929515987cbb2ff610d0d3708db2d898246c36cdfbb3ca6e69acb3502e00e17953675951747ea9425b106d28edad6081e09b307aaae088ba3d94d27f8c26b8018d563d63fb2aac085aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e080bd7f70335e56fb60e17b3b8825ca3ce9130aabe1373604714f7df4295ea1fc220db8248e994665abbce5c451ab422f0ca334846cd97ada9f78a6809346b4a44888864d278e0aff0d9aa8b48669f40e830e6c5aa7d62b57e0adfc4c2963ccd77;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h679c33c0564d9ebe10686a109c8bb67ea40aa24340d80c3c6ea742239e6f284d1106c4c7adba57c72b7fdb5ab1773d988c8af78a569ec4c4b371cc80be84997d28ef7cf644022b098a0454e39fed4808e893550fee2aed42d63b90b92df7b864f2b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64da4ab1cff99f7622b76c85c44352988c3b729b4ec79e23d51983a2c9dabe7e2ac3466ec6c652d7f7ae5c281d7c89b1e25267ea6d8cedfafa4c5d2119bf7eb5f08ebc70ad56e33dc5f2ddc13567bee8dbfee145d6cc1a1a67cedb99e1a5c9a4af9e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5091b5f24cec8da3f059a1920aba495b507436165497f0e6efea3896a53c28b8de23b8e220366b1d68ab8c7514f8bb86d8e47f23cae0488bd9a6250367457c988027ee079e5391c1664ff84b6557895865b4f1cd5f9fe92d2be99953737ccfa0e704;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h966b080f57ac49fd5aa340741ddf216d98405e3ec80f120c4c7f877a8eaa984fa159f881ce0ac3e76bf7ad8b54fce90b5a2b1e7b4c66b9cfc8a20a497da7b23dbee266e6d9918f75a2f48869b90135ff204ddd3af3f86e6e65e77442490ba6abf5ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c54dc02b794510d0979815886b738c0c63f3d6dc49f4c5cf144fc77173c3284497cf55f573c767486443a337dfb28a5b29c26c7210291544df2eadcbe11150ffbc044365e12c4563391ff5db6858517d6ff1764a28fa5f588ef73a4a288da681261;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had78e4dd56c4dfeabde12975cddc2fbf43e1483b8f07cd719e15df9c6b28cabe7cc99b9be8bc9c62ae253fc901991db926ab72667cc8a9f465b2e764ae8bdbc6bc7eb824ceb385b29569433ebc2f59d3d1a466f0e9f65e10fb721ddfd68f588f6e28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h839254bcb274a7ee61517980e39d69b2cc64c18de51ce5a668f4dd4e4886be8a38b9f43419bb2588699f76022174634535f50ae6fca2c0c1006e9d5955177de6c89631fb15e135b1d11ff086539c9880e746fe46aa48048caa731f882488d64b4c6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c8c0dc82ee3902528362de3f14417521e253806370da5cc94624561cc9d37b122eb88efae2866daf07898812250216936181ff6c8d2656938cac26a27db7c363f525a57d7c786f96bc4b65f392b4fcb090b7697347c579ebde5e31571c1de0cc398;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h858f106642bb64b3e3ac8426d6720dfa223f867c3510311d0826e3603097595b610c9f804cb3a13faf31437c141eb39f824644196e700c99cbf9664a42c2058189c5964280573a1bd47938e9821bdbe674a5296bb7c1aea59ed2e38343e3d77ccd2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb605b30e842c961027bb427bacbb0fc7a79c31de8acecb73a7fe0beea544731ec64b96ef251b329451ae56390e35be37aac8605663ffcb41dc75631985d7ede85d6837c2ac27d6aa137dcaba2d352cb1b611a8941153d9bbe327dd5881a9c08a4f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc8c46bb3dab0fbbc4ce19fc735f22947ae8132cc937251bfe64e89bf52331a99d7d792c7b03adf71ef5105bec76a86110f6318ee530b8c65f8d455dd783af6d4a1aa9d7e359496fd35617a3356f170c75b6ea70a0fb23b2863a069163845032b640;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fd3afa2b1bf99328e8761eb2306ebf17f89966154cb05f3101972fbcf74f5084decd579965fd3b31ed4e73d8ee43e94c148aa1b7d18254cce0f4c7015b48e86afadce1fa1edbf7b053291ddde9d8c113a84b500c62bfc3166e6ccede2d95f65b81b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habd8e2c5cad4dbb290fa07988d0e4bb2dfc19916625cfbb9f5f3bb2de3a5f727ed7d98ceab2b7688bb763967a1f31fe098dd8ef3d5ad4cbb2064f3a0fc426bc27cedef8406b0112eb8cab655e3b0a446b3a74f990c117c10e12f5182f322e91e5cbe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9309ff50fc92b1b9b94d104c3ef568dc6582717905decd5809504a02cb8d28132c04888159df8ac73706dded24621cc526034a35443469f9700f95f7f625fb1513e64ee92dff79941343175c8cd228cf0eccf242657934fc061da0673ea2215b2ad4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc1782eb65f7802ca7b4c450bc046f481d25e50a41054df3807142a1ced7d26374b5ffb627b377f977dacee5f305a43a014747321e5f7f800a333e5733e5c62196b1f456f923387e195818f1422e9ad32b98c05086b92e6cb619bc3882a1c064be4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h510282a5315b68a5283bd3341208a0876b87f7ae84270b32e315798bd5eec5e2775d4c7911902b72dbc85a22d93f3cd7821eb87c82771398a4859760e89c20eebf11a3e2d21ffb2c0a3900b113df5545358cb39420b5065f34339a456caa2e854f30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e971000493fb81d214979ab3db108b6b8976ab53979d50f14551c662cd7c1f4f5c4ba96262c881f1aa90405611f5a7d01edc83caa9f4b70117118904f50a1fbf65a0c7082164e40fab64940985b3513ed1393775261342633f75251009e86a3afbd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc871c5b21363868b82107849409105dcd5a37d4fe6249060979b3e436e9e1a1112c489a76e0c157ed2f4d669d126adb8019b37485c9d858561c600ab82a01b438e2e8a1433a8a4b482de845ce5e216b1dac1ba4ca77c3e2113c4c0d8d6c219d8597f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h967be944c3f7c1d738f22aa218f9748bfa6484622a219c7661fdf5499863e5c643ff0e91f013e92b211cf2b32b7cd38bc0ac01fe144e80c7074be32531fe49183b864be7e254439b0c422335874e5fb9393ad7b6184f38aacdcf9ef09177bd188d08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h688838392d852990057fde2ae87f7b7343b86c2ad3b906f413ea2d65c25460963ef0578b52fbad0fa68d4f3dc92c7ba17ec8709dfa6eb3633a2288182283494a654ae07712aac8523870cd9a3d880e358a27ad65d62795e1f8fc74896ca3108e0152;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h547da77c12230e93ecf374c0ca4bb213824c7c7624561fe33731a9e522c95255e1fa5b39a1d57b3efb8cb3f13552e683cbf721eb4e7833b0d1e3db6d260a7167eb9b444242e2eb14ab26c12bfcde17a6997ee3b4d4c46e9bd9ece5901471235db802;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52b4c675ae14f73d31d97018313e50ce28371639dfce87947415d2065de132cb6330c9d50d409d5c24f7e08f96e17e180d4b9249f61d85bd332e492d93792531e72dfe5c167a3e5d24b8e644701fe74289333b3d2dfb8b5b2964e98ac7c21bc89799;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0d79a4d4803722ea42b9ba907f37fdc95eb8837e7053962f73a2c079b56e3929636e2df16fe8fd7a90dea0f0e1feb8246ba0c9ee417860869795e3f3f795724d2bce1884adbdd6d82eec4c7cd7ea144c54c8e568a2abb821b9e46e22ea7031c07af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb11f071a53b174a4010d9cc9733e4d87a425ab3411f4c75629b3f44f144d6cfe8f01ae45a63ab04c5c086630e6e01733a3a7a5b52463dd3cee2e38842941d8b509cd6fefc129cc2ec25d71af3cf001deb9bdd5f396b165fcf2d0d074ae9c9e6d246c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h275ac1b7953effe34807d44e09bf94758446e27ba074a22000ddb6a9a6073f9f5de9c373921441a109728aaf0609f7733178355af5324302f9a9d01370ca40d642e4320a21d18c68645f17201452191ff07f6f43683c9f24897b4167dd7ea2b2b4cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0349a9acd6cffa1b45117e21510b66599ddc2f3c476eaa66fa040913f52a8f5c09f82e21b2963fe5933f066afa68d9f128d349613e467d0ad8ff3753b8a94883bc6f62d5e1b4c6f69940f4af83d2aeeb86a668bf6a9cff7436502dc8da7f506d2c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f813308e38ccf1b4bc2fa084ec8e206bfbdc5c4f6d0158ac4be78d67561825d29a9edf95b2f1db6e72ff3cd20d350405acfbe4a1be865b068d3d441b76b65f08b2bbc77b737b57d8c3788661b9cd364f0089aa8d3561a26c5069d1334e667570538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbefaaa4db66af77ca63890194a7bf166de0ec71defac71ddc35eac98127bbea46ae3a8174d1d75d706640904bc81ee11adbd223e1fb31da0257b703f7f33bb188e47d05b0c46eccae8a6b2a4f5982a8af958018b248488d5d72aaac2aa86d05a100c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdc14f1cf46ed924d3352571293e3d51812e5ccd76deebc3e6b845c606b130309a7739a53733b30bc3981036d64b1a195c2f46d5d48fde95f980c6aee40e1008ed86981fb2adb2943fe982a6f23d5f9cb8c3c5e0feec2301455e68c1752aec41e988;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf34593ad9cf81ac11e230e32914d477743ce70f9081eec4f7251374aaba7709ac019c42d708512f7aecb3598397b54913b1cc33030cdbf78dade4b97e2b955fe05dcd2c8bee41ca4eeccfc9258638f3b9d0777d70be957f272809108e3cd441cfc4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aeccb7c129e8d28baa2d13a41e5a248d5bda4b87e457fdf036ab749fb4e4ad93a8ad5154425ffd705c0c6620dc7ec6f648263b342bbf0dea6157704d32bf5260259a26e831ccae6451e48ccb46f617a8d92bb4ef45b2cd9fad2d14335dbb52df2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h194d0b71608eae77a6c574ad52cfe05c5e640da15dad084f21d6429f61605d9a2be8e45d393c2b50ecb8e0c274426c0de566fe0fea0f3d922bc23b2d987b670f18387cbe786547f78be3259385d562e73e4ba3ddaf03f15ae77cf1dc4a812b8cab46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h458e7c230ca8dad6e28cc25c48e77342bbb1bcd59bb67288923df7cabb46bd8493dc0f9b755cf1d4ca5d18ce7dce32fd41c091b7f3408cabea7c47a2704ad9e8bf57b9351e5f56345dc305b62265dc912d9b8e1e5181576bf4f64e4fecd7ea72bc82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7638d4a8ebcc7088244e509b6d1da17ad5b4dc5a701f27fce5724f13b998da20305d21ac62f2ddfb687fbd032244645c679e896bf5289fa76d1551bc95c617381210a926a022e2a9ef13d67fd1736d7205b60532f5ca597274e6f3133cdf8ea10268;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3561657d3811743e26b145b273996848c6d9580e1b59bb670b94926262a85510d5ebba216865748c12d241aa20ee748be31247054391a9449818e92e2e934c605caa17c2556ec85d3464524502ac2a52f563ab7b77c9424af12487f62a7f5169ce0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb649f43ca77b33d5dc108a915fb2d82671173599a073fdf74a6724ee5597d04dfc3f523a0ff3403f3c8b6bb2287e2b4668f61b3fc77e28197a6c8e3766c864aab7f2dc89997b05308aee4f422830f253bca7c88f046a838e6bfa90cc61c3b77eea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3354fa7c8291690e3755807b5859585ab9cfef61724c632b5ebbd71e780f0f08518efa5fc15912a73c60aced09be76a3119ff7ea5a07769760bf9dd589fd9387cd821dec100d895d3f7e0fa1f612eadd24f2f32e8e4420015e812f2d2b2b8c709e3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h578ea20f61cd5714f6e2eb9267dbfe6ff34ebb817594065a6715a3ba4322bdbf5575bd16fea2435e09db8d6d490880ee523fc8a61f57f79c33185913ba7905e1d53fcd65344f543296bd5ebaa171a21abb05ad5644152740ba032c0ce005ede5be5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4710d732d1edebbddd96c99857b97236d13012878146d058bfd30988089a359f44e963ee6e8e603c1babcf48a69951fb613ae2b8d497d64ccae5e268524848f92ad4ecb68d73021e827c9694558fdb1fe0f2b86d576dc1ad223f0d87f7c80864e0ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2178e4ebf9ca1a37ed457233a02f20b8a60dc45fbb976fd350cfc9c1ea9a1643c1bac3b3d33a6ac6aa428fd9f7113679176aca4ef3b0806d7b4ef074e48d573f5c1ff99190df0ddbb6a0432a5c7a26697e74d5fbfaa9b529ff0b8e162d635784be5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35dbd86c6384ea3c4e4017bf9086a05d4966655a37261a1c0ca1c07ecdbb545ff9eaa10ce83cb4f52ba528963ec1d7011902b9515bead2f773080f233aed17f8e74df0ea3c66bef972a68f395c038a6d1afb308069fd2b5109577a6522ad9e889650;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd004a9512751f0141ab3129ef122e11fd5aa5f34916bfd06c0596813eba778da867e8129f8d25aacf9be3a275193d3b782ec5bb06345a6a1066380edf58faf030efde06c72510463feaec8c2abed0bbaf765d766c69cb20cf5740eadfd77571cdd15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h581e24e497c286a7e6b8aee983a046db1f7e0bee4192ec114f8096730aa2de89ee09d3993e1fb68796baba5e87812cb7657332ff269237b6eb05b91bfaa48d9fd5c969ee51594897fd4d268fa276f741d3fe069cb72321d42e31a8cf97475fb1d1d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he316eebc933cff75b8c84aa74572c5a5ae9f138384660ac90fd75b0ab742456f40623f13f36172f11bdd8c2f38bee2a6fb5e30f8098c86522b6bdd24c789f8055c7ad016b8b11893801147c6e0af81453ecfa6fbddcfc67a035c4564415f8e08f583;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92457ba7811e0699e2c45ce7394bf73f7e75356eca496ccd3040a5bb963bfe0425af354959bac785f0449cb491033caa8e51cb6578ebaec15e7e4145839d57e40fe74781bebfca07ef8bf7206042474f2e57596d538442e5163888e0a8c920dd2f59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1613d062477cb833e4e29d534140a0b72b5a5f3062d68d7c6a703c147a5b956fb594da33d9cd8ab2ba491a6493e16f5bbd27b0619e14cb554015308aa29a9802495baf89dfe70a6d41b0f5d2f7193cf4251b99f21facc98d76b6f99c2b992bee63f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9bc5f69d7f66dc24d816f0aa9fd12c1bdf48d23f2d3f3cb8f4aaa9cfdf749306a9f4757209528e53a6f2b0e3dfeace4a2afbd3d9a45a7ad02e0e28125758556ba817f640b1c2dea066ec2b05f603ed236ada0f6876551a4896d843b98f4e0f7017d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7717c9978d29b54afd17e93736a6a100e7535f62d75a6fa994ae9e1d82140e812fafc3a1624537081ef515439f0f9b31d3076115aa6cd5a3ab0bb2b9dafdb8a4952df4cbe273ec44fdb2f7bde7faa4797a3f08b3cbf8523f3ad35ec5a51a1c0c17db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29183dc19f81a0165c49f49b4612f9c61d9514f4fcdce32d217301061dbcda831eb96f9713658287b5e0304054a366c30a4b4e648059d42e6e1d66741fbdb1a69b755e7f8cd4ec2f37136283fa4713568d79c8ae36ced7818f28a95e19599e366c2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd51a7b5118ec033d5018ba9a19884fe60a160272a678317c6ceb886883019cbc9fbbc3f0a06509ae7c808dd5bca33648c0dbaa9edb644251b74355c9c8a47de3065f2ce04c0828882f3f43bb4f60d77113ef423c795c77a079f56119e907f9266c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10161773d9c8e5b9a7d545ae61bd0e005950bca030d7b5f5fbddf7a3079f8d2574f6518b2fd148609451cd7d6f51e8db247734c8f692970680ef4c2f1bbc4ca4f45f363a0325a8eec0e834bb81c1c5bbe6bef192b60fc55c98ecec749933a9971e92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee5441fcd71095620857b267b52b693d0c6f3ec2d8d4dec59d95f292abf74179962e7d453ff97a84dbab0b1f346329a054a0e44e8d4d9d2e8c8ee4fe5b7d3306d0f0dfee8c0b3153f9b40c69e3de3810d74f5c0973d9efc75ff13130f9a9ee5cfa25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e516ac1035dd228bfa62378f2930b08c75aac94adde0f1cbe79989a50e54f4d183daeb80b8aeefdc6fa2bbc850fd0a4b1888dcf4797e224590f81f606546f2c185d0d4e2ee0810be5fa5aecf570e90ebafdabf9fbfa686c70e48784c71f41a2bf31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb916ae3537dd6bc39e645b5a602e1a40459d00bf7afd7c90c9ea591585f605a0808b2ab26b631fefd1477a1e8b3daf96cd6878a0226dc35db920310dcd54677e37fc784628568bcfdae37e1855cc8c42c4653a440d0a5c834f9083e23ec262443bf7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he724ccb8b1d0f5f8ae143dbc4a3a226bee70cf496f22925531a686478c4ca6153315aca0240e11835cd01c4aba68be2430930a5259e073ee1d8094561a037982f6bce840a21136b6755ad479805794681f73757e6fc01c242dc0546713c8bc97c4c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce0c8e2651cbc1388103542a1348313f38249266fc280f029f88dc115a84455a28b50899d0b36b86fc7f05d89bed582825b6b21534d98f9de1cb2da772dcef1ce354532349b0091ce7f77c74097dfced17adcae6089d0604020e5ae55aaa675aaed2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3c0a66609a6f94ad87e5c74b2a4449aec21e85367debe0fb4c470a02ca3fbb2617fed5ea5c2556be02504bc72394b4010b27742e35c32564d0211f7dd890ebfd2afdeb14e91ea8445a12afd40b3fc3e7c38f14ca5923ea3bf6f05d5f880a8e20613;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedd0e713d99c11ab7c9775f5cc3676f27081859e3e9c6f7a90a2e4b85e609cf8995d71ed800ad808138f4e98880368bb21b6443e1c47d3a8688da4622eb6d68f5b2448f0355967d3aace43a46ae6271f6277ecda615b3c5156382aaa06ddecb6c484;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb96ee69a474349f265d1042fb47a23498576d0fb93ed430a87108f42a49d6619ce8265b9406b7606bf3803abee6c3d60e05a2e005bbc8d695de92df8432acb2424360b01dfeefa331ad6f270ad8990a7470d1bb8639fe3c1de2b1fe01f4891bdeae9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7bc5e258feaa08feb51138fb5cf01f4c03d4b259b25d2d24d30d355608190ffa44d79c45d46dad393ad4252b17c03d4208b922fa8cfbf82ce6c64e698d0401e1afe91ded245a9ba96782d048752ee0681bbe6bc9c69d067ba16cc8ff1b1b8d6f12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f129a8d4fbace699aeb975ba7c227d6e264bd9294a776a8aefc46924b1a1bc4430c34af6eb740e66722f29e28419bc75aede18677e03d1ec7eb2b5dc26d6ed533dc3dfafedb51c16e06e4fdf310b7120f24d9f1a5bc07778970bd5664f918f7dbba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h475426d03d114d86a35a42790bf0954b98060db0089fe86013470c95550c46e4e5a360ce3156bbdad270a4618699d310924e670ce8b2663bbdcba8aa6ff08767f5844bbc297d4a76a69b5bc04e946479ace8456a48cc01dd9594463d46f61608ff76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ca0b5505e3e68cad3acf317cb7de8bfb4734432861dd381a415e260061b787ab101f72a8c3f689e9ea8dfe8738228d05590cffc4b6d4985ea8572cb65d31d0e55c3a865b6b3f19e09d8a57728bb7184c1c058a229bb380972dee446638e8c0956ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3171133baf8dfcfe79116560ad74548c81eb74257bddc78bcd7e50eba85251717040af8db19db26888e95a4126cdc691d1cc61843a94c7e84811732365f7af951ae83edac3302bfa8b16965ba5d485627ff1f8a86ad4f8b2a1c7298e77292085a5c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4467f5e4a140544bd2fd6f72994962de5cbcc2c450ee99be07a099f2b15b190ece0b22b663ac494a1d3f1c754d11c7a7e53fb4f5ed1bc410f7fe72abb58b41d89aeebef537aa3a592b5adab38b8872fb6cf43254b92daf93d00caeacdb4032cf4e55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h339c42272b11df0e2b579af974a2ab1613e90edfd76cf5b28665c81714b7b805309ac6fc9dcdac881820e394cf6ba4bbe06ebfbe0353fa321b537fb96625c9051c4333cbdb62a9acffe11cfcd3747b5ddfe418640235f18462114e68646ac218fdcf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e1a3f64dcd8b79387ad10fbda7b5bc0e670a395e7e398fb01a1eac04c684503de99acdcaf17675296603851e6774bf1ec12c56e4b715835c8c09cfa97deac9a1b2a01ab635a980522f56d2318c7dc43f966238cabf6cacd70d1c4d30bae39c44fd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3f0d32ca7b114f8af3cbc7622e1b0d61deeb78c925e348188b78992b6dfc0f2344678893233fb5c15281f9441f52fefa356f796d0749ade5ac9e24ab3a6dc80db2553f476bea0adccda32c8c295f748c2ec674b152dad5d34b96b89c5a85cb7e41f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb27262950476982bb907daf5acd35a4e6bcaa0b6603f1c2bf469b86eed85244aae919c82f265a02d175d1d13bde3426174f9d3159d48106e42a7fa75ffaedfc75b789a7272db8a222ffd91bdb25b4c2f91640daca83f3d555b1e21ce529d4727f3b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2aa90f35fdb5108bc4e3eb3059eb823718b17f55c401d91e97ed931a2a0852464127f6223d26bed95a6327707045f22bdda1ac8d8d3963e9149a950a96b35dc0532b444f849c8a6cccd6fd2239f22121ddfa375a9c0216a9448e8b830d8011499eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c520fc3e477e69eea2b31940e76ac0a9543afbf9086341ef4858bb1e20a801d114eaaa3f4538dc8642d56a5f22c295dd331013ecf10428074889a58ee7f6ec8514054376a75b28cdf759971cadf91a931dda1c47580d510e45927516bb25217c923;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1e9f7f6665c51e61f20d40be4c52f8d62c51b89d389070179061df82a000a75456f3f7f73fefd14c064724cf87437d3b2da1843d48989ffba26c0cb5991b673e70731c737e4204fc3d8959f1024beaf6940b5beed0b67d80d6de642aed3e747d834;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22305c97cedc448ba72f52012b374b7705d8c4e74bc2e56c8423983f19d11161072298906e9ffb83498efb8b12e3178b09bd7788c910db40975f7f7bf3b6b0c210849630c2243a11082d163a4f49cf0d76c4bbdbd59c4b284da01fe2fe9c0dc27fc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb206caffdd6322c77b7abfbf0e3b228c225406d32caa4a1705eaceffb33f776b67743e8c2152a32af041d320f967b81cbaec159e9d10f01e1856b9253e5458d2bf3719d528c7fda58fc78bcd32572e2057a70722f161a9bf1146f2fa2358d72914b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5edcaf755f25ca7c131cf32e7363965b6225ce386c7ee08f4aedfd24f23e4909b56a6e5e642313ac0c9858cee2f53778d16e516218c3dd21bbf05ebcc05912b5a6a6e3e7cab51bc0e29eae946b51e1f2d8ca594ed3570fd942cea5611ee0443abacb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8dffeca14c46b4ef83c6c5406042264571e14cb5c9202d8ab8f2556cb87e3cb4916df194f4e0eb18beb58b3d61c4c2e00e6cdd784043693dbe7f73a67fc4321f17ef289786a0e994577bde385b4afde3b19622e5eeb189cb9021ead37d2999be3e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f77bcf3a442942cd0a7d7b2d8cd2f2fdd15c26f75e1df2037d7813158738fb2247815d6cd7d366cd2ae9a5fb22aae5830e065fcee8e83cfea5d1b639fc561618091529e155732c69b54a2e16777ce2e7e10863ec21317ac0edde4cd514311462f6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76b1799be55e318eaf9230bb519c01982c7eff38788653bd8287fd9134cfe49071f81ca0f013964169c2a63d760c76e4ae9e0d4a294c3577eb016db502ccac10fc26e83f7fb00d2f84fefc392867bb19331242f6879e4fb02115adeb3e81700029ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12cffc70cb03d33d1e5269919c606ad8c93cd9ade2b34fb9fe6073d872990892bc4d14d019894e2f6ecb27cb0891d0ada2681b5b9e8dcda41299135db9053819227d953053005039514923489563637e32b4a4056b489c58e53a52e9c0a9dbe211f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71a9f7a4a020c3b6dfd234c2b5eaea4762a674bf529a0f41cbc7ca90473b97f7e887bbc021c5a7befd071e65bf48065e57105d45bcb0755345c9680415774aa1ffa09a628687786b7fb223abf7ab906d1b245c3215e95359ea2c4709bcf970d5ec87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h500ecc6bbafd5b42f5988211acb9c45fa3a1c550d11ab632b7497b935beec46b47677a6802b8fb072f3d391f07353c5819451979d7c507b73e2f87581e3fe30be8dd7e0ac5a7055faca8d4fc853bcccf21bb8eaddc733969733b1dbc6666a44bc049;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h742b6c8838d861a6700dc33643382c0ba9bd7adc878ba2075b77001be2acb1c00a3ec2f552b08af1123fbc5994d15bd08309bace8aa10343ff26f43172ce5c0c2977ce71522466bb5b8b58430f61af479838dc454f5f81d148fc30b37026af4cb50c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22eafce9764e4fe2d8126575c88b7c712af726d364779dc3c480ae33fb400b1a24051c7aa3cc7e20e064863fb9f93c7dca5e2d88423aef7ebfb2db972ba2d2cf0c41bc436cd46b52309c0eeaa5d7aec4ce3019e4a888361e51e300ad42ff240f9dda;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92e21eb4a6d9d24819ff7c4b56b75d53b69e82bf2a6415e4ca44adc4e564e2f78110774469efe00b4dd8478cf474c69a29ed28fd52aa3d3993b8dbba6b330ea965080248f94fbcff85efe45576d096fec087246baab5833e18cdc7024b58b92ab999;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8358eeaa9b8271f836d4d808c6481f4941304c277f28602148a0de1faed6c2a905e088a2ee4f5866bd5bda046d588964653f85ee507a742f3632b149689f31cdc8dc48af853824916b736bb5aff874df1acfe8f22a0a8679da1bca8c2b905352b5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20e101e11ac864bc0f089d04ef4412b0ce78d1f94ea3120cd8bd201ecfaecf6a55522cef4dd76462c5ef6bb8c74e34d5913c0812bbeee623f2fd6153fc73ff069fe8d28debafaa87520fe7ef3cff2787ad3fc886e2cd915fd4e6e7072d16f8fa743a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98a895d25ba5e9084fb5f07148b6e43bb36b7cde30be9832efa0cbf6a10814320e08850c1d5d4945118251e0e228abff0d03d830640bd8182854b9c63f3e61cfc5c080b6af16a1b1e64eebec25f450891532bb43573094972eb38a865aa99a70cd15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28f693ad01147f52bcd27b4a0192d6cec30d9c2e8a75b28e30bd8cc712c444c87c1ffeac9f17d27c3af60fd9207780cbe73d0d970744a829836fa02e4b3e98358e7424cfd37090f2b359d1987147f5dfeb01d44b812bc770f2d8cb8723ef70dd48dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8b322a663f5826538e635808755f07ff3339e7c01146b33519b376c8c9bd4cfccd5d1fa7870118299dc6be90dd5c3bf034682c6ca60e247451daf483cad4dab1ebe029f9781d53e17d2dea2ee7a5c2011116d016b402bf165ed9692884e0af51795;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d65fb52635adaada25a892c27a1e630fae8fd2bf6eacd9027d267ded64931b8294be7c37f4db6fd2998763dc54644c0b151a16142d37a1567ffcdb5280464e0661bb5ffb0166d31ec41693016ada30cbdf1e60cd4d0656f31999d7d41702daf807d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fab31ad12d7c7649c9679643d95dbd45f6d1f7c61529fc280d14e8bff23db4813c18585527c043ea0d0e578528cf02e2389f038ef811365f5abac1afe0ec6e94b03a3e6535a95d3e53f106538495f929ccba39e81611d63885b562b165ab9a114a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf9c05a0ebd9b0a9b1c9e429abfe8b642b7b79b7cea80132b24706305ec6365188c8dd53431c0969a992a3a414787cbf544a288f45a920ca3eab7b3d15e3964c96dde7c40ab3a844130d8c07291f4d43eca92e01873fc15c10c0d781230f9d48a86e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5bdc6d7e63f75f8db24af84cd02bd794f1e2ca4acc7c35daf52cde631078417c04caf9528ce1b102dfc2efb8af4181c72f80f6c6dddd6efbc99ac452ffdd28d72ba9c03e048d74122646e51f3a1e7d2ba0f03148da4d30343f9ddfa18d6ae408fd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2af4c3a086908fd5d8abcca2b50d7fafe8c725b014c8eeb712773f93c2a0efa0554e3be964a4208155b241457b17021feb7c5f8671133fcd09b8a2e31d1a36f358226b31c6dbc42e08245fb5ee5538418274dad0c3830785e0853bc9aefeb5d008ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e986007e4400e54428a85ead0c3ee9cec84a0d005ce5a8d2a674a4ec37eb0eceea70bad85d64c2d000a98cf67064a576f3985be575b6ba728e2c104a130b7e702dc716e9bae9087afc9a3b20e65de4532abad8de9c4ca0c6c8558224d91bd8a12fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a4a71306aa4b1ce95de2f43dfba91439927ef377f2c75dc1fbed437cce2368ad52c71229aae77ba98399461286187e625de773dc14c8f9f96286c9432b4f640f712195d3a69514717a55f851a2c8cbca310853e672762418427c59272fbb986217b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68a7cd7b94602067489e4d435842c7d98fec2f24071e81611bc97017e8e20f26be6debc2ecd2502d565d860cdcad20f467e9e5a5152159b532f0dd72ca7f4132e9dc762bb763401db20973876dc60c7cf30381fc0bcb5f4b8bf86f345940dbcf24a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67835043c89a4331c5426a2e5c70d89defbffa1868dfa9047bde4786425623b699bdb60bb3abcac6e6bbb3b40a0e29d89332cfd900b187d72556a4b62a03c96a567616157b8e60b71889c4294ef96d6b3ded74d63d0351dfb41fc76f1e5d2f95c46d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a6f74ae4c90b801cf420f128a2b39e6617932e15da6582c11463a73a58014baec33f72fa775f8c9141c4068019e9ac71e18199da63aaa94b82fddfe20c0b5bc17d7ce10067a0cffaa525224c9bef11f30d89b6b7f441c5d36d59023ed489597edfc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfa86235e95a420307ff2ab75606dcc86c3d9cc7dead58392d648b8e9e08967a43365c4e3a10d62708be52bca87977a8dbe9ad3e60d89ade0c74c9237c816f6999563d502ecfb05fc73a19b45598cae4c8a689674ad1a3f5eb7bbc90f9f2d2ec1e95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83843e618a353d329b99298175c01b6bcdd28a22b674c3dc80371a2ae1a07787d82a595b544d852d4a9a4de922ed61df83ba73c43b232cb069ca49ab38f3073204c88d3515365551abda4a31d2edc22fa8aa5ef845d7fe8fa99e4ef4fcc1a564be7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6030daf6a9fc6071d3f9390d57113fe88ad3f6914b7dd6083053f34dab873ce8bedf91eced6b846fddce45518aa15cd5ac76ac3fc61ccfbcaf8731078e615c38396e2917a268fcae8ff07a283b4a4a2bd0234c317f47b47c62b96b8e32d4f97d2d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6adbd96064f98884a2ffdccb9bce0e765bf7ec038a22337419ecfcc8b8f2d87c55a07f4d3d6896cd0b0f20a7806b46ba0649dc29818370db73bbc610e57dcc77b6f796651319eaa911c071d767d883934b2c5fc92c8d107e121e0e5f945f3a742e8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7bfbdf3f1113c38933acc1f4cc22c1ea38614f79ae48c720184fc1a56886194cb970e5a51573c201c6092d8a4d28f6cddcfa91269026cb423465285884f4644201c563fa44558143463bc78b0abd79fa8e6c164770f6e299896c09623ec426582a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1483462a6cbc2e05f8736662cc42f3b59b0e7308822dca21c20c7054f68f69dbeefc242414a911e550bb302bc101d984e92dbbec8ae771909f067b1183cd56cfcdd84e88345352cdb1d5e6e8077ae1d172ba8b50e7975da060ec2ee98d2a8f6b1d1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h484c4d48961698d884f8bf2b0456994421f350cda1389efb2f59c01e74f659613e7199ba624bdac8e8216b193554bb8f75588131c476f7ec1eee56d08f6d2235d7183ad4b17e11311d81630d6c2c3373e3726057759b5e6d1b5a060eb550c973eb55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58020c46d9ba6649e929e53748af0eee783d211ea0b9b7a39684e02fb17a1d892b0af7561fb001aa2f4d2a566dc0d089717cfc93aca763bb7da4e996a20bb4a22995a4a6b03125384abc4224d913d5e9576706a37e6e55b392af4cfc26f11d0bec74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e09bfdd6577d4e1099d16f763a5f88fa3b8df7ce536aff742d95e1f6a2da6ec15120ef51d01d812e5c9237570466562e4921d08a15cb2b1a749f4c056d35d94b76acd5083bb1af9141b8a04652362e442c1b3048cf5dd5b41a60cbf7109bd73e9f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca54f21608d328bc90dc79435c727eae0157b7cad4a52aa5da1a12dfe3253d310ec2d5b05b3134135f8fbd41fd3cdf9501c084feb86378c8d30625fd0eefb7ec1776fe85cd953b3751930be6d9097e18f28a5a4b0581830199003d6da3385b22af0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61711c7c05f4cfbd7c8bd14b5abd339d8278e19673775f0d719ce7a11c75363ca4469502ac0b7664f9f20ea4d8867583e157201d442f10e9731e84e72ada5843da0a1248d06580174a0442a84a5e897fe85e2066da58ee4baf528584c92ceae66ab8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d2b307724a360cf64f5c5c5d8083707fb29351b10e961cdb3198fa2b9e37337e2585d0e6df5a9a96fec45c1eec886528b35c398428dce995c5e63d54d543e60362ba68386dafedc59c236ea54c1440bb25d1b9c8025ce1edd7a5e1fbc23710fd810;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1706c65c963d49df52facbaf254ae49ac19abdfe519739951fe755191b4e18fd5c69a7081e0b7df66acec4d7f6adebc463d573392f808b2a733f9df06b51f6006276f96dbedf042bae0217e5868a9a9c93b48967d52ad68ab95cd06c59a58ff10209;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca0c66e96e02ba25554f30b570dca40f9a3be5c3400bc878489e4282753ae14d89ae3531e06d0a128279322a94b86bc1d40a72088e0de66bf19c27b68447fc187ee104dd4f49b743388d2fe832fc01b4dd238e7ac363dec2ac2c1321df5313893d56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ac6b35bcdff91294ea7f3349f1a9bf79c1b9065e349775593cdb116bb929f418cd06db31ecf53cdfdb1ef0e4be0c4fd10022afdc0a2dd5f3e8e2f4d76c12845594ca5211e4c6d137cc0cc00099edc1e83f120685a75e303cf26b90e4da2a4557422;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26011f10478f84ca01f9147fc666c57d4e4d2e9d95674a428caa175ecaca6c6f9f64ae26614a8537a8b42c9efa65b8bacee305d0f2d376050b9d1634e4bbc5760346f95ab30506e71586f98832a7e0c7d4256600047214735a3b015fb29785a1f2a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16336fc5d5ca479539ca2bdf1a4ca377b0497257574fb97965475c0e7aa5ab1187437b0168ba3c57dc827b05397c160e7975407265eeef1fface4a443df31fefc0ffd42ddd95eed31dfefcdc3f5895121af7b7ef4b95a72ffc2116ed2dfbc5e443b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h706dbf21700bb017187db9636994322ae527f348d49c193a36e3b7b2b31839e759892ba8182ce12df27f031aa1870d42ec940071c98da6c2842b9cfcbb18d56da2285ca200ab9f0a3767a5ae0b1a77b91a0e06862ff1e0d9f64e7fb975e04f83e176;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf01c387834d2578f09284908ce4a718756a38bc0132e21553ccb2ebc409adbf4440d8fb785a739220ab875797ca5041dffd25177d7bd3e761e6caef9b2d3a77acda70d3705018fc0fc569421dcd85241cd334c4b49c639b22e5d1b955676d6da7fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc0118ac868ba5476a6337f7b8f0746550dc1b578059de0f689355d5ccf77a9ef3fce00ef97c22a85ee51445ded32087ab932483df3f7e119a0c61ddaca06983ebb5230d06cd7bba92f2fa1bf86f2fe8128214e28472434438cdad18225989b9a865;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc19cf975537ace77a111a6c021262bebb2cef246c363e2f51bf96747584790e10348422c33d8b90c1169f441db359b19b7b369cc7c2fb00460a8eb1594fbd9cffae76b053617693f163cb47181ee675ed6b911c103e5aedc58dcaaf03a7778ca6252;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb30ab5931d9da831ef8cec00b220093ce2e99a3f71866f516f3b776e4e054b990dcb16d599dd1970e6da3f0bd8ba597a5987cc378436818c3f2861e2e93104f091da6328b8d3edde21f73604e9236eb0ce7898e6a8a97b5b78e7ca3624a4d3d7ded;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b404a7dadd54e839a6255a9e01ca0df7031e9893ebfa91ed29cd0abbd90947d18ea7b3f860c317fd00d68e8581f6875481049f25011830056f60499c46bccf296030db18a241b3bc6e382e92f4505b95b390923d0041ffe19b29d5869ae38740fb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75ebec08f8d3f2e6b33c0f4d8f885dc647b7e4457d90a0d325b246c4b1242a7a64cb539eb8109847226bc535bc8bbbb88006826e81e402e4a4dbd9f12185ea1af50364e72e1ce6a5472fbf93a8d08012bc389cf20024be974741c730be356a70048f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf418dd9ef6ebe56b41d89be7c005b3df1a4718ab9c76aaaba18ad87a83cf43a08e0f6b3952b7bae482eb200e7316c7ec5f8b896698ba1c50db09c14065778a1f7ce618eaecd63737b55eeaea951ea68091e511708cbc0e6c322396c22de1e69d444e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23dd04ba2fc290d11edd9ea6ee5f692811e411c91c0f466d15e50cedf71ab10c8dbfa8eca21cdc7c95ef43dcbad2a9dd14e1c61d6b58fcd1a927a93fb8b65e1f6ab78a2c7c3acabe70f64ae4a4312fb739016646db2fb488da9bd8d005e632fa09bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3650d607a129d28ea0350f162bd2fec8689efb97c3c50be67a91056fbff2d9c3bf3f841ec10430238da3a00699a5cece81dbbb887f8ea6b9bb3b6cf4f8a4a3cf9d8905deb19a304cc036d1c24d1c46f477230a1c084ad71f5af206dcc3446b31ec5f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbcc545ccaf3d37008815f91d8457d1cd75a281689554fa727898254bd865bf57c0433ee25da83e14e9923afcce42055c3380b5b05ffcd2640cda2693eac3a78a944eeeda366f9c275af6b7f62ded2b43cfaf66f534ab3ccc39810339be0e8f70636;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc296da99f263249b4bf0e355cbb020886ab041352733cb69e7c8dd1292a16ef9b866414a353d1e1442ed098c496444d1de69f22d0c592cdba266b8f2861c28633bd0fd1648688e363478e9710f90cb910d1a3beea6bfdbd01478e9bd7b0af65520f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h970e0efdf76d6f41466f2c9922edef90c45fa6f4a1d01b199e8ce676553a3552782fb3566471f43795280f8e2cbe11cbcf6b1be0b6117e344307cab6aa7b3f2b250d292572e9864ec6e38e4b67eff20e4632a8a2231d59d08e0685c274b84e111a9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7681a96debc2a7b58251c87a244ee7ae75958b937bcd71111b4a83870f88f3212446cb55303e21a2015e4d648951abcd594c784f082943f9e55230b26674ee1ace6aa71c481ddf160b24c53d0e51d7333396a2f08ecb0adabdd24ce759a27c330659;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0bb49b8dfbc9d92b2cbd85aaea913cea434f63da5c648649c00fd5fbd9ab0236847e2a5719461d2744b1a66e9c799a39b1a73aa01bc71f415b18d8024127d721c36e2fd25d1ce3eb5f2f1e699860a80c0a16f4f4ae794d5a9eb27b2041db1ab263a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h571b6c229c3123a24941e9d4f12d7482eac9fdb91eec69c87c8a3f25c4d762c3f0aa4df5bb322f6176f821da12abe964ce048ac04853cd1f967e25bd6752c660ac2b23e37bb88c18fdd9481ef4e1b9dd2ed9ad3fbb3e3660e50a5226d076a8a2af8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8a2e05667b80c9a7fbbf2a03be001822c4bbcd7e4a965eec1839abff925ddf122bd910da3433fda0755c02a890b2875ac3e3ecb9f36cd1891c7025d60411993d78f4db911bc6d825e8e38cf46eb7f7b9bb36ad19543d382a510ae99216f98898853;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd78168bed729288ee31bfab2b31c1ac3d36b49b7417b71f0e56c728c1daa486596f8a643539b23659731949d48ccb662c3328a86a04134808fe5a39f3455fd63ad4b92cd11eca9620c8393ad81e6ff28eeaef392e8e6ffef4d84ecc4ef05445cb95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h552701ed5e0dfef74a6c17ce032619afcc7fa11ce07fbdb62fbe6ba78e5400386e83f469fd6c0dca3640ee61446d4c03157343973131ff0d63f7f17fd9f948bd3ffb0faa61cef788b7b316dd52e2e12c8d685015f21afc5436b01c152205afb79952;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f1fbeeb0081b43e32b120dbbe0944261a241ecb9c0470c43429ccc91e38263e2f46933819c0cda776ac0d38a6821cde63830ec2add9d97c5ab7301b7c8e602271bc3df57fbe2786ec31d4f092591799491d48d86483cc5e4c7801166f983779bf5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97ab5ba21430e8aa39e0bb5756b8af3b631805f839dc792a02028436477af895bc67703aad341ba83a023e9f5cdbcb3f806790a92569c1142a9d8c021019167cef63b8d9019336dd99351f2d90716bbca2ec23487e5056ce9a9dde9dc311b632f764;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c8a45d4c2e63e71b83e3997c8b80da62eae1835341f8a37089baf29db1878c2b92ea51ce47de9a06bfd22dce45f4532c9133e7d36a6945451b965f6772730f03b55cba08fa2caa574bcf390922a05bdde37ad880fc4257988d70820f559a0396778;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82b193839cf4002fb63ba48dd1a4d2fa35accba8e9126006806f52feefa3488ba260dd3f66ce90e53e980822e3cd31df7e523adfe0c79bf0162285a4e2f0700231c47131f875992d9c2d635a26c477dd70e2466db29c51119e0ec93907bf27d02aa6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cebc6f85ce7e0dc148911d38e5fe05a83b9de7913e7ef79866d3af890e147e90f54bdb78cba7c105013a18d1c52fd2449994477fdd861c9ae09eda1a8f99a9dedcfa42afffa7981259754a2852a6cd4ea0fcb071ed92090fe61c225ee4df0a3f5a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0a1a6a3550b40d93f415c37de5d1d3eb6458ff85d1f3a5b4d8a8b98ecd013277d35ec521b62f241f79be5ce9f61543e268f6f8fb0515c9f73f085e49f281a9925c4e42b10b6977e70f2c1d3bb36f51ba3de313beb75dee43061db402b193712d8e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f7a7167477d665c72d9ea01efc07350f6a6673113f85438d3b3c47c0da4973db70a804a9eccc5c7defb7a358eafb2b06abbbaea323d01432fd77b8664ad19f92306b74d0729355be1a97c97bd6804d488b8bbe04bb38da76bbfc90e9ec768986f64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70d360811af89a8013fe929daef76315fd1837bf3ea6e4c49483e8d59b82949834171eee204e6cef112d5d1838cab1b2f3d4ec2baebd880f7210ce443bc5ee24552d1c4ee31674aa0effd2499b6581cbc3298b53d3e49dcb15647cef6b853f32f369;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87f21e91472f447a8e3b334bd23e9d10f263212ca7b81c383a14038c863cdfd8779d33ff4d88c2b3b6f14969ce311b634633b3e3a747aa0aae843630f6cdcf2563ab5d7b1d026caae80902f1104d925c7d34997c6721283c6a52e37b30edce4f8083;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h279f0c7f267410804c748a762bbe47a4655c32c130335612e0abcaaf18ef019c9d978c583f2e10f1efa85cd475d84cf1ebb043246553a215cc320f1d884277f66d9f2a877c67ed22ccc9b74fe52cc1da293323b2a0d4bccbb078fbae6dab3e20eecf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae67398be4ad2ff1218c5338fc54cdee4eb09a15af35ae61cab4399f048946a3b99186edc0150ac0e0c0b85ca8399f6d09c5205763f0847c3cf692e0a604ed1498f8b9f0b809afd13be1f82ea31cda1d18f9d6945bb8e992cc5d060f897cb9ac6cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d91946975c5b2a70c41a9de65a12d0a9274653bcfae41a2c1e8c4e691d608334f3c64201ed12e499ad866128626b5ec8f0991e22b874ebd67d085e00e0c1516cf0a57f3ad8870fad8aaac33b4e03202861c262e73ac77e3d229e9fb6c4382c2e5b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc475fa231b92392a6f4d7613e2d24e5056b8571b7027a7baff51a7a67d7ccbb88f6ecdd06b71e950a599aacb4f344f975b9d170547c69ab027e64cd716a90387e14d070ffb42e249061fa1a57f6bad6098e01935c09f898e163a9e1fdffb9331991;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3948e2a7f410478d1b2396b34b8d17985eabce5810f8a97a8f26aad653059cc109a2ec0bc0a9c8e80ffbb4fd2a475c72b60f168239f1cb648cd3ea2d18d96e1c31ae079151dc11272bfcfb1e35f59d6b0ac95a996d5656d7c10efbc0ad242c852a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h647d0fb21b734906a655caa95988360d6de8259508a71c71616e0431080c5a463d5597f27d56d9b23b01721aa90547b60e6704d0c5f1b64366ddb49064d40238caf5f73c61c32500a29fb5aa5b36bbca85ceba78c5595970e572f1de1ebb3f165a11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha866835d91efd89b5988ad9e16b12f7fa7e60af79b68f1d676fd383a85afac99d1f312a3d4262c5d4e49e704f142344e73f870f110a437822f3f7f55e734eb4ec321318544e68b4343ae647afc2c77c889e0d1bba0f15ffc86e5802caf29e4d2a336;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7c8b41e9a06bd903ece1b7ffc01f313f063677674c8c98d0f2fd7cfa5b5980781b318a5d30110527364cbdbb9a89a411fc495e3e6c497c80582e01144597f8b11b700b895a0e0427fa14848593e95099748b2463fb0633704a0cc4857eb609d0d2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h150748f446e191756f223ad63b660cd1c1920f4c1733d7782d87ebb739d3b170703c5a9ab31d194a1e8c4ed8a0eb9aefabc3923e7d981e56fce8689d5e72a040d5dfc13c28a4c2a7e528373fc11ee3c4e8376d931feb76790769204f0b46627c4c52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34e24350071364d1004d65ab1c15d64c02b2888d0f07737dd63f8afee76082beef2d6d1220ca74e0d92e3f8a1752b6e6a4c8fb43d76bbec1e4b183b0fd99fb6055b0860dc3f84abb823a52765a7a48aabc17c8571ddafbf8993a363c06e700e12909;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3710fa4b95d87a6a11d604eaf6f6a2ca0c62676fc69911eaa3f78b9a0a611fb7e4f83605dbc21a0e9f9759b3914eaf57feecd51969d9107f5ae9028e52cc1fa5ccbbd1549b4e300fc51226e224710fc36a32720ce4b5d573f7efb4200e8eed4b751b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6f97183701f4505071feef72ba911d7d2b3b05bfe0352683d7707ee911f7f60355bc080f80861214c03ff0c4c595988032ff3971bd93013855b6f4f9ca64e40601638a2221b61a65c8a0dbeb0ecdc69549e3c37d4c0bc2a4f47010d9a1592621595;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc01bdf5f00455e36f5469330de3847a6bab110346f2cb7544cee4db0a90557458ad556abe39d343f09bc3c6cc4d099131025c628d53d5400aa0232a4e6d14c6849cf6653d8b50636943ddb1b012c3f640443d6bd8e6f82d5f36008ded5e3f1d5073d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7753e049f40554a41366940108376efa1e77d1b97fdf8091dbef38543046ad4ba8713ff5f9cf7feebcaa38ea89ac883fe5d32d26e0adc53bc1be34ae7291dc35dbc526319ca46aad7db6185178d488459fbe20f14a607734c30a835795da8893c550;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc76dfa747de05b435b52ca27fb21c0aef1cae1786072728c0c6ea568af4c90aa9d591293649f9f3dbce5875021f9339db2434ca13bbac2b65cb38bbe91a4799500dce3e87574d9003742cb0262783c92d81e8c196febfba6d88f08caf2e4396c31e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6d94e1609289e3dab35d66a5e43e2c0b5f58c1290221d3ced9d27bfe5890a7564d61fa17e8efee0e0988add32d8639dd84c7c9c83e0e1dc8ac894d56d1f9b083b30306d2118f042b77438f2f2d87e781ba4bc3c2e549c7b4bfc5a9d6f37076dbc31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcff9e4daf6a78cf2692ef8c6a9fb11636db83885977429059deb69c7a4eb6cd520e2a4a927e96cb46cd8761686b04d20c7becc4233e58ac890188631e10caa2320930df31e7280ed784be42ed1166d0143f2e4aee81acc5cc617fccf9cbb3b576292;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5de41cb8a0ba0f84eb4bfd16a2f70088047718a4bf9fe8ccecd44c135660de46336d8b4526827ee7d93e1f2b3c9996b6ac96e2046fd0cb79f40b74a925b0dcc5df45c163ed8d27e5ba24565317995d53ff7ffd0638b56fe1e46e61eccd9511dd3259;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b512bac8ec2b02dd962c8d1b6de9fa2682fc3f19eb2a57bcd9187be64fcefc6da2b5add075300920f2ba925d34704f412d54a7bbbd4a9bc5b934706fa24943525a0bc6c275be3e8b63d980390a2e5fe0a7fc182ee98da2611ae55ceef89df1f1e8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf15f278447546982a7702ddb8856a20bd9adeed82585a5df06c8317fe019065d589f12153df143386d1249e425f88c7307e9b70ce0774ae2f0372992704cb38bd28475e9121382faa51d55c3cc8649cec081eeb6f1aa2b9be4bf07352fc998652f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bd2460db9fd607baa2a606363dfbc3dfd22943363f410f801f3a903cf2af016ab325f40978b63d2868b3d67d34fd0a0352d8ac7f8a2dbcd1ebbfe0a5b301482f97dae069f13b8adc3b8d96c75590a663ddb9167a1bc21e26212aba22bc4e2deb4d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dccf075fde9fc858aa4d52a058c1debb72734e3d91a01bcd7972a64da2f49d8566400278bbb862e72472585ef122599e78d38a0be9b3a3707b7d132ca7c5668f672f44df1322faf9aa477a0934c0e1015a903a828ae511a71fe47cea20a7e7d489d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc087e5871ac157283df7976b1b58ec75a8c159fd6c4e904e9731172bb4dbba8f37df9f3f058fb55704fb8751ed1b8af00f1423dc5ae31aaa24b8fc73ac26d5baf647a0b1232a79de68090b9c93a2b65e50b6e9f6f8363ea174dca09d9e29057bad9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3fad6b9ea9969dfae5be07eeaf2e24fa902a17a7ee94ba68c9cdd711a57378c293b8eead10c6fbc5dfa626d924b36848c19308c59ae63883b510e68ecae48ffa1bdf6a88fc2193d59142f73f8103a315c831eb50c4c9a22d48927ba52e73b0f048b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dc2705b0fe34d190cc760d3afcea66774d3e3ec6768e2f43c28329b574e193293ae098fabacda93697420d9848d5c4665b5f130f4c6320b01c4870cae4851379a53fb1b6d1b9c6f99b35db57737e7a54f85c5d7d0c4efb990fa16642eb672d5a9a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2186a39831ad069cceab9e9ba735b97cbbf32890d80c4c630c0dc091dd528658b8d38625841bcd67c8c94ee3008abbf775219643bfc155d4888230de2044a9de598263e29f014de39b541ef8ff69eea0e5f87f64f2fe73fb5e1550415a8a79db0c26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fa8ceca15dd4989a0ddc04a0a60cb8ec3eb680a96686d2542875a08d206d02c4d684d4c7d9d1dab6960ad3e8dd85872eb9a13dfd0aa5143d8d729422ddfa9952e39454ca827e9c529c8994848826607f40dcc7a42670394bb96cff985a5890e2bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f71635fc51bbdc889ca23f655d6f1c294cf11ba639e5332a35caf53f36c63f00f7efbc5cd15cede4ee5a553311751007d811f44aec0ee61d2ab1925492904b2490a9117db9f440063afb31b77f5c38573824cee6d738e61e82323f7d43799155d09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hced1484e87200aabe60fe2814d9f8e099c7e8bc2349e320831e33e9744f975f12d75a5cf8d27a08161b3032517ac36e748b097dcea19dab5079d26b373b793010a4e12fce27a6df6e8bfea8ffe45924a66ab080a08454ae9982b9dbf83d1e4a1c912;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5647d6e0778426f4aa7e0065ff38ca7b4574476fa5b462a5f1a041fe05bb07c7335f83fa8a64b18c40375b4142b0421fba7af1db2323e626b8a5e9f62bb7b2422b89d9e8d5e26bfe9612fdf20d2385cc6bb12cc5aef7761f9211854b08de691a991;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12a1c6cab25d857896300895e2abf25d6fbf9dab8677818716e9b81c416fa56040662c5514ae5d616191f76704a196994ea7d27ad35b7b75e137e8c4edc9d6031b9f6232812d7b9ee19dc5ebc4eb550ee8f4b82a23bd0735381399573449934a6b83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0be0e08d104de86a47af4ceabcb5b783029408b857286e2204236f1efb5d525d9243a272473a3540a60c55495cce860fe134b4351a243a9f78a8be15d13ee14b0d0a6acdee9bd9e919531330b42a7cf7c240784929db464613bc8b137c6cc5d048;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7875b499e8d0aa366ac9f5c3a331c53ea60d103e2df02610c5c64f92c78df816ac4a9bb555dfc97d2fd2490c5286fcdeedd786ed99d0953af13980471a2bd5c1af080dda8d94d69815afc6b9cb29ca23f1768c48e16490191019aa8f0b5c51824225;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb954cf422d9c7ebe85eeafa93bd43acc73151adbf2c1ef25597cd1e4384f35250501e4176e29c5178c85451bc1b3f3e7e8c80deea233e16c44bf995ccdac17b64ddbc4c772563379d0b1283bb5d1d302b31e4ddab8bb0211e179154d0e6f531a0578;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29cc6f708897161c0fde02111a11937448a61f664301645692cba317a3eed1de0caad34b745677fd072fef7371bc1c1a0884ec459d800e34a3f7cff055b1b4ea37e2522956205f7ca07f1418501d4042a8f2ef174db04d7593cfbd5ebd23721af8b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e511f974cd3fe4398913861b09584fd01339c8b9f83b325ef771b60cf37d1020152183842fae3f176cf5cc2be4eeda00de94011c52572587499a98af06ce38cefc9ef7a2c93d69dd5e83e826be201f600d4362ba3d9d40a5c14f6cac4a70374f1bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaaf35c42278c663e9c1485f227e1b94d327a9eaa03a2a97196728cfa9d8371bc7aab8684c82fd7a9c209184eebc7cd8e0e5888c7e0ca330500187570cca11a4c7aaa4a2806ea1057d8d7b5daa14cf126f6475fd321a6af5566550f5934854e9bb60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b9f90fdd77b751084f2113704e2692da9d6e794d36f001aa7aee3b46d9a2c7087824e221c1ad4a9faaac479a0703513169dd187112f12e87af3087699f01d93d5dfdeabb58bb048d8bb40eb52149eff3b531440571c104b38742fd84ea8dcd5f732;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb12b2dd221b8fec7ca0c86235a2e8a916bd738cbd1b72e6301481e6e44b87bedd5fa47cbbe6af96de7d98e730604345116c7a032ba26cd92b19338aeb0f93209e29fb8e5c556155c39741800d0e62fd1e3a063ecccc16f5a48b28be589c47f6bcd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37d14393c4eea07890cdfde89a1c1e5d6292058c6f23dfdd4bdf43eced346a8853e95794bbadedf2d5b52043df2fb01ad9e1e2c642b79c8624bf9175e847fdf634a15ca1a233eecfccca8c53cccd9852e17e2644bc70c5b551e876a8fab9c7514ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3292bee12c04283a1c4a813041797082270bdf9007390d71f5e3d87ada060ee636ab9250be898c4fbbdeb3693f1898be1aa2dde93d3da62fb02df633d49cbf7e140f5633dfed6ef05e56d13f9606f7febf0597556c415225986a762a9114239b52bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac16327f578d29fe6fdf2e855e1d6e4e3ca1475f2b015b1aad981b0715773e83e5209d4327431dbfc3b21025d0b704aa473135f7558d83eedf109e5d4c9327ca3cb16e49442949e804b97f41837227eec16844da8fff43590465e3b0da0638d58210;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59f25b1afa990386d74f748ce7f6123606ad8fe2c379418004a51cb97f4c5a2d8ca5a4c3d0b742303e285116705770daf9fef73a2df6da019b996326ad41a4d5e6327ca10e356547c5ceafc67adf8af065a593f81f99f3d30c2ec9870f74b4eb618b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd88dc0bdf8be040dad52e5c87d623dc4d9ce63686d577abc05f30ee639076cae8d2f25052e58e1f9c1cf6fa3a9225bdf1a2d060274b0839dfbfdfafbd31c6e1bc90dd7564a79f0a1fd38dd8ecb3fad4365053238611fb17cb455478ed73007e6f7db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha75cb939200e981d8df8eac6be67f177d6bd6ff2c2094dd79cc0541ee7952a32b38816faabf0336c322becaaad933c55bcaa12a85549da381b433f5121395603644577289aaae94bf31857cccc155690a6a157f29247ea36404a6b4fa2aa0b1366ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h270f33807178ac75b81d8f9f20549902ac72b1b76298cce0060c4c5c0568bad40f4e6254617e6be255cd8ef3fa0eccb1a0e6e27eeeab5e3d458d69f84784ca9e68d99db8b9aa4db237da5639d7db43ff379ce06741f767b1247187d81c9f9f07c0b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb5629e784e8cc1fef003e7cb10ea3605c406b25fdecae33dc4e7d10d585c5bc1d05b4c61e36976ebfebc4b2c444211929d77aff49a1ba113979da4be0e89eef6c58a2c4d1888326bdbb25f8ded210694bd5e30e554dada91d91299188556795077;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5828e961add49a453358e61fe4bc21197810a82a4c43ccdd152cb9bca38c57846ec26fd509a3097b7e40f9cd9ec5028e7833da0b3df482dc60c161e4303e8b7263c1567edb9cd46575dddd476f43463296c42160f31882fb3e74ab6bcc8156f76cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f60c87a039d7e71ed23c9c77243792f877b830e202cc842917d272ec444952c707691a27ff3daa9879f6b76a767fd07a83cfb193c6e5c047b5f1a399046eb3dceaaed49db0c97e9ef824422d4d173caf37f068b25ad5b8e42a1d88376e98bd1898e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f0c18ea339549da224c8f79d092315eb50f0d2c4fae1c91c6efd8d9416ecb00c1615de3edbc487d0dd761fafa12cbcbe3e312646f9f1d479be7d1fcb554f49e96dfb75a1bd44c43715d2ccb3d789d30c0854128a234555c6a0884ce33b412fc7cee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41964560d9055b8fc14be79f3d4228364e39b0a8acdf4507f8bf663acfda5f85f1abd6b486c75fd684bfa87c6c3b0375f0ce5e2dfdadbb756490883f583bc318a6cdeaf92ed5a11143f60719bb16a594ef465a0b5154993a42f4f7c0fcc0d43a7e3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b08508e899dc3829ab158f6aaee456deb83c48a52e71ae8fd560a4ce93cac7d2117c1c94bbebbd0f8313cd55556247fc0191ab3629b78fa7b649835b7804f4d2da3cbb882eca43bcec4ce6b5b1edf3ee6740a11caf5466d4d07d9ee3c6606d6ba19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1ca5a4e4650268b5897e5cc42835a653bd066ebbb684680025fe4e79b17a879843dd0e63253765ed8b25fbc953219dca1ac0ad62b115425f9bb3c803d6f7edc64183c76e07251c76b850a36ef10ebf926946e9fd910c719cdf7ef3444f8061670af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc430803a4a2ef365c80cd8ad6327931b7d8be1d10587d659f456ea534b6bd45e62f7c3f70b36c41d5a15f3640ce40704fc4818a8ef78e07b0fc9abf390670636a4d5d1f8a214bb687a0d8ac43e6e6f4760f5201e59f74ae62e1ab848c64d75585298;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f0017593b68e0c4dfa88ee54f92999bd5ba203056cb8f16b0daec598552f8a48eb5c8f70615035d7b84bdad784af4d1aa5f3df38c29e87b665ae5c14cb100ddced6bd21f059220a72002ab89008d52a0b85e778ccc3e1110e8a849441a595251b1e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ce876da8a6386302ff80f5411222994687f0a1831d1b21422103ffeca582f52e4d3d2e585763153f7ccba0331e312dd6b8ab75105872bda827ab99e41cde1569bac2121e2a5afbe18d0507df12228383b4f0a2644e103ef6bfeb6f3af9d906b470;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fbc55350386e4ffd168700e416c0217e38674a9780db6d3370e0a619a32a088087efd42d3b506e0821e91eb979e7c2513bd7946241fbfbd6b818cdab9d6bbe86cf685186611448c2d5ec96dc43c04c9eb7b55046bd804619ca04b9d7b995b9c51d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1167bc3d7fb87117e8dffb907146d574bd8df080274d6a819448f29cc37033c30d8169edb2023b5d1fdb88975da5dd7fc5e793cf938c3e07549d9392708ed3d78e66812cdbca97bd93a296862472bd947effe495b3cd5f6a0c78edb4cdcd6c932a77;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c771039c64c558e8cec408b8f9440a16e2ee939923703e1e153f07e349425d1b0b381810ebbb6bdcfd41c5a8864e15aae7f0b624ed8e5bd23b83f8e877635a5848ead6db40f249f77dc535ba51c2f093d3a4f290e3df2dbd53a93e329f709284284;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h606b0ae0ad89e9f6945f6a5e2399c1d2aa68d91c0c85d17f1d5c123bfab785706d279dcb7eb06a5b1d522ddd87d6bc11bb40e78b1dc0056577ff2f1d1659ecf5dff41878d5876cb4781575b46abe54d3ba032e65cf0ab6bebf9de5fafaeb3de0774b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h574a0a5c350faa2eaa45c8570588cd29802cb3754c6d223a7d74167dc4b48854978bf7b9e8f5935b615f5f987996718186d4bfeaba135e0393420d698f97ea94dee35eedb692fa44cabf4cb87e898331a1169ab90254cb3f2bbf49afd4622d7a9548;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cfb686e54c952839ee207fac3d3f3d05f40ae56136a4b2f45fdc3de2c458d78511f95933fac983ee373814dc49b9dec15f5f61d83911eff2b6f4072542b3cdde48c8351d63c68f116be9799bd51a75cb81b276d12878546cf99396b6751cdd43840;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39aec3271c3649d37dbdbdd20079a6f0a7d8ea4ff7d309dda0a4f32666371bfb3e2af60de25d68ab71f35e28a75591637a7ffe91aca6aaebe36bf8ffb267d6615f796debfd2e2a739e6ef5d0614c9ed35f1eddc03fd9d7c5599519bcd1dd051814af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53b29c38f10c7b964bac54c1c2e503e4c916e32de5bd75bb6c7731b35d22c6206b908d7284d6c4a8382c3c3f45b86c78fff5326ab6b1638069a77cb0a02a93f82b0cb4fbf231dca6a202dfd512c0ba2dfd2cb49905467e8a23e168a258ce7f9e09e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60601911e7b7be0ee773d83067d9669de4aa47dd368d5a77486b4ba98f0ff0e49012d30236dd4decf012e5e162de70664527e4a192b4e6c61c49ed55c08a95299c28de2be3225b6726f52e364193c1521684aec630906d7a0f3af783b1bc40d279ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha52c1509fbcf7ff44799582c1953325c92deba1d90787cbf6e470fd86354e6ca68461687c2ad6ee0d5913f33bc523326f303c9e26fbb566218ccb340b032fe37c1d6680f40d3cc9c6daed97771bfafde602e54bf8c91dbe40a6c95ae4700ea67705e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h406c2523af575a958456219694d65e28eb0fa4b88af30392f9c4e528a19f7d7b4fdfcbd7cf6f299a5aba975084a94182f1e2cc9d8440b1687623e88f0d5fd17dce4525e9d9c5370c69649929c6d76a8d7b582eab28d62394f446247ca13a70bc08e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6577cad224c38bf0be91e93951c17c4161a431b65452fc4d55148fb45790a4a51c1d18250b7663711727e6df54734f735f9d5ebe856b88509c73aa878047b14db1fa4ea0c07e74a909d215cb1ef7af3e9aba33cff76a787fb7e9aba3ef1cdcf5633b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfac2f2fd91602ad8f6e6943972a7b39595ebd705ca8b62f5beb0057e7f34cad854d3f3c7c9b52981c5a8ceb697040cda49e1d8bf8779d0da45c51b2fdfcbe72468acfe39281474c634749a11869758753c0ee33eef7a38af981f9233891169d22a02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d4e434196aff3a714b1cc8e854994087e9487285c0d57e58d5bc4556b5eb95b983cc2dcf64e3a4cd8a7611bccf9c7c8a8384e52edcd8486a9d349717628960bd73f0174da306410db3cd294234695fc5c3d26cf42a6334ac1656904f64f7ddad77;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6216c633a1c764f2aa229cec511f8c15535ab29d0b3fdb9e981bfc571cd9d335b1b6c05cfbdb14ff0d6283e1c9ce98c4e25e2044d94ebb2be363bf5376142a8a29c2ac156d87bf915decc77ccf9ead57b80157320c147fea03a668f9aad395e1d63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8f0974d10c7af3c0dc0364b03b34de88ad5f692a882bb61e862cabd6f039b78cd8a4361b97ce43ec5195882d4e2b4981d5ec2165e654567a814b65aa6258d7b149665296fc8a28bb3915e0b1e7bfc23269da19cca002eb86573960cceaa7d5c0cd1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4344b3ce742a7301ffd4dc65dc81852d3b45c414a1683cdcf1b6cfab29bcbe95e3bc1ee134e2892ad9f4bf9b8ae8b05367d7dcc9e1ac1f0b29d8ba9d3e073363a946b9f038bda23248f226f52e038723e5227de87648794b4edbf82c55f43c415c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf682ca493cc2ad17ffbde0d6e47d041abc5d17aaf59bf2c2136eb5d07e2d801a1cc093a33e32369b8b45cc7b58c7405d1d270310d8cdc32f4c5635e5fb15d055d9a5cf321284bb61a127e1ca0eba736367d4d1d70e7fe7bf664f9231abb011eb3ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42b6cd01935bc6c4ce94865d2f1fda5aa3929253a4272767678bc2e8899362c124f38ed390e241c86bea9373b35d06845f8dede45e12099aff21e9bd5a7515ed985f871e8030c67b2f8af29dfd21f3532a41b509a75e3cf14e5bc81ec3eecf930293;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h498a2cdd741956abb3e868fee49886b568ba62572edaa5d9ff15341fc2d1dff0c26f3b8a3507f909f27fed7766f83ae727be1025f268d088bc169c71f1025f9510fcf1a7feda643eaeaaa19d910eda8caf6244fb05cd071bb253e6c9eaab92fc2b5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19a2e0f42205aa3f0b080512bb8ce741611cd6ba7a1793774a1d1d889024a28626225ef48ae8798a9bec774d15da5a9700aa9ddc04dd73f06f162962ca1f75b30b74026ef19c682404aa09a0f2d5ea601093192be80646206a50e11e936081e6d316;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ca373cdf1948e39fb127495e1b09a4a615d9a6fcb007320092eecab0cca3dfedfb18d0e4b36d8ea4dcadca648623648f2ce87cf4e35bee05cd6678632da1bcd9ffd234a0e00e3ab7280a03aa167898a31524ccff7253f3be17b55ebfd92ce6671a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20f55e1653ab4cee8edb1a08f5dd5698eb17e7a31677a59889e298abd9ac724ab8884773aff121627e08b5e08b8a8651f79d320792c637340f07cb6c9e06c5ec136265f0eafd49bda3e883798c7aa0e5077499f168018a1db626f6975df135c9db2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h893beafb84056856812bce5314cc5f71bb690d2a23e4eb052f4e480d07e2bfbac72be450f3f3230f8883057591eeeebbf7458ba501966a573148c0129e50a3a5180f38eaa1c84987e2859fa148e7051105f518e67ca9a2071de6072aecc42976d674;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd94e51158bf14652f66c558ba6a8d26c1d76e947b3f1c2a90e03f21fb552ddacee3485d20ebe197bd3a6d31bfbb8ef66377234f9d3e7f7aae5e735f138ad93a63f56897dca6ce656129383f4472bf3ed6b2c312ccbad2d3b272c7b9c10183e36a0fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h536e0d1b2a8e8a5a55f9838ac2909f22bb009f0847b3d4562325bb26d771923b5faba10c2ed1b7ea8da1570f16b12c193a6a073c3e30b147f4b8b08e3cf178da91d624313c29a6e5a6db49a36ccd8adb5e4a226d6c12312bc59b89ded1b65dcf3ebf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16125b9b6b6dee1c481246567f21217a7790058fd517b1c8b4f26f6909c371a995dc6744b426d72dc0e5630209ed462af5009a5d57b8005fa9b26cf890c7c5a5ca736388e842398e99e8fa38e09ccb546ccb6c08d26a029d2619cfae3de190cb2b98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefacc7d9530c1be03d5554620947368c07cc4f86a1c7603d01890df86663e716c49083cdc7027f6bba5a45efa1d9a0ef800441204938c53302673af0c2f301c6bbe157e242606603e73d9abfe09c218c2ab9ed6f2e99eebb2dccdc801dbbaf405454;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcad0661d2b617f83d70471a6ce2abce84a790295996e5c17449149db377abdd48f1cd7c01f04b2ce81e0a655a386dd56b8415c59b4f7b5e811dc4a0ecb09e8ccfaac9ca72100e053b0fca6e22945b64c8b41f8a8b5106be3dc1eb9638b19497f9668;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57d9b16f55730b2e534a5de899092060307f8c925ae64db54ae0662d55215372b1cad0ccc0a496f0d50c91c7d944e0337714328bf59ef3911d5c5bf9c5b02050eadd6faa1d352d85c4aa8362987aa453794d7170bf7cf453e423fad42cf830f691f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3e309dd4adb588ea089ea63428dd18683557b36717a5a4e542c4c59fd8f73faf87c2bb0b9997c9d03564c0cdf3ec5b7429574db156b06ed30db5c9b8f5a94ecfabc3adb24e262af6f5296fe31d1459a3d2d0605f067eb2d5f7cff8e56bde30641b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcac3b650a201780bbc3299892fb97080e9eeb132787bd88375d56603cf40675d0358e43dd0e202e863be4fcd9cbc4be8de09ed8007e6dd650b067dc2caca65d703d72515c1e96c8628127d4793f46f98fb721d2eda4bdf13fb6b25e35a2cc89314bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h998ab801fc4029ba4b3bcf82c38f4a8c7e56f7da15db1654f4739612aeac1057f8f8bfead947c1c9bf00000e83a29bc349335a53c94431fa0e3efac3af755863ed559df00b9659fff85506515942c67eef473477d8bf2454b53d71e39b2b9273a00f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha51ff3e08918a6e752b928e66cd2d903e4c1a9d71d5018b94eef8fc0e884e3e684a7293a4d678fae3bd5d9ebb6ef73139fcc8f522dc7f545e9c3db0b0dfd01f90eb30a2f8b8ec497cdd83d1b5b504723bf79bc4eb6908f81483361f6fd87a9a14c4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98dc1c490e168fb60c5c1fcddf4cd66bd60ecc699686022f712cefe7e1195e3e9823bd4d34da730e67d17d13b9cc192d12147b75b4b1d32296af557bf01032cd4645de42f35590c39c36a10c92f02d31fb50859ebc6ecd4bb004e74d687ec84e8b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h601200f0851a5eea3aece2bfc0c27a8f83e10c378a57279fc70db70b046eba4bf96f2adcfbe6ec41d1b01ac8fc82d3673d0d7a447fffe6db8e671f8753dbd7946e4662cac0744458e1f592f16d6ef514ff8002fdbb467f09c860a95198878244f037;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h485cee7771cd2e6494ed2283a879990acdfeac1c233eb16872414dc5ed7799edb59b5bf949949de8763b9801b9cfa299664645383cbdccc073fee86e027e838bc43235afd2e531d7954c47fdbf6488bb671994c49f32cda68368c4a9f2143f0d0bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57244280007442e97647a3c8c1122ce7bef4195b64a348c9b139554dcc139fe3eac237aa446ee8ad3f98fbfde34c405ac98bf51d78a14ea7a1cc081989a0b4737a5bf062cfc1270f540e54f85b2335a29812054e3651e7d0bf6ffcca9c7b1d8a657e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc50a11cd570a5a650b79990116ca600dc251ee73dbd032b8d5f17a093a4e45f82b413ac702ee93aa57842f3d835b4da927b75ebc1501d7d01ede5e658576834d9e94abae5435530d37fc24859c4ab91ce2c01aa989c71ee5a6e8f1e6dc642b5890fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he98bfe10f8741bb4f67294018ec6d733c2f223b5559e204e894eca0e91007c5b4ee0eed760499835f7e96038f26e73af7c0b6fd4bc7a49ccfb39b586944fadfd440884dd18c8748c0094f341b55e966ad786c87890a25950d4f57c45e6b46f7bd9d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha851ef8165e4001e350486df00903643aec13d467edd1706062f4207bf067f60fcb52616ab98e2dfe6b6d2346fd034d83bc3f1a0001f1e6e3f824eccad1295b1cb6daa98d9e2b1610e61c40c20d37f13d238949898af243cb813e78623902c04f069;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d170bfde5ebc4dbcb0fc0852bc057b8dc3e43a7d1b2b40a34909cb2a126f79232f68d5f0d965f1c47a452182a6e8dae90a5bc49ff2629982b32ea444198169248defd59b871a7c2ee3c663acfa52195c15baa4ff2169199cd7617d4c442c3a7373;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30bf8034a58bfa86f7099161f797b725eca2d1c7a082275f57c76acd547feab716b01d209ff831a20dddf3bead0b4d2b9051c4015e19fe723e5d003d24a07fb9efefd80dc556a9b8e2799817ccbc04d569305cb715dee70dd30b80a0a670255ce7e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dc15082121b19e3a12ea9d3c57c6d1aecdb193c31a989f6d3b09d803e7728c0e2c0d40cbf7e437ec2a839783149db8a3647e13e433841646b885173427456d96c677f74d36e234871299b135e0a64d9b8fad8e68fe0e3a7aa515d0534eb377adaca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e6577cc8b52410ff3b404a42927bafc207fe6ec4e9fb028ef04081f9193bc9b6ee508fbf1f9b5b4f0e70d99bd3e840b59332bca0b1f9aaf58bbdc3bd582932dfafc70c750a1a598ab8c2c1692ea2ca6d2d595a82175aec6f5748b3ffcc52db8c149;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e6e3121ed2ce6ec981c77f7befc8723dbf1fd0565b6d8559d8853f139cbf8726855fd2af6d3c61d21e1895d30efd6ad284818f35467373a916f37c423c8bd8f70bed724ce5ae88a0f05e1f476d43da58eadf72f92846b7b6148f5d82d643d8ebdb7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84f1e65a026fd232a14be8f4a465547263000ad18575674b13abddf9aea74e0ea289de418983ca2cd4b70374ad8952db77e785d84db791e5ea2c5c1bfc0d03117422780389728d2e28465182c41f9820ccdd752c6067927d3e6f39573ac814099472;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc27f3b50e0ae413bce3c569425ca5aff79d883288ef9ef61afe12d5743ae22b1a31d12a613e021dbaf5dc3a7386cb94af3728c6d7beef13af7c832bec4d301b5099cd2924c73395b18145196199433401c11fa6d28aed52403ff07f72db29ddf759;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3b95dddb7e56998922b1738f2c24cab265044a7943bcc62d59204234a778226fbd1d8d32d7e268b6c2ca53522935dd1d83939dcaee868c9e32113be9b8f6e160d408d275af165c88d55dd5a0f231b713350334a43af65db24e058cd6e6d5fc88663;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87e07e8d97bd3ba61150fb046b15c9c10cfeb00b416a5682bd63a58128750845bef2274e8f31e01f0b99f048a362a220824e4ad4e07acb046d725e27ad994a765ebeed4c52e3227147467604bc5cb585c5d3476760582d30cf3a9005ec1d4aab20f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a6a60a196a1ec1c00f7425262c8b8fe6b822e19854e9f80bbcc9dae8851de3a8e21c5374102715b6a8c2fd9d7d72e3f5c152052ecb5cedf08554a016a7c70e0bf909036fbe1776705e364998d41706869d5505189270713c6ecc715c9ceb35863e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb487acfc6934b3709afca6f7c9cf9614c5262e06939e571d0df246d90b7592179f2145133e85bcf429acb3bdb2d15a95858657fcb5ba355262b2519d373bbfd69958c03c66b37ef6c59dff026cec0bce86e4d4cb2bc77abb4ae423db275bf6ec977d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24b536a1b3b22abe3f65ef66c47808308e97b38007705053de18a111658e52b5456021f7c8ffe15b0157cc66d819db60fb8f8d087c2c2b06f8e1f4f69ca02ab4ff4c05061f8499d1c0a66e2e72d77b65dafaa4cfbc9bd6e818cb41ad05186cdf3171;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb8d963962869a54c446426fc423c17a6e26f9d268bd003abe617b18b7333d8b66e956e1d18901aeb2a606c67d45c6ce7fc816417ba05d5ca63fb7c7e2d37b6d6ff0949159b886869782bb87fd7e523548a607daa206f7fbf370d15c67b2130969c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f62a9e8579027833475869e755a3a49b3676b4dc19951ff96e576922fe42a768fd2e1a7ae9d1214afb463551b37ba48037dc84d7ed97024d992466cce28ba610a9f7dee991cb8e48d5ef29fdcfbeabfe618ef3fbf5811bc1a4283eb2cd87d8ebf40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5c0e19e3df2e42d5c6203c860893b82a95f7bacc23e304142370640b05e19962857c939192a9645a52e34273869617fc02247a1314ad3738f55b0d8a43a80eeb60fb5deb4f38da8d2ae5109d6ef50b55a0e2165e4d52e2b0578f5cba59d9453ae77;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd45b088945b04f8c9752a902ab3c561ac80a793cc9a51f32d5b1d4a6b9459cfbb5c24f5de1e99ee9f87f4171c491319b22be6872abb5d779f18f7c97aafc78659b2c2f3f8ed6d2385a0fda24e419f79cc83fc5a55f0289a9e1ac09493d82f5e598ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b48bc802c54c39b20e4abc64f9cc213421485cd5e6f2e38bde984ebc409d2e96db14f6cb98e1b34e33271aa75e2f662d96e0282a378300391eeef2f2d991c73aa7b4562a10c8eef51b94e0ec734acdb169d27ee0b6fa8690f63b21c023aa48e1bf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8314a465c815d018ec057442fe4484559628fc67dc89bb8a30ae65116f43f711966b50eac94e020c9b5634d50c777e006a6f45886ad01b08631cbfb35aabd4c80217d26630a59c34745af5b60b3a7b1ff7d1c076b611e1ea09428f22f8b34e2315a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h606385f00e07cf3c08a7360ead405ef3a507366ec90022e62c0ecf51f415949f3ce2121c3b5cfc02c2354fc70d997520e1bacf1e185e0693008b4897bd756f882828e7f071f44b5643f7626ee2c8764892d7ee5e442763f735fce5ed2754c62d4af5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9af245210966aa14d03efc471ecf1174d5a50ec98676f36e871a20df29f99ee97064c8ca589b01b9b0b069742ee99876b77d9b105675470d3cd67db6d971a868e0d525299f4b72ed28a484d3cf3af4664309488193e5acfb2afba43385a34fe964e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5eedf6ed33d3591e860753e0dce5b0e326889ad34797713252a42428dc1f70c58391a5ddd508945d96ce5a0e51e91df3867a954f9599cca01cc9f2d761c038279d8b0a11b540468f84cd7d187abe782887acb5e9d1158644416ce6af93e0e0103bcc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc81b0579785c13ec6273d0650dfa0f4138b8225eb0ca6e830fea264d4a1b8fb06d38aad49464912fcc7190251ce614d9ae31d9ca618bd589be6d2da6dc684a5dc7f4760493d92ffe88eda264cd0d322c93f2a716fc791c06db312a7f592864411ad5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae261d3dc391b18ba6318c42afb85abfdaeae5ded8138e9d2325a2d937f99000341faf056e7a58e1de3ec6c04c64348048872b5ab9a94ddf940c2d3f0f9168721143021472d9c8e98eaf6161e7b874afbc9765f3cbc3952940010ab7c78346dcb44b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16169be3ce89b18aadcd9a5b3394f9c4f31e8a462620df3e4e2c553a96b463fe54f4dd393a6d2d81f17d9a773ba4f2917df84a6a49f3602fca457f2062ba8cfa840440735137876c31922012f0b71eb1f950d767576e8a64c3f7a9c06451ee170a68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb917d974f8e65859e1a82967b2900de8cacecc15b0d56d110885049782c49217aa006194c89e6a574af707c56de3d90a7328da85cba990888ad40951b5d1b9636c752edae82d356abecc68bcf7b5399ce759c01e0631a8243f94bee9516b07fac00a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec110cd5adda8983a8b980370fca5ed71ec95936abe988abc5302394dd5fd1bb0fd13d116b54fba353cfc9cb6d6cff8977b776dff548070d895cec8ffd32dca2d61273ad72a15da8cec665cf11c3c5e44368d5362f5fa6d099a2bbcd3e7993e68ad3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87fbf1450bf64bdcec278f723be0dc48dc81f575f6227445213f1d1adecc7c6f03362b41e88cc25ff8a04cdd4401899ccdd0f826f69378633911e3053ce06675c627c9b906963cc0faba2f435cbeaade2d0d0278c218b1d4c4313898c2d5acbac9ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d61768d3dd7bdc8eaee9ac6f6d872ba148b77fb12ddff1bfcaebdbef90fdc0214bc7a3cdfffd0c8a0e8faf69a4c448649511edb6dacc3f25197a8fb0184edc771ea299681399bd2fb44b77f7f2ad0790650c8012e0dbf2abdc00bfb36c46b68f936;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd439a1964e62e334d297c4240ced531297f84c58d0564c359d5c10e86705885eb8a7a6ea2341117949df5e7274f0152eb867b7380d7f00b500f98a6445c76f659451d4c68e4a41b7457f73f40ecf56c8b57773a7fe983d722d033e1defc3ec15f0fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4048a7a5cc26d1e93ed3b4a2c422d84b45bf6d47c08b6e36a161eb0bbed8d98513513658144dd6e0d979bc1d8b995b0f5167d58a2725c2da27bb9d2a8db32454fc488bc2c2c94b02b359cb04295ab7609fc9cfaac011ca98c535dd7b52a8f827112;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7496244e7721cec44358452b4195ef6915326ccb187a4eb06c102d42badfc980e95e1b75010475d0f80f1701fcb5cfea8d609b3e2df3357f9faf71608a0359b4b8a518171fff704f79964286a3b73de1d346b4f1b1b432d35f6aa6f826419f8bab25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27d9e302f00f3c154c6e9e5df3307e5b7896823e31cdb65777df53837e90e661162bbdc02c9271a10d3158487677777ac9b7214e0919d9aeffbe10fdf080b9e878de0f77010717f7145365beefeaf548ff31bff75ed86e45d7a6fe2a5042064d4a65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72c3b7893057fd5619a20b74f142f365b38a85604fa6d7e6fb1e587c33417decfabac2757675834ec8b501b2a887a56ec228257e06528888097e5bd39c37f7358528f1c7104d320387bbb6f9578bdd5277cf5c87ff1fec4a10807f7cebf13d603bf2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd68ba3123e2cbc0aac8b18c32d1bd8e412f382884b0c7c0d7b4f506fa873ce4132bd5634850a58044423bdd052eb415766e6e20947abbdd22580e69bbbf2ba20701a4bb144b565abfe1dcca11d8b0445ebe8ac1c590e274cd43caf06c7b438c0fe1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h607ed6b361251eca2fb227e05fccddca1cfad0228a61c2e0716fce43b761d1c5f417d874cd344efa93dcdd9cde2f1cb7d7cc4c84db35ec0eefba628826bed99ced64c67c154255187f2a2c0553c875e368fda6224f334271ae3489b94223cd315a3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbcc7abfbce40beb383db800a764fa509e9093b67f9d1b1ebc85d4bfda686612b734f80a96974f76f9ad59dd1f0d68873e2cc4411dfaff410275fc9b6ad3efbc4251d83c72d8db17752e16ee8840e469caaba52f480a71407e9afec6594d0fb8782;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h985d9c868b67332d6ace7bd2642ba736e5d880b28678ed0dc8635e4974d17d09d7bbe583c0b59065e33b1bd873015fc2bbdd1d494164acb507bce39051f30ce4786cf588842cae7861ab6fd18a955e2de7f7633a654b5b6bb17a25e4aa3edc3e3cdf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h469bdfe723d5f47f7353fe06ba2c7864e51bf11d79a935da0e0d3e55283251d43411f219b407147ec7d2c319d7ec89f30894792e684e98769341432f978f9086097dbb41fa0b8a9482e99b576723d7078a4555ac49953de128cce2b45508fbe74386;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b4d26e3c85865403bc9d071a4f340991ee73f4a2bac17ddd6ac46d048f0dfabb2d65bea726bd067efd7553a11196b45c536f10250e7e2c5b64c845048b65e9417c0323f19a2129ec2a3b066713aa2d1299a9a842b5d68681844e50a75ad91cf5052;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he047f06c62a51e9d384bb7274c17b5766a99486016a9b52de92c130019fc7c492b58f8e9179261ec004704d25ebf1333ceddd5a7e1815347ad5b7038b958cf8819f476293f8db61aaf77403099bd0e6c4a3231c57fe60fcc9c486475ab39f24fb4ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc386177f9239bf37cd20b313d2be42d59e37a6b7183e519ff80d236f03bf79997c02c01f97037d294035ae440be56ba4e533239417c6b24becf583f404c30dbd75f24927f0dd31a2cc65b1ccaf0b5d5e8e9e08b0ba899cb263e175de2809e283616;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f8e39e581736f6becf40d8b26143b9f22a316af3178ac9951758e811b4a2124132a8ffad6b4bb510be27864fc7f64102162412cc8f0fe7fa6f6131f61a5335ac291feaca086f7d0d070241e2d60e492541268eb7737a881f293e7b9cc7939713faa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4023f36a0ed6f7d1915317a4c77aa85a49898d592da1cf1d477d529e2c4873f8035089789511e20dc089b606506c337144474966fb2f7fd623c41493dbbaa34b0011e2ac485b36bd1f990814db613694411f0fc27b1124746c8094296ece0d81f4a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8446d026c2573a7fb495a98feae8d85826ba519083979263f2bd2e020bb133ac23d2edfd50ed66daab95b94dd6ad29c820a4570ae4aefddecfc7971783cb3e731cc4a9da5ef85759ec421e2ad37f6037e007ed3c168a945a0ab8818b26b403f09956;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc991a6264a5fd40c6475788f9ab3cd08ec2520386790f0819fd57335207d809e464c93fa5cd8751b19b8c59a24b0099ea53f28756acdea8968b366cf89f2e84918f51ad27941a804297dd7cb8de38762c2d11a44307ce70b14121aca38910384b1ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b8b64ef4a308c5e1620cd5513681c7c2b77a44d5bcfde9c7d6e9bd41d5afa09483cebb98b0bb96113920405acbd2acc351a9c20f3d284abddbc82c3a42ea0b1a8550bcfe6052456981f3f0cc38080a55e8101e28556ce51e727c98bf8455ebd5724;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd363a31bce5cf3e0d1e33a9a6a610859a22163d260c9cb536432f368dd891ae7a7185c7471db06cbf82b5d6ecd8f671c40b952795629a21bb476bc83b37be40893fcb7368b122f32a60a5f5981d23a491cb8ecd7d46c141785e1da6c313cccb7940;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h345ab34cd06962a4adc75a561b1d0ec8947e7a3e1dae3e6b4cb021920235b68a8e46bfd9d0a3ad4a8e810271506a676ae569708c8eca4606ece618f7b9f7ffc36e503a878fa98f31eff7c11c5965f90c416f334c51a27733da2e9a825e2b03612af9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf2b7d1446351d86e020217608d8d69cbf68313ed3e80bbb4dd4a0537702db839ff0fbe44306ed3733ee91bb14e65459cd5cf5afeeaeb051a7e4017fb88e1e7a77ce17cf28decc92c98c003258c4439252e7fc6510363a46e6274379a28ad4eba836;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h448a1d399896271160f9369e1c080626a28208592cf1469f4e1cd9be6ee16df049dfe03347f05865b8502f39c0f1b86502251a6d96df728452b93ed331a70739d7deaedb16d5b798a23009561010b53aa3f02071cbe6741291b8985094b8de0d6fad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h856965ccee2ad74de44acb7aa39b6ff8c5ba033bdb0c581bffdf6da028c1e4606cffa7ce8001928f323b54b36a1bd3a534d305e6730539a4fa906fbe645f457f69668cc3b688992d029f1324c8461df8f167b4a40f1c38db004aa5878a6e0aa0576;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f522caea9469bee71a5bd7e627f11a64154129ec4742a84abb175a3825040bcc01144fe6af2f78e6b55150699bb5a1b9b244f0ff68a70e87d834f983d3531eede5e90e984be07edaa6f3b825c0881f42d00d186876054f2fce41314fb34fb54f8aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d63c34ba720c9b5b5a4a5fb3e9a49eb26cb98345e3658f488ddab8d4dfb11e4cdfa03879d902980a61de7649277b1386867eb2ee69e327408c00a2ebfd7864e6825ae4694bfe6c75717248b796a55fd5248aa041c17fad8ec09ddf3c726a7d8c6ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a431c462e732e3ad02e344881bfa14d9d1df24955dee098bd2bf6634edd24fc7b85771fb163a18efb322d8b20ac33b7dd02988425ccde95919f69299316f42dd9ce3244a6d6b38ad95d26a8ef440afd56eba006b8266bb086b1d0be8942ed8b298d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe1b3ad77e3af55b28b59d27513da21c4688351558f60979f2a7d545af2910a1bd8857df7c268f4a9464407025d187e070cfae65a0db0fa4f14a831fa81e4a0a9df39ae9e6e23ad6975e613bb17cfaa659606744bfecd3d50539eabb2aba313b120d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9673a7bad44f478a5d73f4bf7d67064283ae0fa9bbe1c6ed424e32b7646855f57966c63303a28ead744baa6abede5f11280d4da539cc2c3528bf72e7006c10f3dfb20e3cc34d29188c1de97de262de2ef7b49bd0e3628f73523e7bd53dda97f6116c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd55f7b5aca76b25a6a35dc3d41ec0294fe9a3a5578c09bac9745ef160317df68d6a974e301d4a87d06646f4b7fb860aad56ee123bd2ce171b1b8359d435c0e10477488587956920bac2df3da8429c63374e44f33aac62150a86ce81268ae7393a69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7c6cb3ea199015b4398c450d67b244d99c4acc29988e1c7b2d210af02a1b04cbfdbeb99655f8883e8509bf2cc6c80859e783e9d5a1e1d22477a5fce75ff5021fac25c7c1b899edd078b5d31ea18f95bc2008318c50cd0fe1115f32a0729203772d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa171e11fa78dec06ee19a3f8a691c99b7aea836431b216db2d987ea3a3a6d1453542a006a02bc368e5c53f5c1fb505748ce4979008c6dda71698249355bc1cf62392d0029c3c5024a646c9c8af3d1aeec012b71d4e3fef263f7da1e6eec37886ab8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f5f7ad599bacd151146cb517fe72daf6424636914c628395c65a26309a13bea482426c474a9c4e16f6b005ee15de956e33fcddc03eec113b4378b73ce7abf9902bbddb05be55e1dcd4ea257f879d081e8dc32accd57f07b2d250c2f98bea0743a19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf2810eb9cea64bd87211daeddff88463fa2f17c9f99b7643e20d795d3710313fc57b302608d7afad7ab60977b4cd0f94578e8a3a3c6a6b7e1475fcb3ae4a289e4995d0c40e66b5df3e08810230b88d66562043a08402cafdc04462623a41561ebad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea43a71907a0202c7d655edaae4e492abd00fcd5060cab194f68a30de0c7ab0820951b4d4931aa1c3a1ddf8cb0777a84419813b3970ef14d4147b50628df132e59720b2fcca4bec3c0cc77bc67853e536c92346aa24ba6be066bc313eae194a2e63e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd034d344a4989785e258dc2a74376a6672223497dac27f627d526247f2eb9d20438deb2d623233f43f0104792320f88dc01ad8969cc189ddbaa0946548cab3a0020775f715e72a6df3ccfb0f0db326e230d38100bf3cbcf114e2c963acbd28a8effb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9c21df667faa9b0acb624af801eb4b6b611d15ca2cca73f0942fffcf8843e2b80d376c3fcfe30e4554b2f56eccfe91c5a35caebc0dea15141020dfbc45758338cf0c1c6a9b7723b60f6ff3dcb1b2ee0e5853458448bf869833007f57e2bde150263;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41a3f3c051064a59eeafc14bc7f52afed15a94ae69cbe8f589a003760aefa818e2459342aa20b1d2e921265f8256f6fe45c8fcaafe922bb67e1196905547442a811ae86388814e9cc2f4587786858fa4b23eff9616e6a520b9f43df3460862963cea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha026a77720519ee0f769e913a6d73f73b6e47acff6ad06290be50f804fff39c03448ab9d53e29a9556708438320a8239898174ef27320a9640f50ceef85b68475d6de98963ac4c0b5d4ead6a8047714ae30326b07713b348b3c036b287cef1cf7865;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h624f2474e81511b89d995d0509b82ed1b32badb8a36a01d26670b7911500c494ecb8867f142324d21dedbb67db91620a03fa4a9e4d4c3e5e6dfd72bc1ca7928264424025c7e6d38833e7c25fc89bfdd98ddae8d0cc24d21374c6e3a6a1bb12ec5a06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcd031e83aae581837fc8cc792906757688981bbcf48dc85beaa13a9ac9d2ff046913a87557fa2b111eceda2eee0376b6feaafb83cb26b74c39da48aa9bf36ba2f82288000697c4f5cedace6dd9abb6d8064a28ea7ab803c605a05b20a1a6a9a5b3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79a0c45f00dac1e61638e3a8be3bb2fc5edddcc1801bf2a4ca8cfd473d033cc5726b0222773ee952732436f49d1bd7f5bda15655263da9ec21c7bb2ffaa292eacd860b4fbb1c374a4de50a2d4cc0cb4085594482c1ba6020a9f8df767bf956259ce8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc35a763c68a4a0e212bf6c9ca229e48c627f8b887cf7ec4b35c1b167085d249490d5b8b88e69356e12ed096a0f5b521bdb6b708bbca1f6fcaa3312d2b2bb11ff1b0d4485670cd844013ff3e5d958dca59808b564965fb986391d202966916a17bff3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98a282be1f1b99db48838bfdb3a560ee64b375ae3096c62538d0a65b8dbbed8cc9a9605bb0f6ec32ab529c1b7aabdbe21e9ba61c8e77fca3becd437bd0eb51e58afdd1669a9812a151598be132e6cf6797a15c8c911281f95e5d1923fc904d9d932a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc100228e17ec4efc0b0af7d5be4cc4e2a80f0071d604039184e0e44bc669029a09baae61672ad37ee8957b95480e6048b7204626d9232d538a3504d5876f4f7c2be44098de7066b552ccf783ff22017329b12b0d5011da40b9d1389ceb7ff0d2ebd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13d2de046c1bc9c8e634631ff4d98352b47345b4c94fc76845881347e36d424e5337282ea698102f38a0255c8fed3bfb2bc08940418f81e4d25524d0dc71916d16405566065bcba0c876d861463e36d1e7bfb5439c426bdce876fbc0075310e05dd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h618ad3d160c4cb9b538f897b2e1ec99b21e80214f738b2ecea33750901eaa6366cbc09e94017d4cca80005607ab41490e5b128195adec64df27a48833bb25efa9ffd9952f973233df88c5b07a5febcfa6fd848476c4a50a3533d9a1898c4d8975e8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8caaa7b5bc968fb86a59ec36acf05786c14fc686f68c6579c2da78bcce0886d8d4c2d812c2b0aeeac12b2d3b4d2f95db5e353320065714de483f71e3711d7d85c0abf3116e203c6a678986f7f409d497a5e6e1fe801e97eca0d96540b91cd57baad4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha04ee3b1a29a266d99312bc8743629001d6416597abe7cb1bf03702f5981cd77f722afd5f730f0e2eb5232e80e4d80a2192135858e9e498634801a7fd49ac20fc37ad998879b08f4880ab480311662ebbbec1d52024b5048ec101e7425b39ea89cd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfd824ba97f27ea29c2c77ac5bfb54f5667a77a49d0fedaa4c7c2edbb95576c768dd7021932b309d7df8f3e0f11677a0f82e1d7d47bad442d3b97628d71d664131391751554392688299b66994cd096139f95367c1366e775f57cb6414f5aaf83ee7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39e66133fc622cf498e56895fed38249b5b64eab3942e44a89d700a52a2315aca62fd5a2935598965ce8acf5c6880bcd907d40f673b44525848b9b2a38a74b2d1a2677aee004fb92447af017db85bc16635c8d354d2f6e4d3b2ab92a02d3b54a8e84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3473b88fddd3674030b6c2e349031bf3045aeecf06b65fe9d0ea2b9020af4530ee4891c1497e9fab979951580beecf16f23ff258c3e1abc8408352383af9c1a563169524d1eb93ca17d4439e568dcfabbee5a4477eff5e251e23f22288dee6145af6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c8260678b362adeefe64a44e0ad72f0c1906fd6e072e18d860207c61025f899bf15f97c08e7bbb1578652556d49efb680eb2409f14aa6f5f8accdd49953d2b80b1f517160519d1727ef3f569d1a0d1bb134614666bbe37837f203ca86f3d290ec4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98126ebee75c1a4fd8711b5de2ed0182a4ba0aad9624dd8d1a9ffa74dae4303285558632bd1658c95657a65cd0d8644cf66118ff783eddef0b25ad989511b99c7043ef9e13564af8b8d8e21119a0fbfab21499e6bd2bfd32d7104fad6ec3365fa831;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43e863fdc4abbda375222fd818ab3a3805c77e83640e789428a632da8580624e1829c648814cbe47eaa87dbd45d4692dabf14f5dbe52586258ab853751b4490d0895eaa0fcb06a0ee4246a8a9905db1d229ff1b97f8352cac70f13ef2d6c07e4c0be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d817cd7b25993b1d1652a1ec39ce45f367ef3114f0217981400f5c0052b9a2c49c0f13918958172e855f11d5e3205baf3c0141a43d043aab44cbcd2c8857b720455c4e7acb16d0664bc4b576193877b571b753d208b939dcfd0000703dcdbae13fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46afc21bfb7d4fad8a1c0e6a5c22049af9c9e4e8a3ea72167075cdfca60121d5b28972e871f800081e5872fde9640869d085419a043cafcca159f921af2d174bd2f0d1363a620d3aa9afd3c672b9cb0dc5d0466a146c845eb09056ac5d6ce15c6f81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7418dc402f7cce305f7f0c30e087a81b57e9713af521406c55357adad7c971daaac520b10bd4a0ca808d6f2202a3dd66d61747166937a5062c266506f38876560999e2cc7d07e8106e97b5eb7bd0128037ae72f81db54cbdae53c999905d45d7c0b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bdb0549362a475baee99fcec02d735f2c96a54b5b0b9b9992b12925a04d53bf17ce4aea4da13c447bf29502c337fd68f414a59406ad79c9355c0e21621c6f51dd4f79a6cf0471e2313aca337ac4875bd422324410af74c3a165b1332106442491a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63af0f1b1788280a8651dd8b24504e4ff0e4bfb79e7c261d5e510e401b01ce3ecb63784454b3625f84561f706b4f1ffa7aacb77c7387e417828e2b55583e455d4712f248b48d395eb6bb1e044ebb5cf8d1578bd9d2b1d60e7f739c176f661f89e290;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb05e2cad40f944f64e095ca3f5d1eddc9c5ab6e77fedc5de0246d3188b151797f7e997880a22ce036bb0f3ea824448d1381b476e54a5b45cf58fd550206adaa9f7f0de1bc2c9de1fe2be653ca6fe9a596ada994c99138e630119a23fb22e3458fab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86988448dc4b0aeb7b1a539616aaf6b6eaf237ebd0c1d12e4403ab72b720b7d8840260da40bd186e5da60d3fb2149efe1f89b02b01d32b0be4b82ee2cd79dcf6e30218a48bd155b8161aa1684b6c2ac5517707f0674bbeaa0d1fea5f5e61799c7363;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcec9eb20d4960aa15c3e3e0a71d60f52b73205c30a293752348555dec913ad2b59d6d993d744aa7514f82ceb55b59b7c15ce4782ef3bf52bed070c66bdd67a8e2b32544847163456d79d0db400f2639e600a8031ae4da6da8dfd0a771ecf434095d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc812914b118d8535b0a8b49a77900e02782820285cf2d48394dcc4042135ab4a6da09306df83e0bf4100d2582ce1629379a7bbeb052fa28fe082c6974d870fda031727f68c5655fc1ee11642ce7dd8d0b92252f3388148ca39e8e3ac7f47353d2cdb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h366faf22b7c7964dcb016ae271d271ccbed0ca1c1d3b32a60e0a799e5d6125a6c8c3d0b4d9d4d2ce99544ef19aa951f69f09d3f86a91ec0b01bfbc2b8d6beb85b9ac7ff1c2a94a3a9802b7f2deaca6d5d265744baac3a8e87a1005d49fac8ee3cfcf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h624f4c972ea4a9c54ff455fac8e9887f68b3c5d38b9587b8a68cfad22f5db92dbabd56cf4376b69aad9e2fd7fb6a794a8d4cccc35c37dd9ea139eaf49391d1646dcabc834b796e44545bea4e36596421a4f637ce475d3973c7886a55bf273d3bded;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc238314c69eef77223ba26d0e0f1ecce95f0fd81d8c6f6bce7d5515381e5401d0ad8ae5fb5dd6a60f12e32bdbc3ab00d8df38170a9ec8980c63621226bd0718e1d0288b909ef4754c0936039c18fcdb642e70a61fcf644b84391ba546233237daaf4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc565f9ca430dc7e733140da1b3e220ff8c67273abbffc7b58c6c55410e9ec956295410bb1c8d68fe6dddcaf94784d5e9c7aa6e6fd073a0fe7e71d82122c6a089f8d3e77e7a6d7455bf6ba9eff6c3a032c298c69103d5e0c38d85d2153662f0045a84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h172a05aed8907a846ad1eba1ae2b7dbb7af740fe907c1bf7449ff9b4219bdf2569a9030e8932e183fd4fbb3bf1d20af16fcb6fbf04429c3b9c080a694ea0f9b582d0ac783a04a916aec8a77efe805ba29379776a6296503dea2621e7365961c4b4a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d577c0eff91e4c7bd8d8357b9639183d9a94b9a351596c58d0ff14a07c771d1c24a0c792a98bf189ac3d9494efeca64ceed7e919be86e24614c9fe5512a97edf573f13d2e65ea833e09381b6874ccf27b01d0bd689cabc4e0ff79db759a5e74e44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he94726c28132c55269faca761005c48a52a4e4e5192293fbfbcf991aea5d95912b39cbe8b9c5692a19ab1b3f288a677bb52485ec3b9cedcb8e858ead3d179129ea8cf7224169417ff1cfa1379b3d27eb2feecfb8ca6051daed68911bc76412c4ce49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b6c684c4f4973f494eb1e494f00934e75688d8d8140fa56e925650752e6975c1edac77d43fdfa18f8c1abfbf85a7020fcdb640776b11d785e86ca26a61e6eef366c5718e3e629213ca9acece5326213fb904435a7e72611dc10699293b4447f93e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h264d741903b55b1af9ad7b07b37b703dca34ebbec091d59715beceb3253dd4a63e28e7e460614b10c8557c60364732d96f96d23cd363f7646e7f17dba7c99b0358e73668b1cc804aef338be0ac7e6aa3e684b1745a4c3773be4fa5da4b830dfc6234;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbb6512c745a8e9bd8084aba094a4604210a37bdd7001fefd5e021511d2de377f6d07935c959ea651298bf60e8ed219e6d411aa7781a119ed2f3b8d80400da48fa53943b96ad300d13f0e4a6f2e3b1966273212c8b3fc690c602633f3f719c6b431d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h674349de272e4178ef29a3de996d27edc0d80e1e6808be03e16cc6f55bfa4be4b53e2506057622494ca749f1b5f6e5ecf813d8d7e5f84c00dada234ce329c3e99bfbd63a9cea368ecb860e1a4a227e974cc9ee648bb5f9d9826fba7724fbcbc403d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a7463db4975eb7e894c1137124f7fc90f60f7f96d8c430ed98f9389ec89c624000a9a62c6cefeabc4443d3deca2072633178a7c102534ce68938a4ff1076289cd9f0643ce7226fdebfda186ce2536fe46bc4afd5fe627b3ddfb8dbaf7587a5190f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf91d647ff64fe6bb04f8311643a352fb4e96b602e4ce6a26d8223c8b00faee816c25c7a0155a164d20ebaa916bf045c5c1ca1d692cae6dc40eaaa08466a7e2a6a0ec9489980eccc40175a0ea9c82a95e58631ddde2e0b34ea5e5a4098e7618488725;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ce67f7fd3c161b0c8ebe70d02217b3db44c69718102cb0ce578a6cfeb0d52d1e8e9a8eee51e51f690e65732f3e944bf07bd459528e4299cffb650672057c93c0409449300b8b7d43143af4cdcfd10b91e6956d6f2bc352f30666703448f638d39d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c840dfe64bd06badc559da99e93e0727d19b956b24baaba61fc7df58bbc6f1efa38f3c3ad6c028d8ec3df0c04bbfe90654c751cbd64cb945fec1c7d1071adce4656c151416b89a93f1ba2b343106001a6db768d7844d244643266546f0c14ce8618;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8e4263384b5a0797beff6ce702b51a0be787cbef6ddd3de5c05e104457cdbb851dedc34696091760e7a004d5f6fc8d212a9955529ed6da118872be0084a5de9d4744e18d3a7e84098b4e5d6b22f04452a8f516532a3051f9073783608365576007b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeff6b338fa7c579c41266ac913e0747bb43efb1a1cc8dca9ee1a9212854b2e427d1a67c4b66478d648df49b1095e0a14417234d2096d5ed29e2c69781335e8ded9e1a89078444c927c2e88578af38e7e43968d3eabc36456d59c5fd71c0e15a912;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h411c70f8106717743312a0669180c5cd70fb05ff3649a2c36af6db670c50afa83325a2b040f44338c51d3a4c0b89b2cfe02e2d7ab39732bfd3e0bb842539a797371e1480c6f8696fe289034d173010a651e4b90cc592aec0680e079def7c4f24420;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d9691822a39c78c3688dfeb3dd2b97f2872deea8ef79d5ac5cc52752510a1c2edd9e1482204963ec7ee5434e4f6c8031c78aaca1e88913e8402717b25dcab98d8792f4d0ec13c5145f736de2509c69c78f2d9b257e04b50c1b5dac87891584699f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b9b386289d85d915ff218f17be5e7efd984a00da7515109c67f8eaa830c3a7420071c5a148773f91d904b5dfb4b650b759c011bb2f02d1e1ca013b9cb3c149c7867f38d37eec4bb2208f4ace87b02ec987fcb69372c2d67f72c3d6c4738faca8e24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef5b27e6209b1376e94f8c58fa1c2e4e6e0b995954f40443e5380be765ace6136a127567d1ac3e2f1058faace02f356704253c6c7d547ab4dab7fbb68190a6386d88e8481f5c19f94ca37e3d43e75f1a8ce847d7f205ad112cfbced3e8c77d6935b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h298cd814285209e15ffacfe09f4da03e607d109e8722b289ca36881613a40c4c283434f0a211cca434d0348bd2de2931ac68b33addb3e22775953437725f42b665248b103a0f38bb8c1293de59e46fd5582cbf9c4244f596839215a62f23e0101eec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4e21b179f2e4fdc8a9d8b1fcd5a443dfce09620ae58f727eaf4bbf7815d6e197d4ae7c1470346ca5a0ad6899c1d8f3f3fc3078b8c46e473e75a58c5cc9c768a1712e6c6edd0d2deeb3111e92e5d94482ceae4f4c4948f3b8e7665e8d8f8b7c53f7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h738135b18c82fb666304ab1c948a526d3a4fc34d8af3b5d4aa9b7dcfd1aee807dd17a12d2b42f14bc277826161073fb1c687ceb0e4482f4f87fc465a3c805f74cf316174e984112b1504b9e009e39f0faddc90d46c5d6332ae2cc14a93d09a4d1573;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb03ea8254e578fbb0004994636752e52b7060f605ee1c39b949a8b7cb284c87ed624c8e64ce3c0f754cae79c37e661540b7c724c2b5597f3caf53df4dc9de458ac72efd8ea14b1c91f0ba9cd341ab19b3b57926aa737cd1a6184cfcd97c36eea86ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cb72a2557cb64690675fdd57f8e4ab76840e9a30113727bd7a58ea1c1fd6dbb394bb22ef94ed52a4094b4a8da88ff36aaf3010c6329a24a2a3245bbc2f2da028a587f728730573769cf413173e2b47677a5ec48a44ed41a3b0295f35303e6405be2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd1822ca31ba5f174a12d6a32a01552381376ded97522cdd84e5e3315e2450e45ad5af33eacdfe83d7f7c8131198d268d8d49a46d44fd1d73776ffd192ee2d22559597a10fc31f4fcb39e6df258e073b427ff05d4520f79c86d13704ad9cdfaa69e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c7cb79842e3e98534448c28d8b599ed354eff6bbae1bcc60f0501a9021d0961fa6669c49a1402edd01f88f31fc5e88dca4a37feb8ea1fd93d0d5b4c24b531e8f9c03826fdf2e9288daf40f7c3567f1c00d44c146c80c74a8e7aab67e1f633e4f991;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9aa8dc2f68537e4bb5241d0130b7c0f68ff4c7a943cc67741e35d6cea6aa0e44e447bfaf5db644cbf6f27f60022e2c10cc852c87b8be08be1268e96a82cbdeff53b40805d03a1ab263721d0d0b250166b260eb9a6a226ec1ce162aa2c1a08237cac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd577edf4baced91f618cdcaf04033fa944aa21805e6f6ca748c8fe37616ce1e028711fe6e7f0dcedec5d6e6daeacde91f68236a779fd751ed989b691cdeadd540d52952e4360d91dabb054c53a4c3597b9e893bfb97470b97f8ae60e1f23bad327;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b865e39be69a7e5e81cbd3f5421ee6353cb7fc570fe8e0cef8b465b1736ba0df700fec8ce695640c6f2443e9e18a1a4ce46d3272622d6c5202aac9a04fc244c43efa0d220316ea93abad2726d39e42d3091e3851617864c517160807c4f8d0e5d39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h372a0c79801d6420de3b8fc2952b1169a5a5bdefc7a0bc7b1adf6b3bdccb45d3d0c7ade8ba19045617f821e825aee5f30ff9fd7249bd878a57b79ee9f5d3044ee4c52465491b7fd7bb0f56c18ef3c3d64f4e6a05ef06c01e6d44a54de62748493d29;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h325e3828d13b6d80c236ea984eb2fe921a29590e4ccc6cdfdbf3cbc059402bf9463752ec498365f737a3d7d8e6dfbcbfebb86a98ff907c5bc1191e12089dcc7c2924f32b7e84b047da785117528470cc9b95f5c149addc38f6040c51cca6d07d9505;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9312c2652eac8b9e201e6c2fa6c28b7a49a8f39b9acd94b2aea1aa9b34084b92b79b9e557edaa62bb4e8881ca6a17afd980778540762e75e39851227991d59b02ef6f582dbc6dffd32586fc47711391cd7037f1ca4773f6251994030fafb3e567238;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb075beed6d53f4c31aaabb6983b8444452a813b4ea69236c3b31b327a6f0e34473bf0e229f4aef824d8ecd497b2b9369e9c8b51a32dd5317c553fd02536ace511e1825f6c78cacb528746584ab05fce92a220bbb5842794ac34e2c1eee0a1e1dcaa8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29786ec9c6b578be5f028b3238e1c2728e3e0e54cfb767a0217ce0fb5ef15ef03dfb1b24b390087e7d7b31f74d9a48936e9c4178112e08e23b22b06ea8e0fdfed74c5b9be1f131f8a4f092734a50176bce8a3a02a03077c59187193eb3d42e011a41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b9b51cdb2c3987844b31ff908e3993c0e3f67fdcc13614c6255106c3f1bb193d10f6f9116c72f5453c15200b5d12ce1c38c0123047660e0aa50264f6915b5516b0eecb69689574dd27324879fcab563eb2061da84b128ae79522451727856b1542d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb92171b37e00a31992fec8df13690b6d40e7a266e415804c45d61d99429d69892b32f6c7d53b10b1cf1f44510ebaacf29fa9afd8b6dfc029bef8444000c633e27f6752622a2b13a75358525631c1a3e81e90d336bffb42eb0695e5713d867b670e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73efb68a78307c9ffb0315fb4c55abd62523109a5a44c324d42791032f178dea9a2a52832034fdb2aca37a18dfb91c0eac67c8d6795fcaeb7ee2f9a19afab5796c8a467eb20b0e73d07f82176a5814b23dcc5d75906d98dbd988a03c39a9abfcc008;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd348e5a40c3e9f1d000924488df4e92657d548e1e4f36d317a2f5b752a37e83bb50f626e8759db56a8bd0b8b943ed301593bc5be2f9baa4e14978c2ebb79a5faf96fca0306f38b3603314f2a18aa58991db1f250e958dd54dbce3a4243d387ff39aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8f18a9244a9a9ee4d207cb74e57552365084bd2b81e7e32b72f668f0aedfe3001357259f3a5933f387e2dfd2d841f2adcee2731862241a9348530fe16e8fe2d2d660b8cb309a4eddbb1ca6c60edc92e4393c23d2f18f27f737e3b722ea0165c0fae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5acfdc29d0fa84805d9a211e3f58cc69cfc089d9650995aecbb783dbf38d702d34e96e0f7d433c96c9ef6fe2d65dfe7416829a5b173f69a20f4711432761ac249462acd96d10672e2293f6d8ef20f0ecfd2c516de79d4270064c1471a038947f055f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb5be8e853e97196e2c3d4effa4bab53cc241139b60a6ca62e775f481eb978c126f81409c5e634f95df9a20b50bc09ae390ad35966c87d412810fb5d7c66936ed71c4062122a8d111b98fd6e0b82a93096219e2922af898aa51e2010e9db985e220;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bbf8c3b4e9da8f2dbe46c428b4f8f47b089e815d8ef1846f2daf30b46c2f5a4004b004a728f4987543aa730d4d5996b07ba3243158ade20ad628f41a9ceec489771803a103f0a00a41154ab5e5f592aa0179fe88d485a4519d202affc2f06846938;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35d511ef38225ae5556212e1c85d60416bd9b9c924c6e79f073b402ad89fbc91fc3630fa60760f6143bc34aecc3d43131d5883a64adc2d0c3bac353ca4553705d8704950c7e30402d20174f3c2a0536ff4878af65543e9d331f1b53aaaf293f662f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd299f676139bf12f937b6ec4cc80443a20333d5a9304c3f0f127ad8fddf40a9c2c97d03611a97ac40b0da867888d9507707aa9069543aeb24f2cf8026b9bf03114cefd4aa54dec1b74d7d5abd63630a91eb66b79b557a156ab2a13303a89a6c6ceeb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35b234e0ea6dd3528ac52abe4e61cb1ffc80fdb84bd95a466805ef4a2693ff801232eb188d012c1e65d20541f74ac8c86b2db77db188aac7b9c5d800bcfcd2ed02915c8a2e7e33f2d6c8653411788b36b026b4d632f0ebe06083350389e0023f4ac8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52afe63754a5c543461bfa88d2ad3196cd30b265b627a2c0ce667f91f683c43c9dc024c22a35d60d1953eef0d2f74eaaa1ce53843acf8dab98d0d03a56108ae3585038177bd4b073b323131608f79063442b4b1bc3a7c5592992a18dcf77e1c4c08f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3fdc4d29db7b72c4045bf9537e09c8237a186c4a9a793ffb662a9789c01b0e8833d96a93a8b1624b05df115baaa572fd165b1f8f15e9c252c5518e30844298ab80fe3cd3161ee7140ca7ec8f3d32a0e92553d8ac351d170d8942b12c37e9f85d8c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bc8e37f28e6a769462e29f826e485a22485b5455100ebb2a10c245d6235e4399fad868da45838355ae039f01cd7153ab46585492cf80f6316b535d6641bdf03124bfcd8e72cc0577c9ffcdae5f4dfddd9269bbd96fbff6548d391b3dd1df2e2d198;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9eccb8da17c9ae603f6e4863141a601ea2e035d3cbcc9f3fb1094a4e1ae7acc436ba12f07261d815c2ba52a3722b897e330433ef6244fc9e6519cb4e7e467cfda7f0cc4d4f91409325d027595aadb5ea5e04c90f1b86fb779bbea021ffbc89161af3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h740ec05218af1da3540bd958e2f97026b2da0bd202e3b8f7a271371a6e72528742c7e2fdcfaf91e6b369d03d6c2e5cf9b2ae3a98488fb74fc0f9a1f2e9eb3edc0f420cec60517a16302a05565136d765ce8eab185eac01cda093eb6583d3078a5d69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7de2b3b10d494b7df6b51fefb4436e7d22666bcdf38f4789941076bc12d4f652da99dec7198c17699a901fa8d5adcd61f77df20dec8b945ce2e6f549ba79064f501073a40c77ae09295fb9dfc48ee1debbc9a3f74daf7e9bcc448d8361ad112d328e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94edf27d676c42bbe310ab6c3707bebd2b18e571b9842707a9df104ff0cd1f1d52dd1dc10c187a94bb879874e39f733b3e4970e515976df4672d67850b4878e261e68417233403f6eab6d0519b66d50533788e8e9c79631db29dec4cc5ae738d776b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b8561c559967b431cd6e7c337d66c63c1bcef3c949f9213f1cd7c81ee28e7fd194f5897a0dac9a94254fe7adfcda4bbdb3369eee1ef554c183faf8b3ed2e3cfd1bc9294f017dc678735d45f7412a211f86f462ffd4635d42a2bef8a55c2991172b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc73432d986f79fccf71acdd83c5cbb5b36d666b8246fce93cba22a4e707c144d3ae6d8fb7997d62b108985c9e15bba0539984910c28f96d5a2fc3b664352e422ac060d3b4c30c9f612c29246b779d9df68da41c8b936a61bc08f1c0422ea80f65137;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49fb68b73699175c6df77fdaf618bf40c1207081d9e09e4cb2f636f273a863c1e15b0a98c6fde082a5e3070f6c0b34de3ca28e218cd8d9e5ee4a44880f0522651bf976fe1c05bf2e77e5271f83a6df9bdc558aa4d5cd345db53aea6c0d16281d931a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39d42c1b4ef3dface2776ba62343f491151a860ab6a591dda3aa468b93cac8a45a8db9fc4b3e08f313b52b92be148fbda824d54ffd3ecb0aa3c0f345b23cdf00a70716a288586072127f448f7570c21601b760b78f465237e28f3e63be752f65d6f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h698ef37f46be98b7bd664487eedc0e9683dfc62c3a67e69a50513c8d79581ae409f50369711b5d0798cf2a02250adeca27994c2724ab6fd487e51d431d3bc711da38193e6c79a9938ac562e455312d2b7d99d8259733641042eb0d672cd8a2f3cd9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ccc6b15af160fabb79eff194369b74fe735b903465f64a5bf524795f23f6837a335b153a828363e545bdb767cebdb3af1d21bb2f0e7749476281a12df86efe9eba00772aed463854152773afa7ccd8ed14b6a4b43024d05625f7062ab13460da6e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b92f0bc81540fec738d01402b12263dbf583e0072b7e55aa634ddb0226cb210e8e31cdb39940fd2dabc602566594d82f3f760c0a1f166f29fa6cdc5b647a890cd928fb3de09f4b5c761970531030737ce250364819cf500354d2a74720d0d9b7efe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f0a0e6f8db0cf5c93e012208b7ba9cc9735b6a6eef0e8ee933cf335beadc7a25dce4e95c4afa978a39f7041eb80ff0bda759a678c8fd60aef5759f56cbd2956e1f3892b639ec11ee6c485982e67ca3f13dc6a3fdf2c20a8cca35af4469f659fcad6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa92e5670c282912d1ff34660f1f65475721bcf8361907697ce57be65c928eb3dc0d5ba48b9cc8559b4e06a8a8b956e2c49da0d75a177f9b65578eac3f4b1091534d1cdf828303e7a68254ee72bd4447cf5d9c055b2b299b01ca6f3d4117a57de34c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ed7829cb3752506caf76b487830e329dc38c4747a79dafe67373198fe5e0a9c691c328ca5fc88c60fc78257e59f87a15ab3c365fda8cb6867895723a5c773c81453f60d978b77f9d4e5402aafa845d0dba6744ab2762d0a12bb77e3bc81e557c21e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf661984164d658c0c36a1487be3dba91c4835ad1d744761b4a5bc5ecb99e3606593d8aec03f04e40546b8b0ef54a0cddcc04b59bf014032259bad5125b293d02d6c43ab9bb0a69b63fb317fdfedb0e6922bb455058e8ee03231e9f8c2a3a7173c236;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2029666adc0fb94eb199ab3a9489054e2c3e81010fbd899f6f011293de03b8e6a152c54f1c8dc70831d815e5d631e2a918c9fdd7edabc1ecf52c7829842f4e8c18ad3916be8ae7a203088140e8ba20e56ce3c28afe60fce3aa8715fd296036af04b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e160ffe9aaa87953d2b0440e78d7025bbb137c73bcf822b93fdc4cf5b5c1629ef366c456b36fc9bf3511f21370a66d57ec9f36e930a569202a1c54cbcd84682bfdae24f812331868b8e2eca4d6078e7fd2de22131f0efb2a5e662106ea9bd74d10d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc5ca97228354ebcbb767854812c1335ce50befb6d93cb98830c5eba9cf351d1523c4dfaaf006a1a85ac85be70f56f46f7473cb7e5e5253d9839d9b57824ee5447de671fdb8e86d3bb83cf59beaaf6c7a62e58e7d7e55e6ba04c6dc2c1b9a34182e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h251a472ba9e4acc2c0f0d1ef91be98c4b2b9e10c92bce2957e4c1ea5f8327a17afc75a9ea71baa4dacee261c6d125ba4c969d1f33dfe2c82643ee0d4edec564cbe2e423fa579e364b70b0295428957271c540b9d5d99d60fd09bcedc911302a28ed7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1007b376ae8007532e63683f6cc0ec829b44f2d555e528b4f3d158ce48dba5389657db411d4ce401679e0a14e5f3c9c42f55136e5e82c5a6d89e96d5f7473bb945393b287e19e96cf9ed3ff7de08b5451ca7e52758dcf2fdc815b28e1741b9b06d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h535192b815292c52c347f79b9b7230896f52fd56b74ca3c3115afdbc65fa6bdc3e95334227493c461f082658dd0977eafcd97f290b7bbe2c664199cba3bbd77b3f2375d396fc02dc03d01c2561f52e972c3be9b290499927844cd441d0ef11c04fb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20548e3a267c1e44816b7d3defb63e56392002ac7447238a382c08a734867892e048c5c19b3d9593a97f54a6e1484ba07555d9ae07d5210d62287c8172ebf923fc2fa0897b84bd4b7fd949388891716f351ff15311a2a4b2d0ae219ae386447b612e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20f9edbd079fb49f51a5bba62f1ac9b5843e2b8fda5f0a25b5cb6052a89b20c5fedf360b3c05dc14cce68d7a3d1985ee07af7eebdc94c133d376f83872cd5ca3423c04e9d7da60d6dadfcd41c378fb38cd0a6814cf7f3985105271e20962b916f66f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bea4dd3e201ec41be8dcd8728ef66d18cd767d0f7f556a244a2e501cfae9466e55bb5361756feeb21a1d620a21d9e3d5830a2f4a12286f903582c3916e0aa6fc91effb753c7abb60ea26a9404a7639ebb2cc3108398a99006c2888db024b29d8532;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63d218cd2084c8e25788acab159163cdf802516d5afdd74e18d91d60c3e0ecf0c46387c68e168cd562f63115aef5c7cb9f8d34294f91a2def5c3883deafc7721a83d6836710c53a1973caf864d6f85b6f631757933eacb7aee10c49fbac137e4cc09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h437a0f603fd30ea5774a80fc5e4a24f9f4cb8509acb9983ca69789ca753464ba639a7e592e72bd861d0546ad163072e28e26abe1355b69b35cf62272469a79410a6c24c896b275d08b78f8cdfc0cfc36a46bbec6549cf210c5b4db4490b39568507a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88754541d3470daf036a287fbd53e1d3c3605e8ced2faca19cc3959bc28be91dad33d25ca3dd73c342cabc3ffbd5dd2abf645e6f8feebd094ec6ea51968a85ec83cfb99f46074ddf94767a12e625abd898cd237a2f7e19597ee4fcac12d4765c93be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8483f8a279edce0de843f4b204bf128c25380e8713f129c47c3e007bf090693440e4e8d3c7e4986afc2b771cd11e2103bd8d769ff6faabf12e0274e0976afe9df16d509f5f971b7f64be4096d76197c3b832fc0ba78086a1de871f0bae9944334e12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h745c9af4bc7d5521a28c181de16703ec3e3cb2e5ea0dfb791ced77332f973dc1922e149bb2395893c326c53da3bf1076c7aa04419641bf678b9dd46df2e45a3c97c9294a028bf73777822460b8b83346a21ec2a025f8a6c24891b3c19582f3e72f89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac04d215463480340052194065048471b4fa6b1f8b761569ba8c38e28a36277c9842341e85019e7c99d931cc40324e41e8d68b21f7c3ace48f6c65de4fa2a1d7fabe118bf202c2fc2384d73577ba572dead7c8a9723bdba29b2af8d4c93d47cbfea1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5c1da4fd542f7c97fd17e3aca3cfeba7caf8de5b1a1c17ea53d7e78c1fdae5bca241d22c021076153009c82f4d326f150bcf6bc2bcf6827aecbfd23f0d0ca445d84c78ed6d6643695aa62437e4469025f54b682d011c0ae3b383f3e681b78d8c9f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5210e7f786ed7745e560cf1299bf8a2d6ed09c6373772fcb19933a19ee1f201f9138f23c2df86f83018a9973821409cfd8832d15690d50a660b39adf8866c8edbbe0fb402b1ef612160ad8440f0c1039cc1756675610ad667cac6755c09e13dc4c8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda45230c64f240a07df52d9555f2385b611e0f5e627589e6614b1df47d009eb2501ffda6ba80fb75c39b9ae4a9a38f020f4a6e95e74713a5bb06728e4392ff7dbf71c7b506178ffb25c2731e549473bce2ae6378f5d32524e9a30e8348b5e7783a62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfafb0dc8cab94c6f435cfc6c67efbe0406abb1a497bdf22c915ffd89b83f15b9d0753d405744d9017c99b98b6f140dc6928dcba8755e02ae8475d984235fd0ba0e3273eb07b3711441f4ff0ecb13f3fa1db96dab13c8955e76d5efcb30a7d1fcabad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84dbb6b8a3f8ee2efef87fbc98a21d36014224eb60312aac5e47785bc0a5d77799a10b47ac447082b082fe7641a9b74aef0e0768622e1ad414d8e34b3ff0809ee0fe6027a393f9f4e9bc940861f422307cfb762d379573c4e019873dd4159b5c319;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf1699c2e1aa8722d99d1f4898cee8d4dae477d5cfeea8433ee19dcb3dc9dc7667606553b630d12d611dca8880e54c8aa496086fdd0f51e703d0840502089128058661995293c5a253c5503b9c912ae890d8970306a586888c8ab5a3898f8a48002;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11db54ccfb8b6d81e3370852e2ee9b441a057946ab83361bf626f5eb05afad60c1f2f49d233161b216dad498f92695a860facbb0bc905146b15e459c8ac46c22b83dd850cb856a08c024e5ba60f9ae35b12a3f5f0e579105810e24c4624ba2f62acd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5850445d7b8ccd99edcf2d5df914106fbcffe1b4c02e3d3a83e7d3b13f16c7bdd0019364ae3536004428ff772ae932309a995096482282e0f95ec9f010ea0c39c2ded760d4fd47aeddce1582c80655dd86dd6bd11a6f601023be08e154eec431709;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69dd6ddffe41d607bc5d23ebca01f885f9c81fc5dd73923dff35ede062e3ecb7484601ddb24e033d2ac0ba13f26651f30983f28bd27370cf7fa97070b37a5f49ccfe002d8b2b8125839cb64330e261d4790ec6d58696223184495b2d2884e6bfcbff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fd0a18c79dcf28b47a6863a7d7a98971f442838de87d9fc44472dd09f151b8d87bfbde156fc012a449fc59e11f2ccfeeb9633457b5f67037d7115b27dc777a39ddcfaa798fa37c430e38114eb902cde56213665910f22de2122b5dcc29e8568a90f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fea6343c3ce7240a830a80178f1ea7a8a5567fa41f1faa2136175f7d99f15460f06568c7a3a193a519f024a9f4558b412485bcc2ba25817201456668e8e29bf956e96a170f607526bcab1dec4d3f1209d11e3a18ad920dcfd29b1e09293fb9995ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4ae4e3df05aa0332cc82ef30a9a28df071d001b81f9dd51a54713f9d47805cb1b0fd20bbc161814db396e7905ff1f2a96452498946a43cb2f492796bf1948ff7502804e656c5151028b1c5ceac6fa3e88447d7c0090b6ef6a8a38b6c3af21b4333d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92017c643de9515e6717ca065310e124bad73dfa2afc35e43f56f9e2c36496561e62b6999bfd03d2009a9136c309b856040739c1b5f273f830e976c8e4ed328b56da92d104021c7a76e4681865a0f3fc7037399ca83cab56cd47fa21bf44f5dcfe20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15f32e3d406076e32db43c5578b835250f623584b8bb168e54dfad734711b4fad1fdc3b1a8362c4958830de779510b7cfac56b8faf3ffb7414c28f145ea6d6a776c5b039a0b2d4dd9c23199a8bd9975e70397e2771eca16af2a828bbaf33e0c23a0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b59810c1483ff2d103b4acdefac513d5a23e5c451038f5763fadafcb9ed0b3f3735de3701f933505bc48aacc64d3baa4887199885eac0015ddd073d3d5648295b91a9929152150e1bf2575d4abb3486dda8a91fe5206195d0e7d07873cae0549acf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfebf49be0694b803a8071b4c6af9915c907d6d791b8f5f9194effe4178e3d43b4135af24d7b95f9b4887c47b2545843e737b74767b3105c1ab8febc7f43ca44fe1abbf51806f2d65674718599c8a00f742f2f774181734b5c7663908c4b2679e0a41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4647914a8d9e646c804ca8a0d2e2930263ae3b7138ebba21bc016915faf6ea035d7cb8352e90164f5a47496711f0ede767c0167d61c49a42ffe7dfb4a75fa8a1d07d0923a22187c0cd83b1159e2d954719d74fc551064454a697e3526221c5c71a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d1615cd1c3232e14002f3beeb5a7febba1e7716e261878e551b0fb2ae2e5bcb63fb8d0703599774ce8cc203feb07343fa64c92008cc1206a8cdc70e3fcda7b4f763d4bbbad9f8d026f22044b4946db9e16972b59e2cc858de1296a0936b06823bdb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b6c22af3419cc72ee8660091156d6065ca6b26b378c153f544dc5856f43a0d8c195a09df792aa0bf9b1590a82e54531d7a3b069a1ccc62d5c5a7a3b24187c678b8e1f965ce4ba0f9a0d2979bd2fd8eeddd84b3237a1f22abad2b3a914289287998d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h809d289d0028fc36e4f96dc17de7963d01ed020d22ac5df48061c1dfc166c630586db78c3b9607af547c2e7a27061717882553f75b800bc5360928a7adfd5e5851f418277d26f949bc8833f02abbc4000b4cbc471c68d955257565bb545d53685634;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h233a07a155475a13ab08333ca10dd1b453d5106eea34112775b0ba02e991a17b36a313ca6a5d22fce93363fa9071263c43ee8e48cb43c06610d00e5169ed8233c3e8b32abb50799ca23b27939e48dfdf8ac55cf21da3a35a5741a568674d6bd37bdf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafef7a50d69d6d2d030e4afc783c8f0511240aff6d384669de15cc13d7fcb7cbf3cec2fd4ce9fc3279442cac985b0b0c1cfb3f0417fd62510313fd15a69fe9e6832a170a916d4960f40129df7764872a6f2b9def3fb233385315f8f887e594809735;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5888120caa1e00915f45b04dc90a9b358e8673d48b3fa443f1803b57b004ba30e74372e63eac95649017a7e68c9babe381e0f09e86a19df2070334f576dc9a05f2db63b72927dcbe0d5c5fdbd192e7ba43fa814f5fdf80e8d6d1e506a43637481202;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had55ec99f839568365ffe653eb8fb0ca1d00f115f5f6419e0dd3a043911bcdc3fedb80d309ec924384cd8346bad50d0bb37461f7bf18501777a58f001e376aefbd0e240da1a9d6f69a128ef1b910cecb4b9d1ff7df734aa69d01d95e121962519a9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90942b03ee698314c77f116aad9df615f1008829cd7a9268b60104d9c15cfab53bc25d9809630d1c7840532a704a70c475eac925ab72ff8a70b709f60dfbec8b61512bccae128a8a9becbf87b0dac58e04e014650a669cbc59c3264058f2c999f4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc505b9771f7ebf9e0ee9c530776c60171bace43e4b262f1188d55a6ba0bb1598770702c952cc8cd78cf632a742bda64f76f264b3697e1fef0aa412452caaa29cfefa46c87b1cefba291caaffdf0f2a2c45935f9bd1ea8ee8b334053df526ac19cb4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2900823ba07a62bca258b72e937ffa2caa54e7d3a0fa5865a34a22e7d18866bed95f8b4bd59fe44cfcaa0d18412d07751963bb94e01010cda8e4da7a7df304ccdec628138a1172789e3c8f44b70312a963cba5936a4502064c26b2505d827028f8ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e91e89648b8553e8c21ce565a00ff9abf841f2107e0883b0cbecd87059031fd7586afe436cb134142690376e38fd1edc5d02c603bb8a62ef3b200859f31b095552b67810bb0b15762cc5aa5c5c56c9f225d7016759f0f742a07c428f27a268c63ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba698c14bb1b79c2c00afaaf6272c7eb00498b6811582e98f85bd0e525a188f45b341435cf44b282eea6b0a5b52b3ea9d020b03d0118a775e24aabc3a617a0ddb38a2da1449fa31bc160cfe4720efbd32dca63b25bb52f5061fc664ffe9a01a8e95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5995867f5f9e2dc95c7f7e1dad55c9e3767504520d1b1bdf17f89a4fb11e7e40b1db93ed3962df352cf17419ad4c72ae7a72b2e0497575a672f995eff3ba978d489c690006bac3229ceab256eeef5236b3d806238f71258038f06d6183bf9ee9515e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ee01672546549c55ae0980d42974d76a7c65e9f9f137dc9eacfc6ce22acfcf8e4f121c3991d2b0116359b88e1c18ba8f8456fa48d3ff91edc2008f587cc2915d00882872337151257496875470c930507c03199c5080a0487267f46e1f50188fbcd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7e07688583cf94cbbe2d6bebffd962850dc7dfed0d449fd6aaf82738bf1b917ea6503216fb4a8cd95aefc63cf984211270fec506bc57434b4e68279c655fede08991f9ba9648ef578cb16e04f36e26230ae344642731e9739a02f76e517844ccfd5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha04afe8b4ec0f6ab0fee073ac2d13854543cecb3f04f1d7b42b238a2c70315d6379022fc5adca74def763917c6505800c74a0e50c9f2060a2d258f4eb5df59c22e87c53b5deacd73a9083b9dda922f8615b6245dff09ee064dd78433bcaf03f71c0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3de1b58b28fabe7a37f04ba3111792759b582f04151a12d1cd95b28b0d98af68cc3de441e448cd573b5463472933ae5db8258ba8d521cf14488e1c393446b9ef0a9d51af23d7365eea5cd7e3ed9a630dff8c0fc5ef62fa8e415ff7f776c30ba364ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6e87e4f2ef04e9675982f38f240c4daddaf18b8d8e442135d6a8a6bc2e711ae3c621236a83aeb4df4ae3f663a71ed179e266d18af25891662bfb32421e9d2e5e04cbefacb4a19e278052f56040a0fe87c8f1a6d31109e0e685694d137cb69b3a2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd49f650b6b09db0b59584e8635331e704e45cf01c1076e09f5e5a626edecdff5628332726e43ef60a7561f19349cff924e209e67bbfc3de5abcb2345975638df0e17b9fbb41de507eb65813473b86d04a10d06319f8f83b517aae1f699527154fd01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4316f038e0da81b6aa34f5fba79b4b905573cded7bafb9e599268d0c3516c076336327ec5b2b15d2c5eaf45d1911e01f8a6724222a7f84c7baf65eacd143abb5ec63f06ffeac3b3e48266680da6ee79e809da63d765b7daf230cb54b266da12e3b2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h814df5ee5857cc439af23ccd83e7b365e9dc5374e656053dada7a35c6534fa3379f9211ed86ddf8865307c7e2244b399ecca34e7a70cc1a750b1aaecac502afc7b85d6a2ad3b1d222eb259843c5aac35fccdc8207f6f1539715d85945ef36f9312e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ba72c35c0af675128f0f21262d4f6cbdc1b4ebe533d3dddc1aee6853e0e694379837923b732fed986d92165509cfe607e17de9f519422b8fac4ba557cb2a0dc05e9769bcce108d7886be7b8c89458b6f183afe71a4dceaec490737aa7ce3e4551d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14b8333908918f7b41a35a8da7e799a2fdc27e094eda46586512da5c8f0c5184da21a5214ec2ab8f09139cbb73b0fd137509fa9719165eb5300ddd19c309088543e34e868396d3117adf1c0ad68ba77137704a236cbcc69bff21c9bae5169389c8a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6770a19826c0aca1d7b4e2263c82279afc3d628dbfafed6d902a05e1cece9a1c1b43197761caa4e5f994797aee7011a6a7e80552163e129d5161dfbf5254c3afab0dee34fd18b76754049da269b001ea44ed47266990ba13cfdfde3cd31a54080338;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h323ba089054b9f194b1284b79e1a687071f4e796deeba73539372802e76823e1027e55d2f8b829d371d934250b629f23c042f260368108faba43ea1f4366f0a39418706f06f01cf9b66220311d80f47ee19ed1fa536b7b30177a4c9c4a9012ae08ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcb7f4f601eb9a0cc2bb923c386dc56da7478c97c7f0717713ffadab6a3a01ecc8c305c59f8ebc17e40c6739a3a9ea2c070eea51d66ad439ad11280eb8c846fba8d423df65e013f7dcd6c9979c908f9b5fa6482739ebe9ab72bcce7354b1465b0c57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf6f5ce8dac0200bb0f5f1c60f1cf514fe435609431e6cb5b64b3b92e6140deff40fe0c92eaff7e815024ad44fd94c284edcda15ef202542bfcf6e3a4a91b730447f84d11fcfe3d98d59944f505ed95b0a823f662d623d3d8b81586da5b13c882501;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he11680a48a6b33a320ce825d5724895a274baf73a598c93d381bf3802f2b95606b08ad4de284191099595da6afb8af13e46172c51500942b81f34682f906b0ed3ba5c2bd349316d21c6d65ef8a23788a6ead56c8d2e3e63a5f378c9e35ed5a9424f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99c357a5acb0fd0a358ec55e04fd433f7ce58f17f7403d35f65ad4d59d0551852fd6b458a80f0b5e8be20478532217e68dfe29535b618cc7d773ce3f73b5406f1f7530c91967185cb4d0c8ceb66febc6b577d79f8bf63bc36294f0476f7d98ffa374;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he16ef68aead76a717839dedf71c45a6be5387373908a9d854c8c30ddb9d1488091e3a56fa883b35d73aeb7c43e21c46e1fa251d7acaf4392686b9179ea5967ca3f1067198cacc4d053d2c9d24942cc650d06fc9d6f57a8512d0a81fd2f6f07810c98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba1c2ec96d491f6da1a882b2addd383c79b73c102c8989fd02f3d643f3ede5a974e9617b594248c7ec7785b31d4cb494fcb4424f9cd28c9f50378741ff5264104ea29c9ddbad8bc83fafb48a92dc4382364e2a2bc28d70df3210f0a2722e00f7f3ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dc451ecebae0297add83c675742a3a6a8b68efe7bb675de66103e8c0b508f9b6a3948efe66e74db5a44b2db597d3c9fc85d6e4966b8375c0ba6fcd73d4fa706b8d1071320aed25dd7e8ba96a01a4713c6e3bfe966cb743e339b6bd805c4aee3ca7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6874d486122e7c9d871584889b9017afafa0a133750c070ab7c834efeddf7cf3831d039f01fadd375eb7f1c167ade678b2f0f80407aba37c2a2019abf10f35d53e378a5fb32c7b492b3c52d74505b71f4bf3c1a83ecc959a80ced86827d5f4c2ba44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd89cbb7bb9b8a1ffb0998736d8e467320338a02b4aa2c141f9435b455abc79b6a9735519681ce3478bd023cbcb48816fa1a8d0be0a26c9a1e1bdae278dc37a8b8d1f0376e6c056bc1de9c37edd3d9150016e6b658f076204ebdf1357c08a55705b0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf02641729cce2bdf82061e8e33e87a106ca2398501426f0255dec98158690db14713b0ad12905be155b02bfb1af9323b3617589ccff11cd257c283615bb233755126bfc9538a3fcd8476d3eb8236519b21d1f33341d2de50b023b5442ea1b8ece012;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24f3c97dd8f0c3f1c6955e7a952723d176056e03f08e73d6c4765a244f5927e33f280310312c7f4c2d40643ff0b764d45d9013f1810e3f81f42b99ccf76c0522e125b001eb7e978c7a619e0846a50214450370ff95e654e81ccd6c3f0b6bdf7aeabd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77b305e34b403aaae76d20b256484e6a0e9be8e8e12673749f1f3dc045935544dab394a7f9e932095dbbb4a53cf09c7bb72c3fa5d2a6ad7396b6c92916231ca202eb2b690f1d3fa7b53ba6d2efa2eff0476678f70b5521eee0418cf09d41cda4b9fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h876798b663ae12bcf1aaa11dbe5b6a16d96bf5c08b084098b6b40af9d07034ef588a186b8f1dfa43b4f593febc951372ff126186cceac6a628b1bc76c14c519290c8585328fdc42eb4f184a040f6d5f1008b00790420784626fda73e222939bc371;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b7209980bfc9d5b323a3d96fee43c383f0c9eed7b4387bd7ed7757bc4cffb3f479f81b2c4c3df54905915390e27f37be9ecf786a27804d7d605e0395ac0d3ae56a15724eaa0040cb081308c773f68d68c1ebb973266d4248049fea782c98649271f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb6fbfa46fa08a0538fd44ae3511888bee5352562db3e8102cd711ae6e84d1ea5c933870afdc7d0128169e27f93c38d408cb51b5b2c44851a9120387b744f277e8d9e447c0300e6deb4db0f1265874da529fc299eb248eff80ffd5dbc4eaff2295f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b6a3875186e52384ca616474e659ff1eee4bb0d4670e07c90339eb52d4f60070c5b7605557d19d5a56f955c493385c4b65589e39b70d6274b91b62de0d466366d630a589953d1fba6abdfacad9d0629b11cba34d815bc109c10e32b1252ddd60e2b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3df4af0114b29f8056a37a1054211f92d327c40e790ea5479b865ca65743af75e24b0b243c70b9524d3f9d834a889692e47fca2e9ab9338a7ad229ec85a0abb6ec5837f0776286360b0e8a11d2e50394bf68115999db446c77b2e61776f9dea4a126;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc019f8e8e126e5dce616423790d8d7a26aa8e472c169fab09ba719dfbae195d38488838f7b9f7a680cb6f26774b947e0dd5ab075f17d1eb4cf5a81cea41555517bbcd926939334beaf4009f58e86fdb03222b1548327a8c49990803a8988e761485e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h119df6c73dabfe3baa9b1009f016e38b53bc392ca58fb9ed3cf785a82ec73da931ad637dcbae9f49f7b21c9ebe724d5038f7dd8fa4fab231fe4c610022f3ff00b1aa454fc6d2b5226554d9e6d510e3dc105dfcf2003b2deefefc083ebb7753cb9c49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5fbd5ff1eb07e7c67143e40136df75297d59ad83722e2743ef185e77b1187d923df301e8324883137305e24dbc74f796a88a8eebbf1d56319fd8c9c51e5287fe3018d343a8d81c24f56887f0d6ce41a5b6bca4836fa9ff1aebdcf61903e916c27aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d3475f6d6e8d968287d418a0225bcbe68fa76522d8e2aaa9c65d1242c33931a369ab3d89eecaefd8fd3265c805830bf9c9443e19efe59604e3e0f5abb3a2c28645771d99c88eed71c3939382613f97c23ec4db11b8b5971c09c6e88742718792c88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24d4df0c8cca92a1e5e46c044c187873f01f030b56635220976b3b5100932b85441ca40a79c0ed75f1b7a56b681f3eab009a59af3c78b1e208af9372c38613ac75dd8281c9a09a11ca04590573fc547620c6a6c3de5a21cc1e7c03d075d49edd038e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ea9981e6515b7335a14ea21695a888fcab0e06ee7fd090ce497ae65884f69715eb1177310a3941b156863b9ca3de89f532ff03f93aefaad235f6a0959b175d728222fc9f06a15fe58b2ee2c5f1ad24f2854b4ef7a87501c0dc8f5fd20383dfb8959;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1d69a0a465682388968cac8df9ee32230b1835a9aad7b270bcfa350a45132411725c88f74c60e455c950ee45d2249f72013edd0ddc2d6a0590f15a4b9e77f599f773e42be10ca3d072c7a69b7b4d59b175acf8a65b217a8a2ed81d6f1ef5cb9edf2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd813d6d720eabe37bcdd41385d5812f03e01cb7453dd50593ac5569231b160181c2a6456dab6a7ff9f36012835e4c638f3feb5a4ad85fcf77844c68d9bc83a4e6f0d0dc9cc684c978a32a13d96c4881738a3752742e44365a1592351a799aab0f4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2cf6d3ec72728a1590190abbd0f522e000df1c2f3091e9b0b78a303b0bb84fa06670438476fa5b8d9af2a2936f5d73494a5c8383a52a88a501f1d89c1c0ee2acd56672bdf8e2a90618ee2e2fceac6b94b25ee652d20d225e2808ab4e1afbc74c1b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd06210776db6a24da5586a67ebdd7348dbb44557f87700b977e6fd094ed29a9780dfe6548123b3889fca438da7d3cc634fdf1d00077d4726ea2d0c835ed79e50ed6951e86d5ef28c1afc67c50d26a7fdb471788e424c72111645f22b8607ebcf121f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7d06d08e1145bfbb4114e1d9dffd2e1b3d17626af3585fc0072814d9670c88d2ef1feaa9d7b8d2d8ac77337d7e62b1881dba436f85639544b4313ff42d90b8b99d33b0fff1dd0e835acc496e4f1ecf193ca31ef4a3c72004562a7f4adda9922be56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c89ac5314f448bd642c43cffe0d6e03a45db9c2f013b57dd59b18a3398ba1279d818ca8961fc9e9fa74278f138cb6bff3793ef9b576febcc73135d5cc1433dee4765a1c14566a4fc01384d0b8312b227a3b5603f927b5338849defe31c6e1d06dde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h404abd07753596a26d0fdf4c5db41b69511228bbe4e42f2cbe9461894e3bb50b7a6eea54da63323c5420b01b9879e0f4fec9d14f5d3df90766b4e57def04b7724d1cdf6517b9c0f2cc321f2ebcfa51e6f0bf85275a73a63495e440911d8e8ee10673;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93aec5689adc640d5cf35b7ccbb614c282d8345b684d153880e9e8742dc349926bd9478adc0f9eee6c3aa53bfdf33ce7ee84f035a2ec0dfed3cc7f07caadc7a92b45639f982379fddf16c07b2f3351dfb50c7ed75299ee7f8d02570cc85701ce8792;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha712c2cd402db607d4dbb09aa35eb59dbdccb9dc02d147c10faa7d971ea41e75b720495bbad70d7ae734c0442ce2ea3377262bcb9d3609c78791df0677d6b463fe6c904403a1d87aebf337022a4e720a9320a74b526b696a19202812be6bb403afcc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef6ad231916b9b76cd7dbcfbbc14320fe4143053d87226c8d2d206185155d2333e562d479bf0fd8fa9dc508ceab89e98acb6db3bbc409c9e403a41d5d4b94b561ecca8d833e5c2572aae63a2e9be647bb4c9a0f44d27776aecf45c00905900633e0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd20554095e4c411a06c1e4931ae164e9ada4860ebb2d63e65b38478f9bcdf178b54f8b6ac4dabffb337f2b137394248db249f98042eefe9a9b772bb635ca07e994e52a4a8c901fd0f3a94cb9b6f11776e04a49ea6e3f2b63f7ea1c7f6e8e46505be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haba0ea30333bb75072a50a22e7bad034ed48791f2a9e6e08dd929f9ffa912df4c18962a9bf1ee41e3a915f7e35c0618ceb5a0f0d8ee1cf41b2744ceaabf1dd026b6744d9142e873f65c7f789731f6ecfe7ea25b225b6248d8047c099410677371799;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h887a5c3bdc9040001c01d0a56ea0e615bfe0d852305e678a1f8cfbb2e8971c7f61f3f159883541e3aef715f6b594f150caf08f67c76ff73c5c94bca332faa5958c58e3ff0f9e3e060fa74741e5290c05450a369656ae9df4ead23e2127200e9add01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58e418ad09e8e9fe4e44ce8e7b4aa5ca2176adefe150a230daf192a81dffa59ae00aa02b37e0a1918228686a55889442bd6e0207addc1a42f906b1ee615ca4b84b279a2e4b7deb592010c13401fa51102bdad9b7d2f27d411284540a389fb7b0ea14;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0c83148722688933e1b52dbe1ed9f685fb8e3ba68cd195071498ef8c65453ba3c8c3c420b0109bc5267bd84e7d5946a2a35c6a6183437543b3f026031d1cb09f0d927f7aae649e1eade1f54343282db4a160aa054efcf1f49e3a140b3c81be232e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5360eae9eecd3b2b63464a6fc7480dbdcece679c072c0805f3011948678b9ecb2f3703315cbcd56d62b5becc486eb284c885dbe2692d017b34ae5a5e11f6ea83cf78f0b3c167e1e795fe317b04af305b1d86a8a06897e9249c60e38a354dcbc8ca86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb2f0ae9ea0046449ba0ef8e35131ba3492ad00c9eca5e1a9029297187c07a35fec9b52fd0ddc4860c28d2189bec68bf18af9b992f54b54704e9ef1b1edbadeba9554d545e977900cac952216c2f5368ff87d7ea51079d1fbc3a9ca4a559a4239c6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2c982b1cbe5760ceaefcbcb7ae05224cb77ae1d0facc4d94723dd600e503e2d348cd219f51ede1a397adaf22d7c79b1bd372f39c9aa9bf0892e242dfb9444a0b5bb7bb5e8f3ecae83243bc2daaf1199ec6db1a14679aa40829937600fdf2a08bab6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3251a74003ad7fe60be04c72569825501abb8992e1a5cd341fe3468e83a1204e383c2fd53c0b4b795dd3a5d9a8efc724f352dcef1abf47035230dbe7bec3bbdf3add1e5463c580dcf7f998e6dea9ac1cbfd928c54246bf1f5c390c9c7387079bc18;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cdf814aeb941d108526deb7abd80e813dfe80edf06f02fe2c3684bd592d6ef2eb39ce91d1312eb2f6c2c732635d0982bbd0392bed9e188fdf2a9e14542330b86f9f89219d9595edb7d880a423c048f4f257af1058ee195785bfc0a62af55a124c6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28bea13aa6bc03b008d691ae63a453e53cc7bb07bb40f92106a15b39de015ce77e9c7a75f0cdab19fb60184201646fcb3d47de9837a7f569ada5609735aa51bb22f3b6d6f1877573eba01e54ffd27ef9f5453bfa4b13cf625bd70202dd00ae63be3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16ad51860b6119b47c3fba6678a7c047e889f64d8fbf747421bb6fbd16f2821b87c8b1fad6061f19566a166f5e517e525237cecc67325ced84f25f3fd8fd7d63e137c30972fc8c95ebac13b94ea43b30fe74b090627d607aa6658922047b807fdb1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9aebcbc5ff6501c260ce3dd3ca72d826a90d5b5fec11fee5ea1bb5355003d85219994364e6e4028bcb2b6645a3d4b558300b56df9644528bb6645b09e2104bb0253f2837e97e67f2de6aa97394a274e8bb7517bafe787a3d1a2b9a436c284c82ef38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e8f9d9f8f6b6d98b881fd49dc2e00e083c3bc3349b7621db065a111a3f0735fb6f005bfa21440194c8ffb48fbf9aaae3bcfb8b704ef71662a09994aad9902d7fb73bdb366c92db809b5a614fc29ce13056114dbe9762c6a5e30c3fd0a6d2f657c81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd57cb9c20b9428de27aa08f55f26fc6b775a3f986392c7c17d10ddef0885c54d507767ddfd16e43b3479bc1cecb530aebb1932fc00ca5d56e79cd9dfcb6819ef4af5038208190c614940c36635551b069e7309df104c0b45dd284a82e2187a56c17a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cb5adf6d6d53b450ccf7f267263779b9bc8002d49e688c36583c6f969d2fb392ed8b5e896b3f87088cf7494770236e6d66cdfedfdc0f9b6f3ae43f684aff9d94dec184e1e6afb088ff7dec470fc434bbd8b6ee5e5232f32135280e40529ca0b25c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ae82b370a270a6c8adb8971c46916e3ebdfe424ac0c4bfb95a7e8c2337211d435c4ac5cbcfe0ccffe66018ae76b2df61f92fdb51b91dcaab4f9d7fbababdd876db7016ac26ff58a5f972ffb116f8b889c603091584a8aa87a478de3946d89397c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ff8f4bd819e073ab20121cdaf451f5869540e86d515e0b9f49b3c1878324e64154f435be5aac73c7b63c337fc56fde69f2cba829379e2c652b678b173ab8afae6c1c0b62671a3e3941cb28c89a8202babcbd7fcc07a3174e2e699ac522256f66662;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c42820dcbb8866aaa7e4572c8031acaded4b903ad6f5a3df5973016b6754e4720fc7e202d8798f5c9b6ade3bfae13d3d07aab48ad36410ceb5f568e584a98ecc3039673bc402026c559801e953733ed1688bf2255f9653ae6d849ba75ce522028a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d7c4b6a68328a7be82fd3ec76413a1a3b5b43e7e34cf8450900d4d3ab8f641e252c80ffd6630203809315a218d7e5e5b887fb4266cae2c6073262a6f773843f12d15de2f73369117313a47469719dbe34ee0fabee8966365807a51317b658f2d0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h935507942fe3226d1c3bf2a20b3e753e9ab79a5350f795511ae08af154fe311a5f1530874eec0ab72e47c2285d25a45f778a98d9f4b3229362db80c92c0006c44c00a4f039a4651dde16d92d7070e448f65d28f9a8d5cdbef462ccb8b8c716ca06f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h768fa5b64e14a782161be73f24874f27982a42e27da0a1733ff33eb579e4ea1b70f70a2f1b874d751c0ab7a26a6c1b43ce579ec96f9b0b6e8d990030b869055d300c4dbb251ce9f266645b2cf3d1b5cd8fe68c88943f0def0fd542de3a3799bf16a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39f8476c313e49c0daf9287e2c4636d2ec9a07989917ffe987c8cc08cf9e84f134efc52f92c36cc59d205349ffd95c0a0f7347d7b2a95eb93b797f3efc2110f7b3e69f3e831e14b58f9ea29dbd653c311f686a4cd181270bbe84e054e5a78748ebfb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3712974107b3a0840d82a9c2ef2ef256f0f356654fa320dcc1141eca2f1f2fc1892825578c043029c694958b88446f63eef51670301e774a06563a45180f200343ff895b4cc13ec8ccf80aad763cabfd6353653e2de18f5bcf1cb44cd369fd0ba3f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ed544292faf6951848c30189116b7ca30ad3bd7032c09e8937c146a39e7a1f227ef5baed53db0fedf4b99dd1029841d75fbba17134f3f6c200b9e99c3f05eeb211ca68fac3d8cb9e25c49669b24f77b77da3e0d86c4104a2d9a1e98f43b4263e60e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67b1a7c7028e747720ddb911431363f6076159bb19d03db08d691dc2a1e1e821d9ae123debd10488e03fc075000011cff07c5cfca50fbb834e09c512a2d73a5288edfd4bcf6dfcf2c4830f7d8c19025719964f4aefcdee17897e81f3c66b619223e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf1802d44e6b477b72228b6f5ba1ae905610a42780617b0cfce1605998baa98654397f93e03ce60eb086f8185faa05ea463e8cd5f715d9d253ada60ba74a7edca67b48040022320fd4a8af7194d8a4f3afc4c89d410672c4cd5dd991735bb9babcd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c202158add66d7a2af56f037f6e36cad73ad45facd87926b5dfcbdd8fc6aeabeb5c1762d21363339d4c4c9ab83f6acd19d8b4d5c5bab3ef6a27e6f19a8ddcf787cbc1adfb8589db2ff242be0610fd7ce056cc6fcdad00b6fe293d0384d23b818aed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e2015092134807870f5e95f9e094cad1c267766559c5d29f9633a847696981e2c097ca4123de1ddadc6b40aa1f78888ee112eb1a8c2685fdb96c736fdfda27447f8e95a24991fa4287b71613087c702a9d6ca6d5f9273b81cc504ddc896f7838475;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20a913c7c8ddc56af750d52c47b15261a6cb04b43b94588c72aba9ce610dce0dd7907d4821300cfe0637d4629d942efeb96b2b7aff44e57976b434a3c1ed9363bcd67af0d651446f40ba536fba2c5e93db3d3284f8b806ccbea3cf78fbdb51f54e47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hceff643b00cb1f7ae16ba3f72c9209e03e194eadf190a61150255c728030662195a47bea94118f6a26a432d510708afdfac6c47eeb1d8fb93382a4c84528a89d0110c3c81aa143bed968f0e3070cc9f9029fbf9c74505ade3c5728b0e71c6edb1148;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3a7e906b394c97da02629e26d8ab1f01bd94206c641fec933e1724504f753ceafb6e006a99b2df0d85885f5b33a567e5c6043d78c2a72bd3abe902e2c2af5d50a5e170d54fd20879d091093737a1f24da8f4f49a069ec6d5edac1bdeaff67eae410;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76697d40b7248ff8e73b7be41f001b1b9c6de44221dca1abe6db7ef84ceefe2301f4c3aedeec0efb86dd6b44343583497bd16f09f6710e24d5c1a895ae9f13aed548e6510bd0da88439bec7bc8163f893a12505d0c084a19c3e7631d133a05c7f22d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf80f52d0150934b408e37a5443961f7a9ba85ed2cba0377553ba3327de24c1dfed11c2ef2d544c1a1d3004549861a5f568fe459db627dad36bdd8be8ef0019f405b9cedd2f7af17046c6f8f58536379eb3f5163c6e4c5baed05313c3cb9f6803e9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22970bcbbeb209bff096c3f6b93406de7e18203ded39a677e4b47ae645e3b3a87fc25669f06a5815220d25c31dd329707e8aa265aab3f749fd5dfa6a02d3c20897cc9fdc51060aeeba62211c86387a907e3eb78d801e4de074a5517fb87c5d1e769;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h683db2b745fb12e7c057afa6f919069179f91e0e74597bd05c82f3434348ea12b86b07cfd32ba60b7cc930bab78f8e2dc52806d95a0d7e06956798a361fae0f1008ff04a75bfb7f05987ec74d1ad07d72bd25137ebe19aff9e6937a55a4d87101b12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e506cdf82107d28317298315b96d08425a7b7711ffb1973f781e77e20a7279cfe4fadc436db7fcae04f438ea840e12fe11684e3284a6397651213af5d7c9bde6f943616af695f0e654de27811e93cfd611e28f198c425138d8bb0b3118a12dae284;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb465fa77aebec73b9cc598b4c0ef68761a91ad6d4749c002384d5d15ac56ea6cef0af869cdd87e7da62b09ea936d4427b9ab49fa9eb770f0b44a51298d4044cb167172a66f6088b3b4d1a89f9816a6478a5159f1b151c7e4faf17e6ccd657e337bce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce7ec6c252be522e7caf2225291b70aaccae853d022e5299e1c4f73063404ff5f3b9491814c3dbebe6c07fd26355f8fd6448a2581978c3561943c1611db2b33ad777458c7e2640b68f8a30b3d2b528dbf8218454515e00fe194669225e750db1efa3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h485394a48770d614398628a712ab074088aadbbdf94aaa2f76e049caf5ddab242ddf08db2b5a396d9dd0016a8ecdeec925b9f9a74c1fd213451c469af0b17880332509345d1e473f876b5526e0bcac1a6eda3f953681571c8f2f3925db375b20f2b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf610b53b508b818e75b4796bacb685e91e1bf7e7f6b2b99ea1dbfa3566a3b6f77939185c83abec2015ce2236a521673984ed8d3affc335c4da965079b6bcae5285e6ab59348eb4b71b0e3d56a976be74f929ae36879523d22808bfe38ed6fb1cbf12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4444b0664d7c8dd0b4ba2b2e018d96ad8cbc6ddfb3a1616298955ccfb076a1c8dc59640b02268902c5e0c3efbb89de4db3d09b193f32ec486f2861189cbac9eac6dfd9a3efcd2ea0bd21444ecd6823ff1083c0b10b7d545e1b0ce614b42d12ce1cca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1815b435dd141a1704aec9a2a8b5e6a5a15b865557e971753c646937c1c94e4337673649125172513dc5a4cf65b025287650d5f288a04790185c6783dcab2b571aeb536fe680dc3fb23cf6dc11d05f64535125a6e7e45876f3198f50523b1608ab0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ff5f19cf81cda8a7379f86b024b991b3b76bfe58aeb578b6f99436d4c867eede33eee361d22e2c4073bd0ff2ac88360f0184efaea5e3584320b80ad2921ae6d131eb4f974c99c5ec2ba5d1f224d1b49a8a7cb6a787f930db708cb5735b063043191;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd93940c6c11397d936419f00be46e71730a4c3e954a678b71c2b91209d9d23e711e3e5c8aa30619b1aea9bc31997ade7b59c34b823ec74480c6eff6832f1f6b1551781bf941ac63d7b1907c59ac7e51c2d54444a2fc0846c6a3be6a3ccbd6b01b38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4f66e6c3741f5ae2e43b95296e08d75dbcc8b9436fa975734d8b17e4f336135767c4deb1ab243b2999d645f9f1f0463415700a5355320ecbe2877c313a9877cdc6702149c1e9b76c684c80f3717d57fefac722749ffe1b3a7e6b05d9750928a520;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbfa0c914ea979030f554514a96d35eb8ebfa9aa5b217f9e969d8f58356c3e2653d66b9c5de7b68b7fa223dde52947c385b71cdd7234d1075d8d5b88d210cb3f14c56504c0d77b1f8be8b57fc8aab097f36aadba8fa611d17de05037a454e94f3c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb3cebdc487d0595c2d71aaedcf2379eb5307c88a27ce127881b401bacd8f6443cf06d25a6498084cd7f5c5d67893d48478566aca0f85577fbe08d70a5c785c48c7f18a008e31d471ac00132395bb8ed085b26fb403218355477c28ad7abd6b6ad90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d37d0b1b1130a63c646be5cb06eb8b12b7c3c49b339319cc25b02b0662f099c173342297ea38fb2786e24c1df0e16e71c30ae2d1d57fa83a0748868c1a24172128b7d73d3879d86c2ad84c0f0b97e11ead78a045e35ef3354c6b493ca069abe48d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4d851ef6c187de4b23e25d5f88583978d750f2f3313fd12ab32fe0d70c8c591f5af20bd76c1b3a7a113794abd8ee9b67da996391cb9ddbea7ba08e1dbe11cf1df50b74828f378584041e3b758322c53ef5f2bdd4e04addd55aff494cede709f618;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e2223fdf68d8ff1f657cb7e843c2b54737fbb3b91395b516aa7a3730d4eefe292bd360ff1346f28999781a33de3d5f389bf1cfe4ecb1f613064f195ea2d095968ab65ee18bceba0cca6fc0fb5e88d1aa2ad972727f8d7e0d4d0f6d963b71c186c12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39e828431938f57513ffff682049b4a0664c16bc1e5426815ddfca5cb5da7abdf301529330932fe7cab291d8e14c8b33197ba0134a5201aa04bf867205cb867303ed9c5e8e1a1a9c34b7ab24d5668504691040a4263b26931b67bb8248a3d2f07719;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb21823ff8d5f64e16517abab51252eefef3e2bf972331113412944e7ab11f6c303940ae92481f602834291eddc993dc341f720984c8f86c9766452c7a514efbd885c33cc09618105f6fe43b0486d363de7239326056740e17eee75845ae97a391509;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39186f895cff2b46e111803cc0d923cce0ada63a66e0a82b5dd5d7fd1873d82abba3aa6909552d57f976167a0ba064e5dd4bc9f43abb5038088f23b8211c1ea3ae3f6568e6363542696609a4a572c13e2d0c880d0a8b4869ef359e66f73cf1326a23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86fdf170c601e82539649e89fdf7ab5346436b511b3254f80d8364801994619125e457c55e4c0e8a8a5f8a1047ce219a5fb061f8fddd1c389ebc5499d28c7b016a947a74aa2febe0ebed31427df19c5f6a6c56dde35dad3fd32dab1f4573d23b53d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15d97ab4f9dc07ebbe3dac95aa6e799bcce9c70da9447dbc70c1e1e6d6d3499a278c5d54dc2d6ec7e8031a9132dd58c7cd0a5dc8dfd4243c67b5d5e49b48dceb1f615fb79bc5cd27e6be21dd50832da188249d8747c10b22388140be100493e90aa7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h250919a1ed0ba285a161a103bab99d0b14c869abad417ad8386673c329d87d74938d94b6f3783eef2655321619371fdd7e81e8286bb0a4af3c525513ef980a8f7d073dbb35616cc3ecf8522f1cfe307097c295acdc677b1be8d0b520261aca90d5a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e7fd177696432377d16fdc9a3f678cbf554ec98c0f7ec8de22c2d8a16a0c5064f77de03deb304f170fbf296af0826a3cd1f23b6fd2cdd688d0a316b07ab50ee25eeac2eaa3271d41e3b643e4468822681ceffd49762fac8f6501f49faf2799c9227;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cfc39081b6edf106271eb6b088c2444d51c269a526540cc68351d40b6ebbb937736cac6c5136ad65397747a5ea3c13f1686e2131d049999e8adeef5eb95db6c405243b709d220843361727d72e43feab939cbd93eea08ba1bb84c396b9a3f75b751;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1096fc64e5d6df09c81f4d9614b09d9aa6d675de3e5fa430b65dcb9fe05878cb54f887f169ede81671a1201096ea68cb328754cf21f2cbd71cd808aecafdd4ecae8823562b79aa47a924affb5908e58a181d18b8d9738f3532eb017181d4adf74614;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ff646934fc55e2cc29851658b167d574451ac42357209bedde3f588757aa6f21d4204f08c1d2edcf7711776f983cfd34f328a1a4363918f4d08500da95d8283e5464a7aa1742d2a1961477872f55d05a0ce27876a93e5df9275aa4377997a0c4acb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c05e60662bbfff90fc71cff563e6c218099623b3c22377f55a29fcc63e649666d214d4f55ea444143b53d96457935b3d8ddd1402e199bf4b1ab3952a579ccddef125a4b0f2e0cbc37718746ef0ffc1f117a033404a42b815af61f716dd6902198c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0b9e4d92ae98d8bc05dc4505bf9945655a347959d856c19097ae478eb0e0ef81c3b6e3b32b7a918a5caa331143d6ead9ba5370b6c664365a89f7696aafa9347793d8e2bea1a229f149336dd61a47cc122e19b97ff10d2e87e3186ad8222c23a32ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78e686d9a2dcadedbc35510a6355540a11bfefd408fb1343341b696c3408bf2c905a9b69ba4d67ae95398bd87869a8b7d0223e7f8b570ea00d38e31ccb85e5def9961f8d56b1114a75345f1751f2879b785109aad4a19bcc5fc1b91ae3ded5000d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb34ddef57ce2784e6206d6feb2ed926e482aa54d42d93fd1c0a1302867b0f52d6a1cfc4d56294a168610ce13397c41e95e8f0072bd2414686fe87c43cb051c6ca82da88c8655ed9cfe0d7543e02f6a67f150879810205fa03bc35a515ffe0967c8ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52aaf69a485a01eb91e55f7792931405f17a8dffaf048f95581beabff3e2aac98ff90ba307a16e7de106bee43a2f21000732e7893480829920a6635c46f104a9d8007172581dfdfbda800b1caeb72da23ae861fc75e5881f565e11a1c89d247d1b6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2e9d279d25c8fac975f0a2026c2af43c2f068fc7be7a1f024faf1f15a67a1ba1a2876004bbb904170549ed90070915515f8681cbbd3c5f05181b4dcef7712b0a0b7d35eb03442ba758ace6536db1e96b4efb348e7f9cfa11dcf8f7333306866ced5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h500bd1eb13d021acf78f783dcd737cfc256140c3a31e88dcbd7fb7f7132766bab40f5f7ea753f534a05a95032497a76a5401e2452d218dcc79526b8e831d13f92b92a9449ddf5ece4dc9fc66eca8a82dbc045c80cae101552f0b38e247a12573e14d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93867e2af23c24648e576cfea0d64136b7ba06a4c3f97f636027e78613c33535bf8e818316e4408e801ca1ddcbd8fc98f9aab15cfd741ce03fe0eced202d0d2d9ab48a463b37f24af1aede16e68b3a235777f2c5c2c72f852a66783347c22f66a68b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ac491a0ee9fad87dc6715f941ca12067aef031ef3d57c238385c2f8710b9b6061732b2ef59a1fa37269b2e4de927df92337aeba51e7061d98c32537fc0599a377e2aa7aa9a482a30a092ee6750ad0d758f440dd85f6e460a2578682fd4a13ee735a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d2ea41e2542292682cb4a2f7f8ed51300312e9b7083f0c7803afcf6025d52ae91dd0be13ac163e0487602d060fd3078f5e76f10a591bdcdf737d0887313358b1946e6ddf747a71d627781b77ef5ef1c8bd0fa54fb6db55bc73f0555f14d372ae855;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfd9aed8f60f4dc59710d351ece946bc03bdc159ab367b1d3d430a014ef368b227ffaaaf4686003a774a602f9bff3d118167b10c11b18084a01006a1b695d4365b3f36e2e7abbf65f11461b4fb64915d07cff3f2f4744187e0f4d0c043d244c4b3dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2c2e242eb2e7599792773a7b09306adda17faabb6a8ed3bfb888b27fbf72601699755b70619cec0302136987073fbfae9d6589b8cc9fdc1a25591811603bc819cea30a7a53c3ec111fe5970529884c6fb7a80c013911765906f4c62f68e41643dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50290d410de205ee9a92f2dcec412dae682f7ddd2614c367ae82c301b36e7a2b6e354de5899508a76a09b76b5fa3a6f69d9ad545ddcf5a0bc8c6fe87392078b21f01a6e55769acc8d3cb2f720f31578745c2488f7c7044f9a209ab4f9f36f0a4a3c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5636839ce7ea45273a43fc676a399d86839e0ed842ba290d54028e6802afe5d2a78d31901a8eec14da76be8905182552ab26a6a95913c7b8f2bb2ffa7bea0f4702986be89592ab343d08b428f209445fc40cf6c73d2a7bad29bef2d1c565ba697fcd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcda747c42c251f6c1bc77b0b6aebc074112bc7c92250b37b767e6f6215834114f6a2aaf2433b3ba798df066ce88a0553dfb65d3cbf10805feeea0e6f9ac2d4355b40581b612277f51424165602cef01da1b931cdb94fd97e7e3881cc6c6d11201cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1a2a0efb2775320e0390b0ae7274a5b5daebc7f720474b2583f331716432f85e6f1987604361ddb32527f0db115436e252de90449d0e84310ca4a7dde75d5228d0015292486db4ecd0de58013ee530925f11eb1290a83a4907dac7ff8de94354271;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46fb9ce5c57d4905b7bd37a7515c8e635586aafab2bd05369bc0005e7550803dd66a1d46820c8f9da8794b0b892aa1291c873049ce2d765d9188610eb4bc3854d66dfaa8deac77e5f4447276d8145f21b71d1683b90585dd7e88ae67a78eea41effb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd86ec25bd87bf02d64fb9895a597fcc5350fbc2a93c8916a736cfdc7a0c4c534ddc683681855487eb580575f2081b722d2df76f73214bed184565f37c1b18dbaeb976504959bf708e3dd58b60826e668dd047078e10dbebe174e7e04cbdeb8f4e008;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84f7a54030851041a91aaff748ab73eb8085c47df0e62d0cf589be59ef9576d9898c2f99eeaa9169db4ed76f8ea22cb0ac78516a6d8e9d179510e8b63cf3c9960bc1fe6eca6da2d646d628788cfce364569bdd5f4b9140b1fac90314ccbf97027da3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40093240d7950dc8900772a1edb221676e9ebd35a3626d0d50ab4b2a6a8131f10dc4334944d00a4da5aa20586f7ea6bc280dbfff0cb017904fa5f17bd4c84254723bbece6c44d3e1310d17c231a855b6e92f059346b8d08fdec7d722bf70ecf002d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6209a29fb918722f28d11e803dfa615b0e25df8a97f698132c5402d4d552788cbd027a09c01269345af455ca90140f846c557bb018247c9da308e7f5f5d105ac185c104e32833361363cff2c22d0fe12ff86e1c9d0ef3f544355c86c492b9d397e9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7601935f4706c4410b45dbcc65e59aa5c6f89fe87f9aa5d3c2085efcd589436bc871e35dae5e0c5d772188e7d55dfae6b899a3b28aa1d32af0f3923cde47ba501dcb7ecf77312f618550ebd643f88e8da645b98217527485ddadcac8fe224905e56b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf96f6e430312bce42cf0d477613c3cb8311474be3ca9c3fa5a3e9a85aa40b9bbc5a6b9745d9a16f5e50ecc90a6e51c34a47a4e7fa75deab332bd9fe9856626f5ca79e788b325b0a3e2c784d628812051a64fcbb146266ccb887a3cd36aa1073f9954;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3053596c83445b32324a3cc27cee52636faac22d8176217ce5e89d7c4fe3a740c3123cb75ef0b032777d0d44cca88014584dfcd2341d0f243008c59bb67b42b00a6aab4d2958cc57be1199fd463341c9f4af8e7a54e1e583588c919f428fcc1ed7d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb07c7aac7bbf8464bd17e33f8216dc4a8baedf93c0f7b4ddd42a48d1059f22e48574558df545af12eff1f1178029e5bd2b271684644549560b8e24604c344b4bb8923c51ee841859c6fe595bd47b6d8fc4360227dcf840c4387508ee09ed0ab2743d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20c1e187fb2adc48f9eb795c40b913d2c165037f76d549031e0f11513a4124892a349d46bcaa718fe13e1022711ecb0fcb7013f0c9437a84cfbb87b04a80fcd252bb123aac8ee96c7404de6417ed166ac635f326bdf50710df66c8e5128dce890481;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc62e6087ccc57b8a7c59de83ed1a75eff8c266f11c3378492efa9959eadb2ee02c1daa12bad08addf5b4f759885265172252f8cd5a5e39f7e43d8aa92971c8a73a33605dfdcf8b87a1d8016d6fffbb54cb5b6fd3e5be09e5ff805be4a98c0e481554;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe24838ce180f63edf9e963ca1c9ca5fbfd33fe0e67cc0d0030320338181ba57c9a347974a422d85ea80355996ceddd9f59439ed1658fe1a6ba267790cd46321e2e42d3d79fe98213a83feb83233107219b66073e04b3642dbaaa1271ddb40cf298f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68250f1d0ece2fde73ef016a14b769fa0a097d7ee5ed0dc8837c436cda94f97a47a26d76c5fff19c882bba69adb698228e56c4fe2657234040323cc14928e065c070d901a102334dd2b4a8942f6c6a26305f2befd8233aa25319d35db914e8ceabdd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11843bf769b01b50d557691c9a286146a4d732af911025935bebe27eae403fe2b01aa9811c2b82f3f0cecfef3d82621ee8eb021a35c97b37300047422f14768b3ba1167da91ba0cef65914b1a3c19f2011d201cd043b15adea1c3e57259e914384c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf36ef77c34d3ac067b6e3d086185823149f3ba60ab11e43fa9dd85c76e6a4b463381399c2f7bff2fd7dde7fda55adcbf6ff2d38d75a32e11c7f0d86157ae347eff91a5b045af5dcba5dbb1da77d25f469f409d764620119e94d10372424ee44d01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h368b7d3cd7b2fb6c8b83d22bc5f13355a0644add11a61cb467d50f621d80dde97a9dd9444151fc57cb0cda5e52a6efb81451e2caf74204e3b68131256ce614bd28f050f22ae76ff0e6092f8163341c15426f8c5ed579f0008dc193bc6f77562c6530;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49996696a751997e293456c9612f1607a838b364e39b83a308bb93eece633ac985dc72cc60a16e39af176fdae4a9a9008e4ccd178a0a41ddc25c55edcf05e298239c675cfdbf5341cd19006139e8ed708f26561c30ab5ea7f6d31de127f59050c38a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8aac07fa0a80e1179beb7b35853f594c29cfb6844aa2303093ff07d16209d755b355a36afb696776d2831e3ec163ea7e52ee7239d0022f489c030ab699f79e68c30691853e5e9506e6ae8141ce19156b6f4c8f557c92e8c161c66c223170bced57b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb134e3ceee0e84c146bc86f982a6f98a286949dde95a62ef47f1cfcb84a56650e23d232d4b2648bda9a5600baccc00cbf25a985714b89018dac5388405c082ecc7fff8add8c4365e52936115cde6139483ec0b31f4fe992690063fc1598dda58ce8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40e51d886a9c1237ebcf4b9739aa9c62c851ec9523b3210e9ecba9487fe29e7870e570465adbcf2a1328362597db82a6b9d85384b19a0e9d1f469e1ee661c54dc4eed261b433355a6d7d55c2e9eac712d83846e5371b5251d09cc41fc71aad74506f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec62602bdcbdc35f386852867755b1b78c5d8381c78d11225460a461151a13399f09add366d28784aa45d27b7b12c1292dabb96a13fca9154a070d01883c09e1688f341cd95820862acb89cdcb91e1a52f4687b51a2ca334b81342d8ebc923f5763f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2a5c989f57b4d17860d2cd830ad8dd8b368faf040d9419331f064af1ee07c5cc780f2ac7092898225c003808d01c47ca062de9ed66329636deb625f871c3ede285a0c6f0b3a248d0babc88e35702ebd81e1c884d3b3a0ba9452e97a708786a76a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb64e92e7263ecfede8c2f97f547d252cd58cd9dd26e4d58dfe66d4ae284342e2afc9b3fead8d3b4eb0ea53df32f9352b167cfc20c87959f2a96d13a650c119fc0c68ef2793638a098011e8e94c35324949dfafce43f98b607ad60d9edef295f8384e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeb53dcce0a257d3f324f1cb75250a694d674d58c4d7b911e067719277ef033f8cb64d5e1264ddb697ba71b2b0316e4c47db67adef24e680e154b9bcbdd3986943cf2dce8a67a8aea17d2a133b686de4479dd8be4be7519c115516d87e96eb67e6d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4800f7b7d6ebd2d28913608c9964d9cf727b4b2814d4eabbe614b8c07ad14d436431edca7fa6a90bbc029e5cd4e44b5953f604fb9186e5c7964cc1799d5d161e25bc6ec450ea1d6eb137f873c041605e78626daf4e1afcc49a99eb953c9d02bb87c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he97a3e8c70e922d4048f675df68f500f3aa1dd3be30abf13e352d08afec567343b0d951da967798685f7450120b2a014b6a3f19f1243a817726a7e6f3d0cea8f13bea86ec426cec16f55d72c0ede6838593bfbe3f2c8a384ad30bc3769976eb956b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94b663a2a495550b7ff4ae736e005be3aadd0884981a4bd790a93ae2fd5a6a979236aadea66c79484f725ad9ca235a8ef2d419b80cb09e44a6e9a5b65c88c0ce09ce5b092a082d7e47afd181c104adb1300fb306b5dd6321e3847bf8fdfca7dc3ae7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6005a6504b771353f3842b010edb6448240e08ad25561a151ec0f5ca39dd72a56cc0e214810be8b92a0facdf99f867e3794b239445830e327e5b7b1b26be746a6bc5e019e15d40a092b00a7d17b060aab5ad43217a2a24ca1fa1742926c402e0e2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37e78704d9de1c65abf26b93a7f4f590bee9de2407fabfc7645b795bda42474c81ba4053ec3900bd9c956a9eb147cceb6318fbab4b078e14fad85dfa84a28ef442ec9bb5a92bdd13122ffda8c999903eee767f8ef705eff8961d40c3fef5e61284ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58f319b38bc59ed6b1249b5034b59f52c2add6c3ce8177664e2f63fcffa9f31afee5248deb32b3330bcd76ec61ab7b7262502d4da9c0ef071df018c0a2ef51f6d81432f8574d1afb4a2c3ac232429fb83c5463d096bab756df9734ca125433e13ff5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6712b80e06a69282b33edc28eb53e0f967d15e58ac73afe90e7ad5ab45080ef76e3256ce41d20030133894b5d0bc4437a50b227a829d8a62babaaee270fe55895810e6eadc350e4723995e0e724f12fb5a19ba88e633d0146b6ef9896dd80c065f1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7cece594f8f3654ac3abe12005fd75e96f6d29e1bb82e43a634aacd64d70c65876c9d447b3bdef0dbc0ee20239d418ee519c1946225507f7a3e9fc8422c66e4fd1fd439b6e1a83f624a0b86e540bc3c0a5536c0695944a1399a28eb04fddeb0a578;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h267cd69701205ccec47c44758d0e02177d950fb54ea39860001d1b49db24df93f9d01b19325f51d66e5a87c3d8bdd75b5c5a5d02c9f7e12620890f053fad0365e8645965b1708d5391fe120d96c0478b89abf23c6927390e59112a1cd2ce7fb4c4ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc91c0ea31939521aafe2a88e8869a43e497979baebdd68d31107089d74a684f62e8110376644623a401c6c1cc214396d96a204b997956a63ff17434b4e456e1445e51d2196c64c44c2db8505b4c73341fb1c6e9659c6bbeff6d08e5b4103501ef38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe1385902fc1a9d585b3e09342f1560cecb25ea0e45dac3f05904c5916bc021d683915629eb06dde18bc59188d766ef1d3885279368ee329c93ee69a68f847e7b73dd2cdf106da0ae65a1a819e9c9de1da4355d68175689d5b156fb433f6ffed3ad9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he33ef383b2c4da6a2f59ad167e3f22e8b2f3a2991dd841b036644ccae574eb30598e47a8e4484ba0e2c98aa5a1b18b1539a4e09f0cec91bdea1a09e2d5d945c16c110cddfbcdd043c6bcbdad68d82b4e2e8216b2efe378f50477d1e9787319af3487;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e93edd31a9ec1031601d9811c3542c91bb994a6117350f1a5acb87bf8e6aa6ffa5982c7684f505468d6bd6a7d4da8d1c10592aeaa311b7e173401c8528a2e4dc81ada353b8cd43ed4875d24a79c772e9e4882583e620c351919494ef14085987c42;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e16ddeed23502482b9b1d30568545568f88fae3922df9627572af8e0fd833161f208686d872bbe57eefae28138ea3f98657b9cf03b190e7bf7e452c07ddcc7e85bb71dc2edc4ac27871c11c966292e9a78aef8d8fbd37ad8ddabed38a3f7c9c3b97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb05e7f2053c986c78fe3dd4c91788f2f34e71b86e6623b3165da76c0cea3fc2df9027249124efbb586daf347df0def19817a85520fd59408a8038eb667f3e4dc29414c8dd055696e04dff746fd124c0264669613b1b6ec765f53433a940d35597a2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72aa405cbaa9df507b843188ba6dc5f81f760e70ad7fb3ba007087fa03b2cd802cc8fe6fcf6219957a41c15923a8e7fe171376551fc32f955ac0a650880286bd7b2a55ae72fa9644bf5edbdfe05eab7106af796742a9baed0ae2ed11969a2c561a3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb53b505b9760c97a929a6e95e7a4d2fa7e2808418e84e4601fedcee87ff629908467056ff3fd965139a23241907abd637a29a686c5d1c3b728e7266db412c4ed9422e186f4971823aafb706be4a0ad09741bba775b219f1edc701752ec0766cbc0e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5e73b222a07d52dd06cb9b5f5f924997cb1dae8c862074fff5c5d94de05401fb4cf3d6da1e145bef9e27e4fa006c433c7bd32cf33ef8ba2bc4f0143ae13368a0092e367e9a7d454f124e04c882eedd51f817c54472e50764531818e022c96f5bc8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8279f172add6375fa98ce090415bfe47cb4a75d326c701c2023c698ea1befcc59a7a45457232710983eef6f88150f58590f1af14885e7e78fd262159dfca0e37e99bd02db1a8e4459bf7d0710cbf8d44fd1c43ab82d57ebcd2e15227e35dcc0f69b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf832d6c46ede468418259374a4239e756f981bfc4568b062dbaef7e63873e4ee911908b27150525e9b258369b3a1fbdececd3496cd6b7eea08f7b95ddd522823534f8fead22974e481f7c7eaf37c2e862a28d71e723d644f1ef85670045b855e9bb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b131ee51b2ca0375f7d0a04b7fdc8243c255654ac259e438a03034d0a643cc049966262a10d75f003e0d93176670a6888ca5b367c3d393e59d6b65b9be91a1da53fd7b898cf92fa105e8d4d7a263c22780fab71e23d48d68d844c98b211dd023ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7548e3286cfab744cc113843fb44db351aa11f1f345163a980daa68db0b13b913f16f8cf7bb56f64b313ff945fbabffe20f4a8d2ecba16c4cd30676a19293d82f790ffe3acdc716aeade5d4461fafdf9f3089d5c5b2d76900996425e7a9bd1d7ed92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a73b8337c73d6d675c74ee63c63068f2d1bf15700904ab226bf34c94a4a9aad139f1931e6455ac4f8bc9f1761987fb7c086454849eba4b3decea7e8e2f0d487bec6da2931ddc9ed7a646fbd53ebef6209eb2b8b8e12b1ad2ac8a1a06d346163bec6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5b6640345af1fdb445812eff137a9402a9aa6d128190037a5d5eaea6c6e24d577cb6897aa4ca93203ace749c2826030bb2adc730aa012e70ac83e826cd0222d609a4c179da45743444446e992acf94d20b53bf4157aceb0b57d20d45c0a7eb4406b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bfd9ab4c5f4a9407461f22aef3e56fd1cc172e87478b3cb5d80473222b8850a3ff7e62fb1459836aba482ad42e19f2c96003b306794a87f586dac678fb20244fddaa52657de335adb7c48bf1da607fce4e9d81a4650e79588cb5001fcfecc7acaa9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90df6acd66d82a509fd759c38e4cd69beffd6fd81bcd73781dd7028960a34d9a27db91b7b86ce5a5cf82a7bd57fed322187f67e470d44c5f51becc0aa0f3b529a5628d4c727cfbff57958b834c68860fa1170762a058cf4fd1ad94919f953417bbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12caacc5c8fe30a639f76e242bd09248b6b22f38bd6f2ca63d19ef3345d2518583c80e92f470cdb640508932dda79d0228eaf75d284032798128563ccb47d540ef06d1893407b3daf18a28e397100d777227cf74ff364290098547a144abeec75c97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27ca09021cddb68fe31944ceef5fce56fcbe6a1afb005437bc6e099ffc061f8ea2a72daee96501f9b5373f8e0608ea1c671fa329b6b7d51c8b6d68fdcd47c3ba6e7dec5763c108d3e41f965f5828f77b25927d972412d6ca084c106cca27e3ced7c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h243a3704ed823e94daf644798fb2b662fc67669252742e264f1290d17ff0465df12be129b1943b06efb8e63aadb60a4f08234cef7fdb5fb235b361a455d6ff4d815383c3d4fbae5abcd2100bb088d34ea0ddc729762fc9b5930b9f70d6d5027e6521;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h109bf71fcd6d4be637df694e0773d896acad40067eea3712867a6db01e9166a025df60b8587745c037ca2eb7585004195a631ad55a0cc3c99fa6ee43f6c8702bdbad580ece78ac224261517b6abbe64cc40c8d5717f96e3d2630d33f4169c3092c3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b043e4ff44b79b0b30a2a95c8cbea899189bf7764ea2cce96f3014350eafc9f11fc5234a963bb70e958a913a812845d6029d49123b6624094da8c66d38afe63c42fc139a0a0afc76742dc5608bcdc1bee4b690bf6d27871dbfa0213cb91e1bb2837;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha27c1ea049e53a55d663b5ba4fecbb4e1ed9c6e1e62c243372b775fd5ba43fde9f0fc547f81c241293e1da7b5920c68d3e10affcbf6dd46812e65cef1ac4079e19a2db0a9f99a126ea0a4501fbef0e904f978580119abfbc1a23892ce20d96ccd010;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafe91f5b25850da12cb94106f170604bbfe68109f75ed5ffe37d09473b620c30aa2e54af234b6a8906c831c02e7bc18cd72f102b5655448fbb272c8099e6e4f9dd2e29407ccf8e78662ba9c161e867876475e0f63d1b3e69b9bf7bafeb17d5d81371;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca075fb89d043bdb0947e486f7906be09b0f8ef6685e3ac22cc376b6e305d670dc462f9674eddf57e1d542a646525a793a5df1758aaed057ac3078c6503db3054d118ca14d3adbdd320ce1340a70e2fa4794927041afd2a7a792de98dded754dbea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31ba0e8f46f2d2073cae951cd8f297e0d52ade3eb98abcf7039f725d2d7b7c647659dfc67dfc0884b646277dd18f52411d6d4349aa68212ca118fcf8d1989f744bcb8db502dd62ed10b964bd59ef10a139178d688aea928e9878f2cf82da6e82e954;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bab20f0e271937e35d065865192d9b0bd326bb365f236ae6ba36e5572ce4fa52002210006fd113a6e1b915bbbaccbb62c15395b13a822917d0fdda6add5375200bd92bd93ba7f03a227b8904f53ce01547d9f72b4a6b282cbe5396195c4dcb691a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24eb91f910df2949135eb3131b1bf560e695c19434eb103be009cbea6849b5612f710eb23837557ecb907f90caa9fac78e33c7d82898721a3e9e3a4f29b68689cecbffd4a2ecb15001e37b826572b9195e40aafdae1431bcf4666e14c2237c88b1dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50e5648b25c31ac48d437fa289cafc1bad4d0fe7f306a72f036f7f4759be73086da79594602e22ded09e04db90a98eb6875ef776730581afaf5be990b3236d288f31b487e28ba08f2d6abe563c4de092596e167eb592fba9fe90744c3cb0b7f15db5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8f7463da4d15f6f1bc53b27ee88319c5d31040977b3aff32e3a9eb5d52c08f78dcf27fa5a56e284ab1f0189b2a3e516f903dc1174a8d79322f34dae5a3a7e9b1ab444574d4416ab66e9d028fea01285900a1284b273fe71123f6d2cb2ab40f8a37a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34f45418e76c810c19f9a85758ddba7560312de525535832d250a7ef3328842b95b70dff23df10466858b7ef6fa0e8c1fd8c2c102ecef4ba8033e2ddbb20e3aa90ab9d53590ae2b521ca0a6b9bf14c9c40ebf121ac86eecf87321af4b7f7db5b04ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he677d62d46c44b6676321090e009edaf99339b681f0553f8bb7aa5b26341b3bc2ee1724c61c677c80ca4d4948d72cd0f2bfc580561cbb2712764aaab91e82c18609137eb1e7eaefcb8255f02ffa42e73cce2b8fc20ca58693758c96f3cddf1960ac8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he468bef83ae837f36ad87d34d713a11206f2d187a5ab230a9c5f15b911663f156ee4656754dd5e32060df2b16b4ab6838ec769082d2058ccfc4ccf782fb192482e6ed14cc198fb730a870b6773a907b2016033bcd4ea57ba98ef4d99258c0edf95a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha39b64f2b58447fc26c7e020749e1b0be3765cec170c6f42472803e772bb1f5c91622183c7ad89d3bea52102b301b97bc22b8bec007b9320f99ba753d5de7a46f0aa2cf5db6154e2ea03025642245c2d498e5b918a5fa456f14b4d3e8575bb260c67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5f6bec7322971aef816007832cd6161423fa543609ccf92e03b4bf6b9b2f730364c2ab318cbc2f7a6f03477e48b4c7434cbe3eb8cf72a5c825bb7c2b3b1e443794c3d6e85fdd9ba59423af81356138bec5877f953c4cab5713066334b918eaeb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbc1fdd61f8595531f4b9be0575bb59974d14a24e1bb4ec6d0906782c1a3cb1ebd20b3e8d908c9c40c92822fc415b688275c3f8bcfef2ca12098fb93cb5b99fcb8767b726e3e4bada48c82f01e58ef4397eca6b7a07f1c7a3bfb38d75343d06187a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94f5a1956c909363815bb12ab319dc51378a2d4061207ffb2cc2589df272163b348909b1e91ebfcbcc1c0e97541c4cdf21a28370dcc1544647bef25bb2cd3d3352bf8afaea7a50bcc8b1bcdb7ffb293f99f006b4801332b87d65bd211ec1a6c35ca9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h114b67cff7cbe39899a1524ee5912c37f4484033952d4455a4d93b166703f4eb8e5e17cf981b6fcc0b34192e0b27d2755a20e48c11e40cd4bc15ba282a8f2d8c5e883ef0e88f1d8387f61ac80b77c1d95480d5cb3d37f29d17befa945479a23f4b6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33dc2638e9ef4238def19fa5cbd854dd03934f8856fd60303b2b8a8ea9205206cc0a6499329d12a75f37a52b35aa8f4944c6ed4bb3e2014c9dd26c41d5f7e06e9b03876081bc9965440e7d05e4958eb84a64b91cf2e6915f394b30bcf2aa8c4b39fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedea76106a6a969079f7cafe069c2c6b89667601c019ada5e4b256d6f6bf8baa0da3f2534e62256e636444d7a567d9559fd6cec01e1a80b708777c0ba36f6d082e5279e1c2a2476d3216c4fe02fc182431dbd5c8171d11bb49b0e29707c49b0768a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0ad70eecaedf996697628e4cfbdde769bb42deb18ccef8a0c9d1e872b461de41c650441c64abe5a87953f4ec4914888939078340c31083081b506666a36f1bdfa52d853641681f379e937509d80ed8017b2658ae4d1409df86ff145b18f7af20f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf482682676864df2480fcc5cb5cad84e97e5121e0d8d043d6a0011c8ac3f5c9b97daa25c6ef5f6a9aa19fc868c1259c91311989e32b22ba8017a91f3566c885c366310ecedea4f6192d1ad54af66f953827c5f634fe06f2e812367d35f78312975f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37da35ce33a0edeb8f7ddd419e6d9b685c18a45e175935afd52441d535d7190fcc69a25f9ed22b019ce719dd11db9b1e06e7179fd9a52c1dce23d097cc0820d17f0a8ecde529803eb99e4163236e50581e15965ca520ab322491b2dd390199c89966;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c928eb65acb4490e64c3870cc64a4fa51745372b335304083d299e34d1e47a707a4292d26be9fd5e01c25acade8bfb8ee69845eebbd1b37abe72757bbd12d029eda3e7ef888b2bfc7ad6188efa2875a51d4eab3093966eac3daa1dbe1fde06120a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a792ae4f28a571d96bcaa1618d89ce814ad4bf1e96ad1fcb2af755d0a1f230865e8783f6912b373b537bb2609574d63b743975103f287693306965c7eb44dcab5ec47140ecc44c4cd1749ac23f692fea287e91c0954b4d3cc8894748f56624ab16d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64131284c3573c1e7a5eb7d639d10de99789b83e085deae07f68cd873c2ccad9468efcd48050065e0473f928b47cd49eb6d57fce040801a340ca6419eefb40f0bd80277cd584fcbf2645a02f98f19e0c90262576f7aaf17a2e93545c665973edd0fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e5d885f84c176398c9416ec0cdc2376440089e45b6b3816f0a1e920931e38ceb2029736692a5509b56efbc86dda64f5b4769541bca7fb684235af3f89d1c60076a7f82c6a0b912930727c35f4f1690b91714cfce87981c4d32ae8065a5e82254ba7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4dd741853f87df3bc6904cd43ebebfbf8ff68691ee24ced91f2041a151b199ddae90ee70151ba1ade475fcd1e7150286e50b48f1a7022a25e229acb29f0aa3295e7e66f00cc27ad683808cdaefcfce87472c7d63e7228896ce9b8ddfcee55556c639;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb275fd9bc30f6045e31a834c9dfbdb94046d2eb06021d65c6a5908b70268fdb7123e0ef9da9446e05776eedfa958afe6fb3c32fb841fdce11db4b327a8417d99a83be3295e72a5b9f6c531511d5df6790d38ee9e1ae545b2f5820b90991e77ac6df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h334d0d3bc9a6319235afb66bd4a12236e61989dd94d468c28c7849415d7b9034fa6a511ff77f69d1af1c51ded67c5ae03f0a145640b8f63168b32331bf0665a9ba8445e42b36dc7baa76f01da0ec59bc0f803ff89a3089ee3ff32e37f8ac4797e523;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d96adc7a739ef1a83b4619e9e00e8220d8af43f0639ea1c9b651a3ef7c2474ed210d64e3a4275738be83ed45575a43c74deffeef70b805e8a644f3cc85286bd5e4c44d5d9712a81af49b47f0bc2b3753b9419c0c20b31087d15a3838a4be0c08f97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h853c15124c3c8c70a4d7e84cc37052f51ad428286ba6ef4fb0f61a95209e926f078bd50bf1391e9a3b7f38a5074397e95e4cd5f94e59f7297cb34772ca14fb042dacea84696e64a11792647285db274a83957f0fef78e09cc3237ad343c0b568729c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c2fdbf7cfa564e42fc9eaa509104011e9f6d52e707d3dbda5b0d6244b04d198aa57b7a4903c66d0d5a0b7f0eb4370879ab8f91c10513f5eee6b12fd1b1d6cd75371c198ba35ff7ab0a3d2b45317d52200127ab9f1045df28535c9a1625661221b0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h355cdbc666fffe14d01fd1d4897f82c64d3a21412becf6753b52d2fbd9212ae562369e4c1fc9390a1f2c50c8bbfdd95754f00de6566525aeb2956c460ab6bf44192bc1f579c0981e1cbe6cd2493781e8e033cedcc1c4867625d3b3671ac700d7999d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6563e30e912462d0d1e4b5ad21d13a10855c0d4e8f816cb6ba721d54eb389161a5a8c011f69d47eefa15ea5fa3dfaf8d48efeda8b57255130a9d11a911b40bdc142cc09de27e05430e1f9a30c33e1bdcb8ca440998fffa299988ea2eda021d8fc998;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8dfb8c30fc49d0d0583c1e77f3f90b0e13a4c49baa2d879d0688360ec535dd532dcca4893f5ba8a5f5034c9265b6f960ad9c2b00dcab52ec361070d5995ecd5b810c497dfb0bfa85067c7a9337122d9e8ffa14e3ba0e376ac784793ec1742f53376b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f23dff96054f9b2e759928b72498b2831effda04cd578160c24a47ed61c6c2bf435fa08f1ada9e82129c7f84e31c29104cc77228279269f4739396bc3d5447bbed6819381ded2c24d3b64da649da23884b62ed50a277fc936fb0a59547a36ba48d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafda718d4de29dad2185aa165d6919c82cfaaa367eadae4ad83a8eb2d2fd3d2fe0f938a95189cf2c3d3a19d47bdc95b813ed927b3ed81f6baf3543e6df3ce446b18ccbb18ae028ac0cfcd24d16e7bfb02328e5da6780ede8e311489abf525a8e478c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c81a4865d57315ead89cacf5dfdebf0430b690febea0150c5a1998232f514f976f8ddc3c8a5d1eab979eceec17f6766983d1f247f38a10d77b16358c08efccc36b58f049c57e8a869eb30881283b2dfe4529688e7afee2c29ad82f232f8de91b3b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4495c73a697ce9fd5248a4b3ec7b6e0d91415b49537724e15299f6e87de9e98a7d5e79a065c52311cd70b2119362820342684825b77386db6460601ac08037d910f8f7a8bb66aa3e75dc23dad0850be680ab6c7aa5fed3a40418cc1a9bcebb79daeb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e2c01f531742669088ed62a40f25ff59dbdb90eb0f030af37b686c3b009bc2996a2077683e37dc55106915be4beedda2f1bb100b832984f5b55a8f7813f619dfceaa023522d4eb0d422624125d0c2210c4561c5bd7606a186118afe6d836e82e998;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc89ef5344962f5b15c9a6a565ef266f40cd982258b188abb0bddb6f7d9d243873124984a1228798c2ff173dbc7fb77218d478d48c4cce470971e36fa4d17eb0c9e22fa146d44a6ea068da3078ab0cf9620dba8cb1154299231939576599d2e08e503;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf817a109b0aa1418a6a0aa32e91378268c9d5922580fcf160d16bf86a027303f791062561d7ee2695c42844a99a3a21382d4addf928d86cd609118a93a2ec9a7ecd831af5717383628ac613bae3ca6e55f70fcd8178880340e515814bb2a3979757f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50c1309cbe053caa7859a8623e0d09231267f88cfb0c40930f734465eaa36e307133e468d49a45fc99e65a66f0d48b515a7cc84050b005226f976525450ff9d6d0a8d89dccd65fd55b10d29cc5a7e5390ab58892637723eff22b4ee559944f77ca77;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74fade4667c4a804e2373811f560432838b53de617661eeb818e810eab71e14d4fcee0fccad288be43b771ce297379380c583c1a8b05dfdbfd865b5fc4761b140ecf36090e6670e9f4194912258d6bdc9e903b18e8deec800fafb29a537611a3ad43;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fede92989d03f9479a7c416d2b7d69b0de49755d844e4b82e0e34bee690b3511703fd2d8e63a920f113074d5ea5db4a2a037702ff1518faf500e0007cbd5f1c3b25bb0ceff066bbd4a2a3cb8f61c856ddaf5b8dfa59bfc32af8a6c1e100e603741c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc698cc1c2fc84e3a81b7f4cc8cd96c3433fd19fa0ad2e8db336985b085b9891a7561fd6b381883770c0e2facef701e3756d5a65be69826eb398f6f4e20a0d6154e4c443893006596c80f3c36f2d52edd58a46e17ca5b443c8ba0dfc26bd6aa6834f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66e2993456d84ad5d87ee57214f3e8ab4ac38b504ed19679af2c20ebc7aa6959831b93041b2dfb08dd3389f972868205802f94f50fef2b62ff840c6b654894aba4788ff4e45fd09546d019f64f612edce7cc8a5131ca899cccafd8a326b03a24c6d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3de797bcf4dfad63d241aef32ed01636fca30014b81b6ed87281eba1dfdaa5f45e646c5867da1ebf45b08fc8ada302374acad55ceb9790b2979ae35197d28869f0c1766539d878ec9e9af6e9ad20f3cc8aad966a1c628471ddc08ddbe8620cd2cb72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2af480fe118e757fe25f8a2eec629b33d1be2c82e2b9b7c2dfb61b2595574269eeb1a0e0bbfe0d39dbcb77d766462e7e11d52bfc2f8b03f27d6940b4089339c25984214057b2baffe3aed81db54168c4999e5053f1975c722c45838a6adeddd7bc74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc85fb793ae4a48e31b415a5b4fabe25a0f8584aea30b7126dfc1f57ab7d9b859fe2d27b1db015e6f7cd9cea7f99f231fa25f16798aeab4c3bd4a00887885a014e5b075f86d4fb8821a5cf1e7928758ab95d6d30b306429d6fcc61c99dbab44438a8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21e3262001006f80763d942f91310f1c8b0bd1c7960b45bcd7c7647cf84d9aac4d87ea0de7359b95943ae10aabdf25b9ed1d1ee9a5ffb4521161cea81ce9c31b9694c1e5b985b4e8ad0ca5e187cad185bed823132e72802baad8279e418e9041ad8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b62c52703403227a32eb5843cf84bfa411ecdcd86e3bc8b7a867fbb6f5dc01b934dcbda7d7b3cd0a2810a0f571662714ecac02541a6f70af7c80d07de112384f1b566de5401ea9893002996e7469f2f782731667b805c0054ee16dab7b0ac80e4f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4eff250ef2c2be10ea298fc042412cb6648e170cbe54f33a2c1cc6a73c3de47f61b07f5f5760537143d56421f3862e63dfb83fb919d659a1f8096c97c9d99809ea559d51d516668896418dd22a994530c86e56c17b0fb688c780243509fe4e758c12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haee2818157947ef8cc947369a3ca7f5665af77d08d5df96f7c881fb626dd3cd2a6b8fdf470b0d1b5fbd9421107bee636847d7558bddc3dc2a5a9638f2697d0bb4d20654183bbe3da6383fab135a14ba291a234b70ee038defc5aa4ffce3de532a388;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22b2046de0b158404f5beeb11536d4ed0225550723e54fcdd6634bc03ee8d9241949bdb95714efcc0fca4acfb2ecc0f81552e6461f760e8c37c30365281579a7400e933a1ff645148d27d551543989a70a9757c1eadf411943553282f450589ff730;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd46fd72b6fa1b3e09d5b2f2bc46538a4a691836812f266664dedef93efe1516a69913f95d43ecca77de6a40778e8adaa402c4244392ea860890d455deb1b48f3ed25233fb4dc652f14c3a67b13bd5c654118d2fd75e65cdfe43cc4cac65f54496cb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9c165b020303e1cdf0496a3a3350f02e6b71efd553c5792ed7f4d6b99e6218c63fabb4592de1863ba97c708410c8239e357754f5bd379c5feb86bc29c12ec134e0075ac6666e78174eb62737d721df749650f5162a9a0e2280350f74d3d3579421b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33447cf3d58fc62aceaf0e902fbbb0c3f44e3f84e01bc64b3f087e3c23bb28cc11984e323d7eb8ae9597860c46b0269a5b2eb324e4571f23e1996913c60b06d90b33dd85999890394d97b00e9c69b057f92e75f820e17f5006f6b7a3a80e8c743b9c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cd6667f481281d9dfec6fbbe0fa1d3bda4d98dcbd889b616932199104f0a363db2cabcde016abffbabc331c19429f12b099d77fcc2470b58a55957705a3335705be1c6e778112728d246d1a616a3e2cb2e9dc705e52ef7835a17fd5213908b71804;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8426e0901eabf3f4ae708b6d72ffa0e59e98ee0085a8641b09249e4af78c8d49a53d8bde44870567cb79d3b4cdd0d909fc29c326ee41278d8aa36e1bdd2105df82ed9b341ab711545a15fe447d84db3e0d3c861c831ddf5e629591b17496c08bff4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1aa1267530b990edd99cf6f04d15c44bed9940bad3368c7dbc2067a09d14bb3978e0fcaef31ced7fa79a042bcd8c7bb132da1e714da1a1a0799fb1ea52b6cea4b1d36598439f30f50e6a1e4265582ffe626511dd595e0b77143dddcf2310ee8a838;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h603db7b4004395db3070aa4c132a0707b5c38d6fe4b687e8264ed533b6e4cfca2544ae9f2e2e2d218eeb74dc0a6cb0eeb3a6f2bc9725be5e2b03448fad217fd8667b3b702fb778cb895033e9ad27b52e14abd22060eef38d701a517a147618641b27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71ae9ba94862733edf9ccbb55d3d26d555c46d8ec04d695df042fdb7fab28e630eab1cfdbbf6307b3f69616aab0955ff3b8e5f005a2dc38298cd40bc14e4b1781c28803332110d556d117b4cf18f48232225c5ec5bc51f496ce72b4fa32c151fe968;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cbba0c05e1db226a019f3d18a015f29bfe51bea33c47081a15bd84ece4aaacde2213f492845f4df133aaaaa2a5c7d718cedff32a6ba955d392c86f308bc771775ade60fb20f5ee4c0302942f74d735a1b42568e0d483cbbeac367de23e6f095ec4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb27500088a164d5399b4c71889e4e5c263804e092ff33c6a82e0fb57a73d10b9d6e8215e8d50fdec1bbe226728c52cf9f76bd5273a5ad67598647ade8812f6026d12e3352d368e6f4ee6fff0f988642ed4dc49f10a706d1bb13df574aa4210df39c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h981829a975ca2c4a2fb055682cd6dd3a2c9bed7932533b1b3a909c9637e3801bb72bd78b0e2626c3acb1e629c90ac9055ed990f1e73232fae10abae39e8bb4e7337ceb8b610a7898bb36ffb161aa68a15e55b94bebd9bc7ea846a9852b70969902a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63bb82e4030023f32fb1aed91a5dda2187fd7ddf88f69aad30d2f5d576656ce75e9f485ba45e028d055a7ed1c6e5d7f55d2414915e24e610d0c746735d44a7b036fbb7b3e2ab493e3ac407fae49c2068133d819542cd7f69bfc3e29a2516818701d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5be3648836f04ad93cc7d6da92e505a92f78f805552d794fcd68136f53f28ab8c52ca4494a073ba6c28c36fd5d30f59a7e8d63ef6489bb66a230218d9acf061424f73bcef4de217d9cfab11b02bd5988f24eca98b455caf81c9e3bb03f586ce7467c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a6e8c1d7d31a80c1d88d2543daaf186e0b4d05d70f5e246b34420b278770e734d18a2a9b377444f94bc62297f55aff15f6de86b57187f4437a654865c08c3ed25987687a17dcad8ac0e8d68a5a9e2d287f4a5dd0e7c1536576245c349b677f66b75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16a9f2d14a45a07331a3dfe24cb9d5e4401a5502cdf635f366c336de66ac6c57a953017b91d00b88dd0a3b51ff42faf2dab5415cb3b2b71f9f6b7676221238b4cf7bdad7b4b5fad7810e6b58ce58049780974a539ff666cff9189ac7d43c6a08d17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h538783048e2350b2a51aeb47408f6b70a8d186aa6bfb879d7974b899ed0b5692a16cefa0b7be65c3d7a00fb574e58caf612a857052268712d0c030ee14ab4b4cee25c59dfae7c205785ec1c40f849864b97b05b03ca85bca6b70557e9c6e70e6734a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd408d4a1a9f08c4d3088c8855c6ba9c6dc807c5e2cd2b0c11b58700c91e748bbbd555e011ea055fd862bcb67f597c39fc2c5c35f556b17bf8e87d8ff6cb28d199d5e708ba5100974faad43e3fb1194bb402b25646732b33e14f81f9a4e531bb20595;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf5f9a34dcf6bd8da1ff9414b4de401e3f64c46419076f8d6cfad4e59870798d3352aaafac479b1fbe2a4f735b5ca583113c71b9f0158f47c2df7d9106ed76cce2c1940b626617fabc40b07cfc5e51ec46d14205b465e3f022a358b5f6bbbc65b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h614e3e7d2ed45bd7baa2ec5cf33a1cec7a938e3f5f498fe682855c8e706fdc7767c1a48aeca0f52da5c0379a1ba8caa34bc27516bc890887bf30157ab8c55c851484842930afa447e4efa47b003f94390c72d5ba96a699165d6aef30031506e9363d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc76c18988a5f74b8a0c98766c36c9ba6a4bf72e89021a5365dcfb86a9bca7f7bbfb77497ca0a67026b7370168b208a5ed1ab46c1bfaf6c0ab9be72f38d0a0e5a24eead0991025ddb2c3fdcbbd5118f9933df280797ea005dc5ac16df90ae731e3826;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he842b7bbe2ac602e0eeb6bf76801259f9ac11f870d7f6c75ec077da7b4639e817265e7bb5c54529a95aa089b3a2beda5c23f5db0fcf0dd4b0ea0ca3df78a9c33f2637c21d7e680537ac7f8bc931e3db368b3692c1d08bc80d3dc9356eea5bf3583e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca339efb987b6bad44f6f4c2105527a59f927a33c19b22e6d82e62e741075fa44f86e7145189eed492aee09f9b09e63053deba37418e753be1dd08fc59ca30e4e7faa6370bfe97c1f5dcebd0d0f0618d695ede311abc2cc5d35699d241c4405daa8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82f0ad30eb868afc92f3bb976b810803c2d00c0974d88f687861b7419f4a77eeb5b682c40da3b2914cf5a9ba204b46378faf90a8588435ee82ee4f6ffbd75c66fa4dfe60c06c2a89c22473781556455598dd2143898264342e5c457060aa69f366ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72d43ff352628be9f2ea2418cfb59c92f1bcb3fb5be480a3c25d521cb292d165b012235ab666360bd7933cccbe406b24912cb20591610aad4eacf301afe7a95b7ecee4c845d20fb0cbd9a1a3485aaf23b39dfc51cba849a153770a1b86a9e38cc36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52eb287ffe352c473415014c4c11e8fb0c7faab1b4e0346e81bc823146462a0e84c4f40f7553914fae5a6f0ca61f78c49b84ccb790c309e0302e89aa1ee41d5266f90500242500553d63d376c6573149ad443a4e9e569044f43bd51b79468c925a0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f91612db50c129e2edca26276db04209259cfd8e10e84f530d87463e810888d37340d2031562f74d56aaf8d3120dd498ab35d253d03c783d90495f53f2928d549c71ea9d84a1edd9b6a74403e20693fed3ce73d1efddb58b96da79104b930626596;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf89e9b332a57422ecdf5f6154d36fb421c78a7550ae946b1755c307a2a588b723802d22e152b63457cf2f5fc8b5d2f2c1b8996795c3f65c62d507b38515d76b221d63e463868c0dd10322a19803bd839a8588b763041f57739a6deb24f80baa755cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1429e0034d3f7cd50f8ebaf8a6bad4014383f5943482ee1706c4bfce4208c1752804ad3ec8ca71014b6608bf779a81d7b36b92cc881361cc02ecc6c2561438eb8d9e69696c678cd8e3b45409905caf48ce196ba0447a6caf415ed17a8bd9676021b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7fe9ce9d738606d0c0389181bc8d8397ab5ddd9cc184df5f8b52e0dea441ca56c16dcb33a94b80f178454fab4f69c04b17d6927a4a039a7d65f7c7d26c64ccdddf02da32a955aef695cb81aa5afd5a1d13971ea5434708eb846c09080c4f52f2762;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed09e5401b7faf7b67523a328c8611d10d64fb3b06985eef12c3786c00c3efac596b024972236d35d0c9c016964c60e7a2cfd6ee77e398920bfbf91efe4258b66f113efdf7de137496b610a8555999fdb68d3aa46b7160acfe92c99399902a1ed010;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38505e6d1b1ac3416252a8c6ce251a17519254e022b3465202c1eb21b075f037632e64edc9a88a519169041a8c20b12edcfbd85279e13c733153666157ec27a999b3fd4db65a0df60c404cfada0b437d7fcd36eeaec2fb4b901946c377e3abb3c17e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d22022800a0c22c8ada4c0988897faf104b5c9177c8a20022e42f006cc1bdcaf7690934c40b311297705201d60a5b3d1cc4b5c727e6b6d12e3cbedf61daa8c162a0d1be036703ab9f5ecac46c6d5cab4ee4e49e4bb52d8ad1554524e97b870c943;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4acde6f7d860552a356c628d2e4156fc4a7766399413daff9220960751af8e78d292e371affb2fffde184b3297edddd37f074c3235d4172f479f109439f180950c35083b48003105d82c7d90998b89033c1c3f88f90f8cba522753fd25818d72757;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had419615adbf9bc25d5dd3ee453d923246db38e56501f13e32aa5710a836e055fc51c42831d8f9c7e77df52b4814a20fece138a25b306fa5c54926c8cdacb405fdb9fc9b051d0f72b48a9bd9d116c2db9d233e58ca5d1cbc1a1996d0735bc9c2d26a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78cfcfe05b4c7c57fa2506abaa7927bbf8f296c1d53a81300c9cfd345ed1f9091a997eb35929332da4b04d4a4c0589950f761354055a7374abcfef4f5ffec0e922336db685d52eda353d93a8c35df02ac28942ba5e4d385db2b6b67ef1110961955f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2d9f7b7bb450eb3b238f4e48c60708e259023b077d463e609cef8f07534eee2ee8f477b2918b65880e7a0430e17459271c4c3ae497ae63a8a354aa69810f8dd0a262e388800083b2f28f00ffccb4b5af4a35bd3ff3d9a64c0a6bee835f704b48995;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfe572fc74a5a0b06357d9aad8fe5ef6853731424a10d047f1749bdf3c014e0dab9263df9064b4d45978078606f01e7e881e7786f5ada963e838faa41345b502989c77d51f130a5f8ca84cf801460eb3db59f7c1da9230e59daeb8239811b7f6dd41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa6f028ea37666a1e7a378e6a5a63e70fb13d0640a70548cef2a90d666ea27cfa936ec9ff5d7488f13b0c460b1f19ce9486b1bb6a84c76e1d6f92464e798d9feec5dc7e9158012cd91c8969e87bf65304fcc0a02dbde5c7418a0e8659dc8caa29c36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h821ffdb6811eaa8e49b9e6864e90866111852f9abea710cb3b3517b544a8e611755995f8537d813bc8a327e2bebdf222305850ff72ccaf31f0aa4647e0d8eaafc8ebf3ea23043d053119461de56267a2b4e630f581522bafd17538c89cd8a4360b01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2122fe41de89248f6356a52c7d6dd9540f045cb0da9a9fc7170f624df3b9e42df467d1de1333a88fbee4db3f83fad07941926aa4d63c4c67506f238b04bde613dc1cab01db70c1e0a2521c68b2c27d95364a0662c4a4f0a97e493acd41a6ac41d54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60c8b931f613271c3b99942ce1da83ec09365b214ec85051a3d2e08959bfe12269083d732e009ecd322de28b5facb63ab931a43ea22b9999538f4227f93deb13629fb1ef60827138bf73e9068c5939373aaf6aaafab3ef507a4000af86ff48d8533b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3af8101d96c2068d7c900fe24b68fdee52b6ac96f2b3028162a535ffe5320cd0c44a6095cb651ce0c23b5b233e482dd35c83a4a2c8671f43a6db0e3de9bdfb581a9faa211be9151421784cc01e42076ddbed73215d9af462c13e02e223fe4648520;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9247c1d5a7e763073ad990fa33676456783cdba81badb877593b9cb0169219586984bcf71484b3273ddb147dd82b2bbea6ca3a048245c0f571cc4c732953d1d1b18610964e13ad3fad90c2f41a1d88d58516c262b4b03d408b72f7ea975cbb6aae99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ecd83ed94da23bfab42b8ab8cde71af3f08b99f8fc0dbfbc8a6b057a1f24cee62b78dd98a9d38106846d0ee28f1406be5de3e9e98820c5cec6b9c743a46dfef1cf6fb576050099c10216d0386dc8d0ba828127150def0c90c587dd9de0528488119;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79931ed433abc2512cb002c3d9fd3b246e867d4e4a09ac5b1b1d591ca441e5539190cecc9ac2ab01b4a9b7cbac1a6632d3ca03193d3e3a670e8832573d0f1d15bce210e1d1563d4d4556cedfbb62bcc218a43429fec3fc62cb296c7924517e8a4024;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e710aa195ee8aeec2b6545f5bcb3caa7b602a0a1ea6038d049cf43d984810c6fa8cdae3a47a54130ff6ff0857453598bee019f60b6087185b042c5ec745aa3f77503b82705e36ddd9a2ccf22586789d8837f49e675b71408dcc64a415fb405eb7e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfd1b9fb7efef018eabf016336fbc1c075766b442a46bb763b57872e7713e0208d6b7b879ba2219aa447c1ad165284fe1951131f1fbffbbab721d1f59be3ad3900318f5423e49c25f9bd9fbc7310d9719c08cc66ef649f2fba032577cd795d3bc1a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ef323a5221a28c94183f97ab21d5380baf29817dbf8b0eea8a390101b585fe32a5a75c23922f71d6eb8ec194e3d91e29cdd93310db635a38d574862b9fd1dd0090195dd9a4cd3aee866ac5bd4cdbedb5c7c90442c717840d009a7084b619925d940;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a7a75b33471a090ae670f726f7aa2f9a8e529a82613b54b3bc760fdb2ef4fb5b4cda82dee678d9f5a4dafa64e6df825f4fa757abd49eff132c8c0b00ebaead9daa8315df7492b619eea838d883f7114cd2d7fed95069b4cc634bcbab9630fa517e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d95838a2b13b2f322cf696309a535f50f45c22212a58b7ca8e90bf71f2296e02b065a7f9f1600bc08b25b140e99698479b86e16319e5a1770aaf9cc3c3f3e324466a5cef82ac4bc464b34732f34d00345f8fc2bfaeb34f6973a4f82cd40af120a00;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cb17fcc93710d16472e956b128d37d65ddef3debe4e33ca2d9341c53b20a29bd9bdcb9b2d4919250146df32cffd8a14f8af3361778036f5f6f31e9ea0a69fe636bc409a2fa05a5045313efc6d90a718b8f963c9622cecd3ffe8a06b5309ba7f030;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf41313ead91678405243d52a20b21def0a29f85e34ef86c0269e30b3805e01c3cd2b219684733459c9adc4ff7d0ce91b5b43ff533e12b02a31a2d3242aa4526f43cd330fd9776873b3b2b6e851d34a4e1d22702fc254e07d4778d86a4e17f77733f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1efe9af8c7f3c4b053e3d2ee6de1485e7057fad7beb075cefcc5ee58d7126fdae6649009f43885d99664166b79f6a986b24283215d155d5413487b40d2208ebaf445c3d8c0861bf5bc6c37ec64ba7649d9803b79f8a7eb9bafe648ad3e721c542ae9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9375b8f80c8a47e013414dfd65f978393f2b56ef71546fc2a9b63b8b69f3e7e6cfaad4e701622858b2f28ac76b9a9b7218263b5005fb95b7816e19c339fd942924aaa7d56bb1b064605ca9e44c7a83c7dc6af511ff0dd05a68f0a7320993b6e21342;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bd39a3bc5bd590f1810eb92d20f3f5702f11aaa53da65acc37bf4931fc98f49938abef36f63a4217afa05d1d6de03a591b2cbb188546e47f191d07c07ba8a1bf1aa45a4cf0cdc5507b767bdba7016c4cebda06a279019ce597dd6fd37bb16fbdae6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c1d414bf3dd37ee94bad935c92129697f966560b568ab73a6d5cb703246402cb604c8fa03090eda4c0d0acda36605fac37d45fb1eee1468fdbf428e6e4c68807dbc13e62dc4d317ba46c901262f5a2ee26c58e28b03b1fd363b77c9d4f1f42dc20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f9559aad18e3184dc3f576f85000d16552d79a4d53c0a46e56f761a9282455dbf5a230f32da7aef0da0dcfacf1905d5ad24594ce8f44e6da9c732f46f8eaa958eeaac3925ceca31135b6301d4407c3eaf22fdef60ab081dc32a2b9a62c0d226ecde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27828eef59831b99f616c36c9e1f655a339041bf6832c20b7ad192ecad4cd4f091c6289f62827f66043c6be8a2420f619bd571a6be7b1b25f0c130addac6a8361037138bdc8486fc49a61b143922c2f79208cd5c11ee4ab67d2e5fccbb36844d0cd6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8b57620f194c7635762081b8f2c533df328467b5b0df70078b32a8887c25c0352747814b08a137e5accc2c87e56cfecc3dbe03372ce145f97ddf44ed18703cafb7f0520ac15161f66240c474f68fe3a5ce1c6acb75c3d3c2f5a0a94784b94c11a65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h167fb87dd09a1ce5407ea83f55f2ffc1a51b5bcc3d6ce02a1414023584b7a1667d85293b5a41a587000ac6a49b6a6fd7b54610f52e1ca8bb19da7e93ad820558f246c2b35d201859ddb81b2cda11793e7623df870d195c567047421d9188844cea1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50ea567e64266bfaf78843f22ee42cb71ccc4a07953e04d8079fb3629846eae6552db0dcf4d9b8f5f3dbf06599b81669b163af60a9f2d20351541acb3875ae1193be97970e301f363e290a5c10c64bc88b59b41a16958deb4860bf44f7e78b0f6bc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dd446ff34fc94daf853a7e3accd82b10250eda15e656bdb2273aa7265e409855111d42d8432718120c50eb5541a029c431c32e46d7afd970393d55cd19c7acb69e62f2190d5e36cf181553101786570e196638a0407f73504630d5f74cb90fc661b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcaa2ec305688c324ba13163dbed2d5a7d6b2c84575ebd0038599eed6bf4635e9082a083778c8c71e5a77ac1c9af313ddb76170ab7635cd19e43b2368d04c10e8ae0375606bea78b45d84357d33a7807f13da1e459c1194732afd2738aba66c8fdde1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6922bcc3a20201d5ce175487f1ab032d07da5a060dcce771295028c4cbc09813c6d847e989cd36599a46bbad4c8a16d7f237df3c03936abef3750fe0b2a8cd0f110d9c21ed26260a76bc5bb522dc08210e70f078b8cf97ec35af03cc9e134982258;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fec7ff49caf31550b734a2febaef23a11627863c8663cb865255329a638c2d56ff05fb26e486f66efb1d0d3c855edca86308576162e9233bbefc6b2707b612dad60119ae1307bb3de1030bd05812cad6912c9613533bdcc9b3797398c03124a265f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d761d4671ee6ba36368804352ed658ec809f87253bfb0fcf7cc8a7dfbd55c920bf91d0659ac501ea7b11d0b5405cb848210f6846e97684d0ec8df011180bb3141105ded800c78cf1a8172749b70b6851e69ec44f92da04630a177cb2c8dfff9394f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81f9e5d82d89f963b8cc9cce5bc1c82bda14c4f4f1b7e9fff0cb8507f18b82c5457470398a3afc502410a4a84c56a2f75346f14dd0ca00d0784782646a7cd18f2a24ff7f088baefcae7e878781059e2c685ccc57fef328c1034d924819eb1c2df8b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h670466c7f49f0c45fd2bc83f3962b1be97ec2a7d40b91c785bb5cc904bc8905a36693e70f75283f063f1f0e117e78912a1225bf6193cf6759e2a73707c5937544d80fd70dc9ce9e2cb452c6d354b88879aeab50abf976364e1c16ef48f4e3c5ea942;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11dbded3ecd4a444270a443b8f02852c7da4b7e705948f2df6a5fe4902333e6169b0adffafbc0f67586b01471abb5bf8bc46ca53277b7435a8562c26aa2e9b469a78c36910887457389895c4d9cd800624ca2e139240070f056f49fde9de6b3e81f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb7520e806038afdf2ab55b6c80fdcca27aabc3a17bdbf771ad90affc50007753e59c52c64035d1e58b04c2847f29bb562b80a8bd81aebd5f9dca7209247a71c490ab768c9ab6b032626ea14f5650eea92f3be997de2ed1fdc7464613259871ec1e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb45cebaf442d62c4044f20ad0aabdd24ef9286024a53e6744e6cf78bc8b9d0870e42945098d77ce4a3650a8baba64ea32e40de6936406ec813a906bfe6a7ce021bd0eb5d504e4409592a24854f28ea4059bb08deb4551c11bd7f4168476b1520d27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3115cd783afd79d42375614ec8867356b4c84800d78d590435286213459e50a8d864e81e90a7c76bbf052264a2af9b98ef605c1bd48d0f4cc3ee422ae8b139b3f930e8de93e67b0896cb14033ebbe6b33b42544702b6d3717b30151bee3dcb20f2a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39860c086c4f7d97db6a99525916232f435d7d25b1242bea644ec4f44644a613db7c651dc6e29eb5266613ad2c12167011b2cf929f7abeb6e23f3a6db4cad9d19712b455f38a7b68362a73974ca4272b4fd805eebdac222fbb4370822ad4a51ade93;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a48c61108c3a13542d7986e40778347ed09f95a319a48bc2e91818702a141502a6e160261532ba2d6289f93fd14bd1ef7da44ed0b8bf009da6e0ef5042010491145e9e05f7f2df66c8c1def5e4c4c4787f946172dcfbeef6064ebaf8ca22822a124;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e55bb542626c0af054271b5531958276c79494a5d3613d5dd56d1c26701ad1c84b1b38066ec7f7a35f18812fb3d755c4e5f184ed5b45d007c7417f0e7b8d69f2b8039e4db55d0886888f9809c1b568d597c1e9130f54086bcce361c6e6dbd443b8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7717f95ba923859a9776c04a5d2b63d1488bce58717cf4d543c916105fe583b21a912cfea23cbd24f167b0b674fa027b164690c7952919fd3202a54460abbf3de7f92123710003eadc321264296b7d88f795132f43afe5ecfd2c12001aa926c321a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91f5e0935595b1f7f8d2a2df700237a6be1d0e7082f50ab820414e7fc5f31a8529c1ebdc989e78e4a4455163db587fb4f50c76f285782dd00364f6b7e7f46b533face6348e6ecf7ab6e3c1e75100d2f35861fbb29fc8bd7702d4e03f378cb028390f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h248cab19602089ce5ffde716bbfb063fcb48127235ad79fd79564b22e23785219018ba4fd825d0b8bb989b27d1dcbd776dbc5bd747ba3bf1aac8d193c4e2b0c954c30acb816c1bbe0ba10d3c2a3f4bc4fbc58f6aa2529bab6f7dfe4bbdc27f4eb43a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33565541f737b6e7697b061ecb3d9c0029e637b07c7d8d744153cdcff32951a7bf2ab58e45c61157c3f3f10b555beb7a43c96d1c15bc5c9b271177ad458bec5c1c014069158f0c91a8769c4c7adfe41dec184469c06af802ed63f7b83b2056fd6353;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9840358b802501959fcfa3b705881d769bd15577864c342bb7ff3c384877487aa6b317f24fca9c6578a88654e33951982bd07fda8eec74ea18df47ae7b3b19b3c1204649158e7a84b35fcf07d0cb89aa027f2091531ba362411668f1b5530166761;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb609a94c1fdca72a7d157b1167d148d60b9d68c8ad3de0504e5452c7066b008409e174c87fb9e87d90921746007ee6e6cafbeba6f8f0403bcfbaeb47e5b762ebf35388e0ae9e09db4bdab27a4fa884d1a90b293d255f3d86b6fb5ebb13b58873c28a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d6be49cdc74744defc4f5d7a548ea3405c7ec72e9476727fac5456bf380092aa29da666f55b6b3cfc473fdf3648a99ca58b5ec673e96df819ba537b15552018d48b665fbb94fb0b2bb157647999ccfbdcd7c518ad884450cf12d6a47b633da0f1bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd76a599832842fbd1b0732daf753eec06f0982a2c0481862b8edf9493e69a64e3ceee178a0ad556bc0f933a264afee4b02e8618083e8edc167d6fc519fbde339fe1f6e12af9692861bc51368fb236e21f41e800d37fb310ab3fa47eefb3ce272adc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6627afe87b44aff04854ac97c45b25e0bb7b92b79b1cf556b546cdf17e907abed44a69eabf223468c2886f00e4c48888c55a8c7bc7bea32aeb111fdaf086b8f101196e8a34a0f7b9842f9505251023f4f7bdca22519f5c6b57d238e6a2a951a1c73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf5562982007df0dddd6e394bf18e46a07555ed57b59c9fdb31b3e20ab49f3c35a0bf0ee673bf2b58251f45533c9e4a41728a5c6a47940f46776cddb5c069ead95ea23193e31943a498ef1512aee436b5d0d41212358cabe238cb3067b0503210c7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb78a3008f1204e2f3e53afe07c0cbbf53d7aa471d3d0363d506d3ed2e3daa1cb95c570d184a39a8d16a6719ce36e267e8040eb252c70a90073e39bf5a0035fcfa61e5d4c72bd486a074b4bdad4e973fec827084a2f0646ca698f9f3db7795fdc2f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77eddde3ba6d1a358bce5385b3c5478cf0dcdeccd5dfb0c0a3b402c280afa0312b3d633725b3e77f2e60d9ed01f1b0fd47e8bb82d24e39c7d154849e47ca79568f77c30c7ecd87ad34cbeedab3a68148b5a739966188209c63f98f76e9b6e98b45cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb676c1828a70a79a91de3a7982e5b4031d6f72c10dfcfed0ee651f96b844c635b00c7314eb6aeeece27cdc88b5bb3858f50a6fbd38c80de07ae3312d91489d89550c3f70041f215d9f4740bed3085c8f8f16052aa8b167c44d8b904122a00def4cf4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcee19fc4feb42d3d863e453606e31f7d64da9513a3f4db118f0b695913d158612e3e490bd3e9162c16be455b6185043c2ead66cfc314e22eda623a0d6e98df449b3258787b88ac730cc259f5c649294ecf8c09017bea0099f42433f5a749a2c3751c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb116ff0d178c5d2b5f1586076ccdad51fba2e4ae983ac2a42ef72179b6e5735218ccd05dac240578ae00d6b0559e6a0adc0acb0c450fa2dbdca86eac568d2966cccf1fe0564dba717791d8d273122ec9f22e9b07a1a14282acf77c5ed5c121908027;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h427b9b9a427e78b2713e2d601da43f64fcfdb25e2b434286066c0cc0505200092b58199a68f51d3a314a9468f0ca8228f1b09b03ed94810751343dd51f0f3e9d96232580ddb9d6a8b170c113911cb7fe6ff34a6ece1208bce646527fb63dd5cb3c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeed21ee6ffb6d7a71972ef2ed499644446e88199ee0b225914c50e925e140b3c3425a7fb90c4d29876303095c6082622566ea94daef7a02f42f5fb2468e3a00a6660531b11b5922a515c8457d5275f3e5e11c81769cceab59c8a63831f407740;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c774d0c8771b537d9b025745ab650fc83f34c5c9e4191e15929001b024a4a630bc94d7593ff0091d6f55bab80ffa371a2625308866086e2311d18b133ba36574bb06965688fcf2b5f650757563bf20cdca568f6dc274dff6341524da665d6e7f63c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe36e71eca6bfd66063b5d186d93b9f792d7fc7bf01c653a752186a042e12132e0f8f05712ca8b8a88865218be74a5030c17f9f7506bd01cf0b3db6ce4a641ee873e2ffbacd87e20a0fe2125bcda618b93798c4d18282e7fb75916f140dd6b2445ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38c464dabf8c30734e82e6903ef963c44c7f570f14e28ccf23ea7e44c4959ef1205a1e37673db872cea47ed6a8a88911c35eb1ddbc6f9e3cfce12130fa6461a78446f8db116f65f77712587906174b45f7a74a87d6abcbb319c8665c07c7de567159;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h482e28133d67c9caef56af2d37eff50afea663845dd29737a12b0ade8520ad7b14de135f3ce3532481d0d7928418d9931a8fa3237e0683fbd2865d017301f1d8c636a4eced87abc65690c752070d601650dd199e5bdef775b407093c13d507395f5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbff7f48ecaa1aec0b4fdbeebec6b153a9dc56b4cbeae6d0ddf555b86f2f1629c1911c79f91bf77d882df8ea68277448574ea78456f91d1f1517d60d9c7fd4d84f1f577ca3ba92a16210ee81e5f04196e06b816c5ad34c4ee61d60ec6cc43e6ca068;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16b4c0b2278c319efe95165d3e3352313f950d409a497cc42cdbe119a294b1727bbceb60869236b0e4a89f637f5761c92cd749f430daac2add2df9aa936be8fccb3afa0fd18bd161ec8e6c8ae8a6e8553ecdb26dac2a7f84e0cea3d2eb6130a768db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha17a5e0a11362b8203af115fedb7775e951eca449e06538801ca53fb1418fcb4aea382b89b9e841594b12cdf8460fcccd59a093547d3c3e210d836b6af7f6db36cba44c5268215be7cc74f5f980d8e2e3e381a160edfe5b9a82a578924203eefc648;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c4d2ed43b1efe448d82a8864a14b64fb09fb234bf5aebd624f0831588bcdc42ae786c97cafdd19c900e8221732cf71c1544c3b40ff4d099e07768f58070414d92c3394cfdd231b1b2315e64fc7bce36a1fe04eebd7567deb39827e2d94459a6681c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3910f57131ee82392cef1a2b037c2f44ab54d4eac95cb23f97251c548e68ff5af2f47c9e2a141e770e8aaaa0528345a2e879cacd3f71757703c6599092bf6d479a3674373345b49f75414d44f0f52cb2dd1e3290bd1b18060781370895e6e2401d6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h500559c0f939403826f247b09342fb4d040caf54d06250431b0615e5c3e7d0b2c17868bb675a3cfdf56e589c32b92dd6f0efefc8fc11184d8e745489b5d1cdddac3f7cf35050a38400c2ed8aa89b119b1b232967e7dfd4347dc7f7b368132e67f3f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1fa6698e7c04f785826f30fb2a6def171c62fd0a686c4d4a796f00288e2e07c210167e09451ec8d0d58d7c3430d7334a0fbe0e8d99d42ba89cd96db87fb9cf0cebc8fb83c153c3495decdb5477e2833b9c59a945447aba744c77674a9ff67d67494;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82afe7c9994dc15c7a6e201200bf2cd2335b1f0dac9f073077a2d163e5e79b71f0d027e42f6606c1dbeae3a5b9fb4c8b7fd13d8bf48fc84597c2f1d4977eb99238a5c5e45a942e8b9784e308a164fb62980485fab923ec7e2600d63e5d55fe696fe7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dab5fc7103091f61be6f2d21023cdce5bb25423ffe536efb2a832eac8500e78fffccb29bc8efbdf0fa4c279cf6004e0f24d6cd8e21159862534fc07162a76f2aa1908a4ebda3a0a51093102b80c46541bf4ba9441891afbb996e0238d5fce62790c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h399c81133b52bab96934f46dda8dfe203fccf4e09aea3d215686ede2c0b30a283491c735d56eec27405c3e7e137b1b587e76c1aff18eff725e90c0e1b333d8c4f75ab8dfc2c0f95b8d7fb625ed4b8ff371fa24af3edc303fd1096c0e4847e29c4d48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h314b275b07194f5bf0185ea4ddf731699062775ec6f157c9156bc68f9f80f4aa1a87309da74ec03ae3965be58a21864ec48d3b537ab8e9f3e0e794d844d00a416a830953b6d9116cbf4972ebe25b73f0ce452f9249a55de522ef4d2b56d409b33da4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h846b4919d33e8b1fd5668f532896099da3c251326ec5a98b7df29d8a04f50bb5badc2742202ec931da521648c97a42a73eb7eb7994633be6a19facb0ca852287bdaab59b17618f62fc80d5e0ba8c26d71b6a2752724a545594f2ff8b95dbc130d2b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23b5fd565bc3e45a57e1e0bb82b0d97d18a81e2f3b77812cfd12f6bc71c3c7b756a6ee12325e32a0958ac61bed771edec72f4eeab7044b25b7b3f6ba40c100c6eec60cc26cd40374b53c9dcf6f88e8fa891e061fa819b94b209a299e309915d2a788;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a8ff550fe46cbffc843bda53941ac1ff15c2bf4039d361a5415f526c06d5656133f8d5722225b4aa23bac2309830c0cb29b5994a7ec4c756082d83abfa739ff89d6071b5042f8d0e452b75aa3f7ff3190f7c4237331355ff5b74f7b77484d343036;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h173514439d904e7b7ac0ef16d61a5450c976ebe7ff717dc49d33e4d080729193806e850a727300b27a836ae84e0c8cecc17ed2eb0faefee0ff72f6d01b147d75e98c4fbf8199b805c026a9b52e849177eed665cb7267f26ccde881fc2eed8d9d0f60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha675617b73dfde4eff24f2fa53a4d91b00dca8031fce5d5040c8c9b17d3e9ec2ed0a4161ce97f1331f7c35c9bffc85c2c059517c89e750a218ba13e25e977083729af4a99ccaccf9704dd74bffef79541b280bc39bf4db0344f901975a222b49e598;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f48b0d2d8f59f67679f2d7a3836f462b253c025c512b6f1207cccb015671877519e96b1b6cd504087853365396453a1494df315c3ff5b758a5e7b1795003748f05773b80de2955b6b14f4298ad48b61e9dd0e539514a2c71c771fc319e07331ee7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdde4c9d49c8074f70bf6b5e9d30f89df7618b19a3b5a3ea329755dab2dbe22219ac788e09e4ee31e766f7b7e6cc5048882a438f7c74d5cfa55e128eb04f6049fd77b0269b07bbf13b7d11788f3312387e5ddb11c41cbbeb3b9a3d205003ddf9048e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4a330331f2c6ad7c68adb02c54f59a3bfc819914c6e6a83a1865729df9e2f8b6ab9e654fb3071b08c0839d7273f3d7842df85ea6e945f8997cd0a5e0a883acd36ce1c78e9ca12b93562bcfd862719a77d0c2c22cb28d0786b17f46b96927b86e4cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c8d995e74b7f208a28d0f10fe4392c1dec769a08c1ab61e879e660c7c9b1c53fb83b1357c3e99b08b6f650aafbdf64701e108a1d920d97b202c8b2a002bc0adfa17a09931083b9227017120deb783da99dcfca13f6fe8eb424b063655509f9308dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb8ee9f9422b0311137afcacf774783e00145d7c6fe01ea12983158f2f0245e1e288708e1c965b16b06604bd7dad18d15ab1c67df8f64f4aae2cac6b20687246f2394240285540e97b5a6403e97fc70f01316c70f9f14d3a25d9a4a04878ff0a6b39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cbfbc9f26c88001c078eeb681b575c221426daf881f35a72d282c8c3fa1227fc7656762a1d956b3d9f87fef87ffbd9bdbae7bc22c85e60ad79bfe3c8ed18750447e1a3154c89c2d54f3e4c500490c6f92921c5f1157c93879d07b4289d1b27c5a04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d16dd04c3e2c7f25dd7da5ed1f4d2ee901043afe227e4037b156894f4f12ad5eb8e29767e1c5d26d9ca6a21b1c3b66d3d2899469eb86131baf205824ef8a6334245af4b2d56a698b37fdb295178449b5fcecede7c4cce1f222f5d7df3ab773b91ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0aabe4c28584e753deab731c5cdddf2d1ae41a0aab126632ebf6c4feade4ffb77f146e141fc4a4697b855f67653a92609f9dd63ab69f02f6177c25e1359dfad3a5e74607dc1c4e83eac6a0466d97ee88cfef1c8663d5c6df330258f0d67d5e43526;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63e429e3a8c52f578d987533d2ff55b6458e584cf17f3dcb1377ae694732f8be6e0a533514d760c65236148132aa61f381f0cfab996341c3fb6651f6b7553fec32d45cc0792e69848a8a9647b0cad97c7a71dba9fd6401c567b865cd595c0e14e75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dde149e682cb00a265a0613fc492fceda26b2c0d72fe4529e294287d62786819082d296714e23bf6a05901518f9d46b5034ada924a6ec6cb96ef1795cade8aa27080f26541b8d08f367df92cdd24cf6352159142d064915869b385bad4c239afbad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb518bbe0058edacc0c775ddfbcc661b6faa77fb8c795afecc040e35ae958c06e2c313b849b6a7610b7d6f45245296a1203e10e47324a952ae427d0a267dd432a8d67d4a82865accdea2277971289a8d96a2b6780b28e3702f1d1347281e40a8ef161;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2934c3583b5ed5298a5214544b20f9ee3cc25afd0b49fde628c3041f7ca2eaef5cfb96a5de57936357d91c268f511ba682821ba5747da980a217fe03136a578a1312d245e04f4c8818cf2b901fed710d0812f43eb7e78290c1d7234e7003e0b36e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9f1f8e3690f75df39b4b271a7ac30b9b4332577fa0e2b42e7656d116c5e694b6a36a529b2904698c752246328819beff8632039c8d4ecbc300ae9d79ae91f2d9ac160207bb285d0802b7219f77a2ff6c2582af35bc9a42c7bf9c9e36df4664870f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75eccec7140ace07f790c5420c99b9ade5300d273dd96e7e2998c914dd947eb5af5f676d2797ff5215b90fc83c9a181d40572e051acd7f8eabe269dd6ff83efadbc3b88944b04f441347f1b6257111f1012ccb5f8b2ac9b5c238d1cf0473280df3d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1745d2da5ca39f7b3a12e4e6942bc7b93c7246cd18b1652af7fe1841f52af1f6a3b849249b1880aa15b6d09cd87bf682b1849252202bc44e78ea5cc80834c11eb1ec279232cbaa54d36afe95fe5182401342b096909ce1a6fcefb45bc316718c8aed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f2b3f458ff745875bbed7a341e5898674ec7c20f9b8c56f0a03c2219daeb70cf38c02a3cf6858ae5d851746dcb23314b593122f2ddc385bc9c985baac23b3dd57ca86f03ff0d8da088707b71fdfcad351cd491be93ae86c19cfa8249f523c749bd6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he185b196a86630710201b25efa80f83a743eb79534c168093886014461e14a30938666918c551e6603a97860b169b7f7d0c911ea3b6471e6e7d7174ba50fe288e44acf93b7095c2a8481d5c880022df7d0e5c5221e13c2bc867a2b15b0a34909ef21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfafc1a71c7cdc3e34a4565bdfcce8a836b087d2a088ce113551605a01089f8d75ffa56005e2dace3aae2ca75b625e89fd5908c6a576da72ebf4f2da878627e8f8400341d07c7ec7ec75c4c1b4fea24da4b24319d57eff21b32784b48033906fb0da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5c11b3d24e4e35bbaf11579f9288cb4b33bd32437f7bee305cc72735f3d194cf1b7ba889bb6db167270ccbff8e7727c2291aad3553856fdb510f7ac17bd1ade3b3c0fd0e891ea9a392f614bbfe09d358c617e06fcd0999763b4edce1b94d865f770;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he48251145a246cc4904aed1d021d47a48af88b26142f9bbf86c86a70a4571378322e4424da7c7eb3f51e4c74e0f24358090c4a547983cf00ce8e261e203836aed3a7c30ce697a26101a9b2d6605f3256a2548b4e8fdfb31bc99e964025f44f9ad5a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd77ecd04e6924cb4ac4018cdaab90b63776c236db2ce3d2242f0bbe3a7a6505ad9962a2c7b8293eab00201306aa0c87efa9448467798fd5fb1603235aa7915cdda2427e674e4562188df30b0e229325ac608a1bcf29dea97c0b97807b1f530e55ba2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffaeab86f223ee5df0bc0b0cda77a4121d16c71c6870d97b0b84c094d518385b4b7cb05ca6056f69f7cacf4eb19681178ad9ba6a4a620f06b9a9cf123c17cc009c15bfa76e1f9b1989692486b159444e9b69084d28f9715125c5933c9e6e49ec08d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6db434566923cac1b3e20923c6b6ebeadfaf44e1096fb170be3ff1e9d425e002059dbae9bdb8dcba46b53ddc6c7d109af9f851f6a3a158f11ed7f03d74b839733bffabba63bdd6e6555aafcda09abb0d9bc41dbc2d4d3f9d9623854fe06baf2ff8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccad7e31dcd7fd29d395e3f71c102f251d56f5a34388849b9c9b5abc896eb963d61ed4993a04ded619b7dbf384add1be0e14b5dafe7e8f4b1928e032953ca81d67a99f0302dcd10cd8fa24bf45996c8b74ae88f5067705b64a92fa2a2efa59f61b73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4c93687f35ee808bff9ff65d194e0ff29d5b6c526a2fbf7d58235100963633e930862a3b529529de163ad53ac7c076d7fba5edc2fd514267686433a8c58360cba981be3817008b11fed974eaa865f6f1d9b3fd52a871a968ef3b74eeece2e8f122b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2724cd9d943e1448daca5cfd926df3116902b4c9bad32579b95374c13441f2f6825b709eab001e48aa5b792d0dacc166ba220d19844e4d6686438840fe64d18d111de29dff72ba539b6bed952951600bead13745d25321a704eb8bad233ac595a17e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f2537a7e89f17d83120a7b322df74de1222e33714bb4d0ec8b4619bb5a893d82dedc24a63d155f86fec8347d7877a2cf7956cb46b2ead8accebf1744a14a14b147b198dff10a46598b1d81f5d72fd06a31e2fff5671199b06c7f8abd91e612e045e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeb8e95d737c10dadb136efaf0603c876def17082edf8c63ed8f6cf13b65e5f585fe98010b3d5da2f8ceedddc967445186a93c01c64ee37135831d749e6c0f233d14d08231d87fdbb7eae230623a226cc068275771385b9aea468023c4c14a630aea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5723610073a53a1e4feaabc794db8e8b4987c5c246f6515446da5b25a4aa352df47a0ee5b88131e901e43bda70f0c113c990bae68f853f8abdb14ce183027c2c4b3b6ba7199f04cc6d5885789c047da3c4b237d41bd64c9e44083367fd679027635;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcc2e73b324e9355a7011ae45efdc96aefdec3fad9bcfc251782ec5472a8b9bafdf01f105a6fbd4b5586036055a5a93e26e051e770dedcfafc1f4e9d75911911adcb84f1a7818d8aee24e45901f7d4542795b9a5895e884dc9654ade67c3886bb54c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddac3819f38017c6b32fbd44b706569c92254f2ac23e45df8f39d8dad3fca08f51afab3f91d01d8a3cd1185020ce251ef21f2f70df415ca6150161103fdfba58b03ea6f36292ccd4ef9b77fea444d378409ccf1a6468f1e01f137e879490c73e8fb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff42775556b0a5f5d2fdebc8ed0e8ad5bf888e736e56ec4af86c92e3f929352e81fba893d32cf741131a34163c90d67e510ae52d02fa117ca31349418fd1c19ed09982fa8c3bdeb23fa8dc110d295cd0141d956e013ec646bcbb7346c6481bcd07f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f1454d5c65ec16a5ea1099e7741dea669d8462461d62ed536e48fe41c6d0fd3eec74c0b1e2c423eaccd2da918a957887155879fb803cebfb48d9a9a467c75084ad0ffc970c507100e6690b279ce7d2eea1965c6ea7f70154c0ccd2faf5459470b3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72b767fcd3946f5536c347b9e6b1df930a5923d8050ffa0baf275b5c224e1843f40f9c520783840ca31fecf4b7a711cf5feaa0a921f17889d56e1bc228dc29b2026a9390bd73a1c2c7a28f1f85d7c07efc00aa766767e6f0be5754c43e233680ab56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e3a19c8fac44f681499f21e03e8e2ff3564bf66b1285c58958ce26087697cc4c8bd81f72c595141c37f8804feaa3c52aefc8ab66f1fc6447ddb635e37d63672dedcd7067cd6125bc8804d358182063dded3c2896e21a914c6ef080cfeb2c6807b21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9534be427c853e32687e4417d17e38aebf3379b222f425a2138a97d3e3ead731e6e052eec36f8145b59b932b07c56cf56f7f2ce0c75547b7e87587ac0601afa484fbe0c7b3a0bc09a584c3207a6206a27471a2c5175a411ffa00ad358fa4b1ba97d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc385ab464018b8a5fd5a0f9dc184f184dae8103631dc415566b01eda9dd0c9fa2fbf94caa77d9c7ebe9ab0bf941db946afdcc6234959381865befb626ff2ae6eab12308ee8757f5af0e984256fcce10f075f2f71e953e02d40d18d210b6161f60df1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fc48d877e4d48aa268b305932fa0e274a842d377dc721890023f23b58a2fa38b58e8dc2ed5f97ff6546c17d37dcda67fdb975a6d452c0c7dddc9bea3e66958a1673f051c8d9dda4b6ae1916138a40b4e276ed705f062f271725a973762b2aea5e07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdead4b0c6ce4ef2fde44c36fb14232353c2c4cdda206cdd6f90ae13315347269c63f090d9d11cf64850b72570ecaa11a840d538cfe5ed08552a991b86e1f62afe0389c1bf4225ea06c7d437e4143e0a1a58fcb03a05483894ff9f66bbb275c374a76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbde45b810496e6094e6ef4118b2a29fd756ea6c9127bdd7d504b8edf6e2f2c46efe3a20c843b2fb84046dda2da8a114716378b0f7b7bf6c2e1378a1f7a593a0b210f8d1f0a8006a11ddc8c137e5cbfee5afb2ea877b1cfca22ed52184b5c261102f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cd5a84405da24498ae1019d41763eadaf51db3a028e653fede92c582df0591d92d77aacc4638c956b91746ce5c8b85147a55d713a1d1856e367d1b95ca4a122522783eee51eb5b4484969bdc7ea38cb253f82792100ce43ff5c1aa25ac5c1bec28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3442d2dc0f07bea5b5d4311e05eaa2a7852fb2be228a9bc60dd58aac3e5b80c5be9ecb157f41187c768c1d0eec368a8270c2c4469dfc747b5ceb1a6ca63f50972e960b4ce911251af0f3d60c09a5b8bffb264491e0c30d2ce0f473d9ef3183558a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc92e8ae7fc141489467ae5c27c934159863f7f6e2352f41ce765acba4d94430b8bf52d3026a001eb6ae2310ea2772716422ffd3334d0396bc270bbde723dbb3c743b87d79b14a79e13ab640a55713719e08771aca8e6f784d168a7ec4edb015c725b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h273ff35a72027ea904a645fd659d2192e8ebcd78daca1d67387b0b006461df7d10552b4d6d697e2254f8605ebbc5c03923d27f6786cc749c9f65cf215eed35c256a21124113255a2171c444bad21d1747852852ffb0917af0e42a8cc79805d4e446a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd058b7c87f4fd1af81c20ad722f1bf95ce271a2558e283bce93284c566c5528f9dd06705a41df58ade392fddfb14cfe7ce99fb04ad91831ee7cf654f7f859c1fd7c3b148ac6ac2de3710e93fb7c9b7732d96d3d0e438515c67052d5fa36a83431d69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93d71d39f2fb0ef74cc3ff286b94605181ad3284824857fd66c2d77303b89e0b65191ccd12c1696cfbb2961787890564c148fe156e0b0e58a5b1b219ff5e2eb9c1da6a02cb54f006059ba659f2caa9623e43c91e6a734372d8ff542c021cfc23a788;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc40dfd2f8ae16e78518b211c91a9586f6a0832a1f1b59ed7901b3d34bdd0ba12f597f4fb6e051ac6dd0e8f94b5fdfc08616fefd06bd4b2ba8afc83f9da56f23e9ec144c27b72e80eee65e6a400fb432bb07554919054e05bfd78025f10a0b19200fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56e9b2d391e5424816102244679700834c6351dc14a103ecf55cfe700b1e55523be97660bdf288523b0ead173d427d551f40f0e6e2c0887b5138f49162063fd23b2535e113c21e6aa77c58638d115b7dfefd101f8f131bf03a22fe3e18ea11278431;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha27a2add1aace258639c42577e18ee2dd4c991e48076e355947b5cf6858e6c72f91f3718a1cb758500992dd5be3e8c1c40164e70c1017920a3ddcb44867c60b4336087cb35a2541a82dffe2a30cc07f1dd00422dfccd24c5d1a653f54c53f23c34d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h479482f6ade1c8467321103e75f8648927d98a4d149bc67ced6ccada867d3c81a76c9ddb1c4d20e43c421bcfd5b23e34ce8126672659c4c6f926da973204f6143ddb6ca8973dfeb6e8fa5939cdeef19765b46a629441f9082e135c24e00e85acb735;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h711eae03cce6bdc0c1afc46acc812694075aff326d4cc121fe82f5d2aee6821a5399ddd7248639d7d6c6dc73dc9930d9739a8cb5855fd5efee0bdee75d2d60d9e6ca13504dd8e5eed4200ad3d7d210195dbf02c2538bc0b4a8fbbd6ccf4696e7cd19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffdb3ccad7122c12be9d7f43a3e62d006a6d37f348a76c939c79be2974f432ba5927f29325be21c518a98488eb32ad84f4138f50e64465387eaae537e0c427fe9fd3d78c12b8b3a490731cb8617594e1fc38a24664a1368a0d86fd132d962bb3d639;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6be0e8c28fd78f6437d81f5ec339b8e279d10d48425e64ab4160788acb17c82982deab740506b45f3ee6a5aab4745472940adbb8957e3609d44dac6368447bc037582d351a35e82efe12b5fb169d8c9d1f88a06e99a4688ef074b09b2d1cee1dc459;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a24a5ccbdefd9a2eda5c96cd995c791354dc698d2fe3e20448befa9dc09cb5564dc611c91aad22f8ef4bfa731a9905cedac260f4fc4a049ecb9dc8cf036b6f3bfd7f5761d77823dadf028252feb54ab6da7d14569a80e1e7d42f29cba7335e52e83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55728f2c6954326aa95b7b58f0f5a6903dd5e111e6c83f4a572a0e30fe442861dadc530a65a62ca7886b0bf6107f550390af8dcd17eca3054e15fd9791dff4c0148df7e24d652e929b20037738af8b66657ed9b888f6074c27d8ee50eb96fcb196e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b723df60fbbc793bf042e4c211617628285e90e0013445605131b5fa66700d42d5b5b547d8524623dc6a18ec4a9dec0c96c36a4020dfabdb07c16900ec593d7507e670319b4bf2ccb4d41c6771e9f1517873c3adb4bcfb776831467a0667d20683b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71c6b4593b6418a2c10f93d5a2dac16371ddc91465819139e51dce58d8cec626f569ae128d8a55bc673cb47a51d3ca1947b83d9069515e7e179058ae7bd0dd08a2fa2968ee6b910d94ccfc372d864edae5db75df3bdd7973330c5f179710bc28eff7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc9713a14d18fecb2f8236de1fb82c77d28a85dc92ffcf4830f37544034900795e86c0e0f08293e5553be09ad58fd5f721f2e2adca4631b238b765d824f4750ab3b9cf6790d0e5ba5dc82052ccb8b00fcd9c30d82da1cd035556031158321da70aee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf303d99bb4540d5a243d3ecbfe439969df5c9fa3c8a203f19e419a1354d897187cc664df4f4ce1b00e288604631841eab7862843cd481d60ce42edd842ccf33e479fb8cd81aaf3db152d3c5f3011dc36253caa13b0dc6e1ffb60abe61e9522c68624;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h232444d389a34ceda55c735f5a167363e9e3916e4638cd590cd6b90d2d72b303c026784cbe9464ad3d872ce78053715a07df27731476415edbbbfc507ded7fb8b1f6fa65d969058aa00ed63945be48bab0e40b97e30c0e9c2af0cf3a605017bc3049;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he89ec7c7f734deb858a1e8ae28239f04d7fba089026df26cbea3ec9e17019ccdfa2ba3cc6a0baf9960b069f972f69b78d27c2d2d2176978e56ce10b59226e56b2f70d658aaef8b1d54ffb44bfcefc28cf6ca16f804afae34d41a6a51f779396ba3e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c339cf5efb2670a48eac1001dcc489053218f49d97f39495fa4e120629737db31b8f9644d3cd9e21c080e42fde63f608e8352b18d41d1267a95ad0c91aeef2522ff8695a92c912600e1c312da52f5f6d87122fa8b5da6cece608b36cd14e53aa010;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7e5b3487b7d7e50f314ae2587aa9f2626655925c67ed217b8e298711ca1fc28a5c0c619ca016d0d99ed6b86853e3cea2d2d313d356c02cc2aca65b1fc12c540cc558482ec59b4bbceeb1eb094de573b9b76c40a44d5a681c06a25fd077c12249482;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a4f3e6d433bd549c30246ee0efe5e3679a949dcba69fb821210d463866593837fbcb7b250956b265f87731a996df446fb36814ab7b5b49f035d07dd1bb95ababccb73665e2a214e8d2a172e6f3ddc8a4e98ad58f0ca3ac70501351907ba3264f360;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc13890ab6574e7ea5c9e33120a8982bd8688cb1f538d277635ea9d3b6806791df50559f95b327474072903e17af60bd0287c2b1431fd67033487ebdd170f7d7394f7dd8385f53e7e28babc948e4e38ad74e498eaed08f596efb0cc740546f85db673;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9277be01be14758e0989f5a260b0baa0d5b15e3a2e6b3048b47fc131837396b2a5d756089ecd7e7f00da5e56e1c00b2cbd9005de32f88ffa12ac857229694d76c50770338d274ac53295f1830fbb0580b6db226c82debeb16f0f2c6ee7ee00ad71a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc581c79fd264f3aba134150b5d3abb1e4b6f25fad9d9394f37f54830328f3597a8843323ce6edbcb94523810f4a35ee46a6237234f3a414137babbb777127856fdaad8b72160347a18c716f4e6b280a62dcaa954646647d2970f06fbff8d3dfab34f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ec5e844253c76cd43d00b45904debda2ccd74a2e62be7a5ff0b6b4b1ba0153d0c9d04f24a564b81e86375bf4375990b48ed945f007dccc1cbcea1d83649e75fef09e9c52c886869be787eea6d98ccbd31d96bce71fc3eb916652a02c56128fffdea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h176f28ca9ef453a9afc67d94ef0b454f4bcd99b1f33a44e7071fdb77b4634f7e26139f5be912156675f1482ea54e5b0a498f2ce39e389579be807de7bd4ea97ec3c42c08d0ac88ed13c52a520f299dd56e60db6e6e360db7c64cb1baa4fff20fd169;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7970e8e46d4ab3ef1ea03634863a5e735f116af97410d0db6a810008d09e7cfab3f895fadf22112a77ec8f8ce3a9d19d32223d8ed8d41a892d766ec6d4fafada93827e71112dbb920fda9982665ef5ba95d4309863850259cebf69ee6f93d6eeb42d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4125fa8b20b13731967b2786202f712d7a4baa7944042f84e8d0661465d272bd2105ce8fd9026de38b537030795d6c528959d697c3baeded7ec9061ba7da0d0c58a1e7246c9b901553d7eb5c36bb2b65549516b2df5da7533e232be0bed11424b3ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96261422d498b46ab5202dd79fff951e98873e02522e1e2124b9702bd2c1f37fa5e127f5286b233123f5db1972e6a759f2cbeccc0dff52e5e4cc504933f9bc6a7daa6d3024b67d26c04695026820c5eee87c90a6cd346882e5fa1788e1425c2c813b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6199c426771a07e230190ac7b0f80923744beb28263a658044d715d40a7b91e75c0839fb03f26f7671f2531c4c5528432763ecccd9dd15406f0a83a9c74c9aebcc7f9af50312f4c50cd6ba8ed9fb85763cbf35f9fb86cdee69f764b884ba6aca2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9af3112daf02c206b67c5299150b5a2d1ebce389957de22d501fd7b25bba3fef8042c3bf1ead2c277f8790879d4c58bbabb2d951f4f1e959ba8bd3efecccb7fc849604ff696245b6792b516aeba10aa231da77aeec4aa548d1db33905d6f4f715ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67a0e735be845c5da01855c914dd9183d4fbd538e9b7678d852c588aba4ffca1529f2d3f847f56d5c3cc82aebfaecd632abf590a27c5aff9aad8120af0d95c2223d8a9927b45e706e05a830029c1c1b482da85177bfe8505ea78da47f2720d7710ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2e72f71e709a428fed9448b0c309c756185938876938175eb6c358c7621bdd52cfc719f88f4e66553ad939d2b7afba180417687ea639a857d219ae004d07a154b3c4455b1560604d9202bb66a08f91304d69f9c22dec73861df722dac94cf5bfe11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha99bd5ee93dafbbd39774f82bb61f7daa03c9ea40e4dc1cf86d734aacc9990c2e99b118162ad573abebbae2beae0fed8cfd91be29d94cf2f81762923b1676b7422b13d4d7d861d955377a2e21daf0a248781912d3dd73f96e03bcb118ccdcddd514e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88edfd5e8dab2a82499d5bb2c4b6408a1517eb047ac80680c8970e12699be24acbe54c72159c3db12d012ce22b75e3a68f4f97b0ba05ed97ea9ef0d65ffeebf5cd1918a779c5c47abccd840493076aa0f17b7e1cfbb2497b2dd5f2221a7140ecb8ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3535e1001ce5bd449f5a1a85d8329edf4908f83beab762a1bb2fcd46969da319cad3fb1eb7f0f5d7ee8a838bcf3991432c5ff2d3c6c6ab45940204dce19299ef1b03f5932cd33f85840b3cdf9f63dad34a0144c0e80a3b1512e7bb03d25164c16364;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd39820f83a188a3461bc22fe21a274822f0e8236ae784ef1c0ac87e81c3eedee9388560ed6f3311e9d3552d789e747ad322b7b6d48e804647ed08aed9d3470c1a63f842b2f47075faacf2ca21408c1ee9b775d64815967644565111f9a5ac25ad18c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcefa31c47f6551aa289173cfbd79ab23091a710d62ca2bf2d78795315ee5bdd7f2d9f86961aee4a4235f75a80bec77a36e553879125435bbeade6bbc012940a5cedce38fbbdd3d2243f0be3cc2212e44fd51aaf40ff56dd658c70f3f1ca10c0da772;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc87435f17ffb2373c9f8ee5c61965183e998d817ac73c9a634becb9ca4a14e3585b80f0d1d943ca0b54cc80c43d1328dfb497234931adafad02b741caebbb845a261fca4298ad37292dd253c8ea39ce01136c8e0a786498ba1067f08553d3fcb69d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea6d9ec1676e7fbbfdc644278617db4d7bfcb478cfa9558a0f6e309d284238e1758a8db14a3b2857d8285dd5d1fb1bc9831541944593477f93e5456c8b41aebf864505e6f49477c5da95a703b12b5704f5a62e947df572bd0ef2707e2147c84f9dde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h293a0441cbdc16ece69477b02606bfe8a712e0a933826995b49438dfb79c349478928184ecf3e0a8e46a3d0993803f84ce4e8fe7bf99fef396bec6e9119f9a06c674a70a671fc3c9eb2c8a53c2f6ad78f1aa3c39b3205296a8b16ca3a1957a81794d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67bf9deea9274b25658390eb559e6a44dc231b65f631d375e4a7803cdd3d0ad6a18c68c3488cec7d1f0c540a8486f9191891ef1222dc8e63ca97d76c42a3ffb417cf1c44b7fb56e3f85dc428b15801a4513f163024eb945821c9f36723fc2fcdeb55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0cd13a93ff0a980669e5e659c3d2a3400104b73d1e37710237b33d7fa6c7395eeee1cc1f064d1c16d5dec142f1db3f5c4599dcb78e1e0fa88d5e402a92eefe954240d383d9ddc80353ae9306d28e64e2b4d8ea189dde3e81f573639f1d75420a2c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ce13993ad705cdf71688f2ce267e3ed14c7ecebdec6f60766c24926a4b03751873fc387f31f273615d377967ba556e64be4d97a85f4d32e450b708c43c45a6d9487a4ea972dadad5356c69af1d4adf240057d2d35a844716be113505ef8e0f1dcc1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53f44f9e277c9d5c4846429c741fa6be089934977f8ab956c8a83c1e7cf55364bd64558d87c031faba310edd4b571c81918aa3bcb261a3fed6feff93a7bca9966fae4a6f16fdc5e4250333c4782e54b98267876f4e3a0b67960289bd6bf72edb5876;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b4a2394d16b615e6bf061578cc3cd267aa4b019ac997291050e77de9a469a5a0bdecdc4b23a6cd13998c99b083ea935be7d948c733d4d29dc72d1014657caf46b65f22c08b5c55fe2f3ffc8d863dbab201c3a0c492507541513beb8c23d18f8ead7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9621c8b8e792bd3e993bd108113999a84821a85a744015f299ffca47d5ac120ae8f04c92a007c4a1ec897840755591b1b67187166681907b1335cab478698077de4105d922bac215e0422f0c9899e9905bbf75415d4b74b19a97103c7cc243db2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7fc45e0899467c1e60480509f32af71c9527150206fc2ce6978fcac446b5af67657581c5c7599693a41b1d9fa9698241e59acebd864a02715453462682b0b1f809a7977e7850c3476031a02acf3db75ba4a7fce4006789094990f108141b182a28e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2edc0880452ac91b908a14f784b92d1d052ffe25fb477fe4fce25243b0995f96dc0579abe5027735074c693d7badbcd6046aa7586e8b25ddeedd9201f78f182f065920e027d7e633a151c4d4b5510b54a1f0d086562dae90f6844fc1d45d9dcff2e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e25ac73d70b7ecd3690649afe66db332925fee8c247211ebbe42b7331ade52b564aad1d1d9c8108b2f8562b4e6ff1700603c5306bd3b2ac271abb57a8814e281f24461c2cd5f63c04b3cb9aabf82123f3683869467ea8afe5517826ba2af44ff720;
        #1
        $finish();
    end
endmodule
