module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    compressor2_1_486_32 compressor2_1_486_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_486_32(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [0:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [0:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    rowadder2_1_41 rowadder2_1inst(
        .src0({comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], 1'h0, comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], 1'h0}),
        .dst0({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [0:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [0:0] dst39,
      output wire [0:0] dst40);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [126:0] stage1_0;
   wire [137:0] stage1_1;
   wire [227:0] stage1_2;
   wire [187:0] stage1_3;
   wire [225:0] stage1_4;
   wire [217:0] stage1_5;
   wire [246:0] stage1_6;
   wire [223:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [187:0] stage1_10;
   wire [219:0] stage1_11;
   wire [281:0] stage1_12;
   wire [204:0] stage1_13;
   wire [296:0] stage1_14;
   wire [171:0] stage1_15;
   wire [264:0] stage1_16;
   wire [270:0] stage1_17;
   wire [200:0] stage1_18;
   wire [299:0] stage1_19;
   wire [188:0] stage1_20;
   wire [198:0] stage1_21;
   wire [250:0] stage1_22;
   wire [177:0] stage1_23;
   wire [211:0] stage1_24;
   wire [234:0] stage1_25;
   wire [214:0] stage1_26;
   wire [158:0] stage1_27;
   wire [251:0] stage1_28;
   wire [235:0] stage1_29;
   wire [171:0] stage1_30;
   wire [160:0] stage1_31;
   wire [150:0] stage1_32;
   wire [80:0] stage1_33;
   wire [21:0] stage2_0;
   wire [106:0] stage2_1;
   wire [50:0] stage2_2;
   wire [87:0] stage2_3;
   wire [90:0] stage2_4;
   wire [83:0] stage2_5;
   wire [93:0] stage2_6;
   wire [109:0] stage2_7;
   wire [107:0] stage2_8;
   wire [74:0] stage2_9;
   wire [88:0] stage2_10;
   wire [91:0] stage2_11;
   wire [102:0] stage2_12;
   wire [101:0] stage2_13;
   wire [138:0] stage2_14;
   wire [135:0] stage2_15;
   wire [103:0] stage2_16;
   wire [121:0] stage2_17;
   wire [81:0] stage2_18;
   wire [109:0] stage2_19;
   wire [127:0] stage2_20;
   wire [78:0] stage2_21;
   wire [78:0] stage2_22;
   wire [109:0] stage2_23;
   wire [99:0] stage2_24;
   wire [87:0] stage2_25;
   wire [98:0] stage2_26;
   wire [96:0] stage2_27;
   wire [74:0] stage2_28;
   wire [120:0] stage2_29;
   wire [129:0] stage2_30;
   wire [83:0] stage2_31;
   wire [64:0] stage2_32;
   wire [45:0] stage2_33;
   wire [35:0] stage2_34;
   wire [13:0] stage2_35;
   wire [7:0] stage3_0;
   wire [17:0] stage3_1;
   wire [31:0] stage3_2;
   wire [26:0] stage3_3;
   wire [43:0] stage3_4;
   wire [48:0] stage3_5;
   wire [42:0] stage3_6;
   wire [68:0] stage3_7;
   wire [37:0] stage3_8;
   wire [69:0] stage3_9;
   wire [28:0] stage3_10;
   wire [43:0] stage3_11;
   wire [41:0] stage3_12;
   wire [40:0] stage3_13;
   wire [50:0] stage3_14;
   wire [89:0] stage3_15;
   wire [61:0] stage3_16;
   wire [49:0] stage3_17;
   wire [49:0] stage3_18;
   wire [49:0] stage3_19;
   wire [45:0] stage3_20;
   wire [58:0] stage3_21;
   wire [46:0] stage3_22;
   wire [47:0] stage3_23;
   wire [40:0] stage3_24;
   wire [39:0] stage3_25;
   wire [31:0] stage3_26;
   wire [66:0] stage3_27;
   wire [42:0] stage3_28;
   wire [38:0] stage3_29;
   wire [59:0] stage3_30;
   wire [39:0] stage3_31;
   wire [35:0] stage3_32;
   wire [39:0] stage3_33;
   wire [21:0] stage3_34;
   wire [12:0] stage3_35;
   wire [6:0] stage3_36;
   wire [1:0] stage3_37;
   wire [2:0] stage4_0;
   wire [8:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [22:0] stage4_5;
   wire [20:0] stage4_6;
   wire [26:0] stage4_7;
   wire [22:0] stage4_8;
   wire [26:0] stage4_9;
   wire [28:0] stage4_10;
   wire [20:0] stage4_11;
   wire [13:0] stage4_12;
   wire [27:0] stage4_13;
   wire [12:0] stage4_14;
   wire [47:0] stage4_15;
   wire [28:0] stage4_16;
   wire [34:0] stage4_17;
   wire [18:0] stage4_18;
   wire [28:0] stage4_19;
   wire [25:0] stage4_20;
   wire [21:0] stage4_21;
   wire [22:0] stage4_22;
   wire [21:0] stage4_23;
   wire [30:0] stage4_24;
   wire [16:0] stage4_25;
   wire [23:0] stage4_26;
   wire [27:0] stage4_27;
   wire [17:0] stage4_28;
   wire [20:0] stage4_29;
   wire [22:0] stage4_30;
   wire [20:0] stage4_31;
   wire [18:0] stage4_32;
   wire [13:0] stage4_33;
   wire [16:0] stage4_34;
   wire [13:0] stage4_35;
   wire [9:0] stage4_36;
   wire [1:0] stage4_37;
   wire [0:0] stage4_38;
   wire [2:0] stage5_0;
   wire [8:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [3:0] stage5_4;
   wire [8:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [12:0] stage5_8;
   wire [11:0] stage5_9;
   wire [22:0] stage5_10;
   wire [8:0] stage5_11;
   wire [10:0] stage5_12;
   wire [15:0] stage5_13;
   wire [7:0] stage5_14;
   wire [10:0] stage5_15;
   wire [21:0] stage5_16;
   wire [14:0] stage5_17;
   wire [12:0] stage5_18;
   wire [12:0] stage5_19;
   wire [9:0] stage5_20;
   wire [10:0] stage5_21;
   wire [11:0] stage5_22;
   wire [13:0] stage5_23;
   wire [7:0] stage5_24;
   wire [7:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [11:0] stage5_30;
   wire [10:0] stage5_31;
   wire [10:0] stage5_32;
   wire [8:0] stage5_33;
   wire [7:0] stage5_34;
   wire [14:0] stage5_35;
   wire [3:0] stage5_36;
   wire [5:0] stage5_37;
   wire [1:0] stage5_38;
   wire [2:0] stage6_0;
   wire [6:0] stage6_1;
   wire [0:0] stage6_2;
   wire [3:0] stage6_3;
   wire [1:0] stage6_4;
   wire [5:0] stage6_5;
   wire [4:0] stage6_6;
   wire [2:0] stage6_7;
   wire [5:0] stage6_8;
   wire [4:0] stage6_9;
   wire [6:0] stage6_10;
   wire [5:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [4:0] stage6_22;
   wire [8:0] stage6_23;
   wire [3:0] stage6_24;
   wire [4:0] stage6_25;
   wire [11:0] stage6_26;
   wire [8:0] stage6_27;
   wire [6:0] stage6_28;
   wire [3:0] stage6_29;
   wire [4:0] stage6_30;
   wire [7:0] stage6_31;
   wire [3:0] stage6_32;
   wire [5:0] stage6_33;
   wire [10:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [1:0] stage6_37;
   wire [2:0] stage6_38;
   wire [0:0] stage6_39;
   wire [2:0] stage7_0;
   wire [6:0] stage7_1;
   wire [0:0] stage7_2;
   wire [3:0] stage7_3;
   wire [1:0] stage7_4;
   wire [3:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [1:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [2:0] stage7_19;
   wire [6:0] stage7_20;
   wire [0:0] stage7_21;
   wire [5:0] stage7_22;
   wire [5:0] stage7_23;
   wire [3:0] stage7_24;
   wire [0:0] stage7_25;
   wire [2:0] stage7_26;
   wire [5:0] stage7_27;
   wire [5:0] stage7_28;
   wire [3:0] stage7_29;
   wire [2:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [3:0] stage7_38;
   wire [0:0] stage7_39;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [0:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [0:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [0:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc1343_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3]},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[4]},
      {stage0_2[3]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[5]},
      {stage0_2[4]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[6]},
      {stage0_2[5]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_1[7]},
      {stage0_2[6]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[8]},
      {stage0_2[7]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[9]},
      {stage0_2[8]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[10]},
      {stage0_2[9]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[11]},
      {stage0_2[10]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[12]},
      {stage0_2[11]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[13]},
      {stage0_2[12]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[14]},
      {stage0_2[13]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[15]},
      {stage0_2[14]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[16]},
      {stage0_2[15]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc117_4 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[17]},
      {stage0_2[16]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc117_4 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[18]},
      {stage0_2[17]},
      {stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc117_4 gpc16 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[19]},
      {stage0_2[18]},
      {stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[19]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[20]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[21]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[22]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[23]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[24]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[25]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[26]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[27]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[28]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[29]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[30]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[31]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[32]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[33]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[34]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[35]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[36]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[37]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[38]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[39]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[40]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[41]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[42]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[43]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[44]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[27],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[28],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[29],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[30],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[31],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[32],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[33],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[34],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[35],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[36],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[37],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[38],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[39],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[40],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[41],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[42],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[43],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[44],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[45],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[46],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[47],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[48],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[49],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[50],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[51],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[52],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[53],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[54],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[55],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[56],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[57],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[58],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[59],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[60],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[61],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[62],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[63],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[64],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[65],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[66],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437], stage0_0[438]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[67],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc1325_5 gpc84 (
      {stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_1[176], stage0_1[177]},
      {stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage0_3[27]},
      {stage1_4[68],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[0],stage1_4[69],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[1],stage1_4[70],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[2],stage1_4[71],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[3],stage1_4[72],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[4],stage1_4[73],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[5],stage1_4[74],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[6],stage1_4[75],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[7],stage1_4[76],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[8],stage1_4[77],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[9],stage1_4[78],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[10],stage1_4[79],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[11],stage1_4[80],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[12],stage1_4[81],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[13],stage1_4[82],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[14],stage1_4[83],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[15],stage1_4[84],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279]},
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage1_5[16],stage1_4[85],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285]},
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135]},
      {stage1_5[17],stage1_4[86],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291]},
      {stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141]},
      {stage1_5[18],stage1_4[87],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297]},
      {stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147]},
      {stage1_5[19],stage1_4[88],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303]},
      {stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153]},
      {stage1_5[20],stage1_4[89],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309]},
      {stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159]},
      {stage1_5[21],stage1_4[90],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315]},
      {stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165]},
      {stage1_5[22],stage1_4[91],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321]},
      {stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage1_5[23],stage1_4[92],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327]},
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177]},
      {stage1_5[24],stage1_4[93],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333]},
      {stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183]},
      {stage1_5[25],stage1_4[94],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339]},
      {stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189]},
      {stage1_5[26],stage1_4[95],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345]},
      {stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195]},
      {stage1_5[27],stage1_4[96],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351]},
      {stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage1_5[28],stage1_4[97],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357]},
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207]},
      {stage1_5[29],stage1_4[98],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363]},
      {stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213]},
      {stage1_5[30],stage1_4[99],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369]},
      {stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219]},
      {stage1_5[31],stage1_4[100],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375]},
      {stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage1_5[32],stage1_4[101],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381]},
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage1_5[33],stage1_4[102],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387]},
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage1_5[34],stage1_4[103],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393]},
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243]},
      {stage1_5[35],stage1_4[104],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399]},
      {stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249]},
      {stage1_5[36],stage1_4[105],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405]},
      {stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255]},
      {stage1_5[37],stage1_4[106],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411]},
      {stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage1_5[38],stage1_4[107],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417]},
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267]},
      {stage1_5[39],stage1_4[108],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423]},
      {stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273]},
      {stage1_5[40],stage1_4[109],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429]},
      {stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279]},
      {stage1_5[41],stage1_4[110],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435]},
      {stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage1_5[42],stage1_4[111],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441]},
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage1_5[43],stage1_4[112],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447]},
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296], stage0_3[297]},
      {stage1_5[44],stage1_4[113],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453]},
      {stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302], stage0_3[303]},
      {stage1_5[45],stage1_4[114],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459]},
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309]},
      {stage1_5[46],stage1_4[115],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465]},
      {stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage1_5[47],stage1_4[116],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471]},
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage1_5[48],stage1_4[117],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477]},
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327]},
      {stage1_5[49],stage1_4[118],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[478], stage0_1[479], stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483]},
      {stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage1_5[50],stage1_4[119],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[51],stage1_4[120],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[52],stage1_4[121],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[53],stage1_4[122],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[54],stage1_4[123],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[55],stage1_4[124],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[56],stage1_4[125],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[57],stage1_4[126],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[58],stage1_4[127],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[59],stage1_4[128],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[60],stage1_4[129],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[61],stage1_4[130],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[62],stage1_4[131],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[63],stage1_4[132],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[64],stage1_4[133],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[65],stage1_4[134],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[66],stage1_4[135],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394]},
      {stage0_3[334]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[67],stage1_4[136],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399]},
      {stage0_3[335]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[68],stage1_4[137],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage0_3[336]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[69],stage1_4[138],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409]},
      {stage0_3[337]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[70],stage1_4[139],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage0_3[338]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[71],stage1_4[140],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[126]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[21],stage1_5[72],stage1_4[141],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[127]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[22],stage1_5[73],stage1_4[142],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[128]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[23],stage1_5[74],stage1_4[143],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[129]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[24],stage1_5[75],stage1_4[144],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[130]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[25],stage1_5[76],stage1_4[145],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[131]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[26],stage1_5[77],stage1_4[146],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[132]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[27],stage1_5[78],stage1_4[147],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[133]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[28],stage1_5[79],stage1_4[148],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[134]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[29],stage1_5[80],stage1_4[149],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[135]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[30],stage1_5[81],stage1_4[150],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[136]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[31],stage1_5[82],stage1_4[151],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[137]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[32],stage1_5[83],stage1_4[152],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[138]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[33],stage1_5[84],stage1_4[153],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[139]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[34],stage1_5[85],stage1_4[154],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[140]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[35],stage1_5[86],stage1_4[155],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[414], stage0_3[415], stage0_3[416], stage0_3[417], stage0_3[418]},
      {stage0_4[141]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[36],stage1_5[87],stage1_4[156],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422], stage0_3[423]},
      {stage0_4[142]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[37],stage1_5[88],stage1_4[157],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage0_4[143]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[38],stage1_5[89],stage1_4[158],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433]},
      {stage0_4[144]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[39],stage1_5[90],stage1_4[159],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[434], stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438]},
      {stage0_4[145]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[40],stage1_5[91],stage1_4[160],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[439], stage0_3[440], stage0_3[441], stage0_3[442], stage0_3[443]},
      {stage0_4[146]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[41],stage1_5[92],stage1_4[161],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[444], stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448]},
      {stage0_4[147]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[42],stage1_5[93],stage1_4[162],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[449], stage0_3[450], stage0_3[451], stage0_3[452], stage0_3[453]},
      {stage0_4[148]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[43],stage1_5[94],stage1_4[163],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[454], stage0_3[455], stage0_3[456], stage0_3[457], stage0_3[458]},
      {stage0_4[149]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[44],stage1_5[95],stage1_4[164],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[459], stage0_3[460], stage0_3[461], stage0_3[462], stage0_3[463]},
      {stage0_4[150]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[45],stage1_5[96],stage1_4[165],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[464], stage0_3[465], stage0_3[466], stage0_3[467], stage0_3[468]},
      {stage0_4[151]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[46],stage1_5[97],stage1_4[166],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[469], stage0_3[470], stage0_3[471], stage0_3[472], stage0_3[473]},
      {stage0_4[152]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[47],stage1_5[98],stage1_4[167],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[474], stage0_3[475], stage0_3[476], stage0_3[477], stage0_3[478]},
      {stage0_4[153]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[48],stage1_5[99],stage1_4[168],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[479], stage0_3[480], stage0_3[481], stage0_3[482], stage0_3[483]},
      {stage0_4[154]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[49],stage1_5[100],stage1_4[169],stage1_3[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[29],stage1_6[50],stage1_5[101],stage1_4[170]}
   );
   gpc606_5 gpc187 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[30],stage1_6[51],stage1_5[102],stage1_4[171]}
   );
   gpc606_5 gpc188 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[31],stage1_6[52],stage1_5[103],stage1_4[172]}
   );
   gpc606_5 gpc189 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[32],stage1_6[53],stage1_5[104],stage1_4[173]}
   );
   gpc606_5 gpc190 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[33],stage1_6[54],stage1_5[105],stage1_4[174]}
   );
   gpc606_5 gpc191 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[34],stage1_6[55],stage1_5[106],stage1_4[175]}
   );
   gpc606_5 gpc192 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[35],stage1_6[56],stage1_5[107],stage1_4[176]}
   );
   gpc606_5 gpc193 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[36],stage1_6[57],stage1_5[108],stage1_4[177]}
   );
   gpc606_5 gpc194 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[37],stage1_6[58],stage1_5[109],stage1_4[178]}
   );
   gpc606_5 gpc195 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[38],stage1_6[59],stage1_5[110],stage1_4[179]}
   );
   gpc606_5 gpc196 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[39],stage1_6[60],stage1_5[111],stage1_4[180]}
   );
   gpc606_5 gpc197 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[40],stage1_6[61],stage1_5[112],stage1_4[181]}
   );
   gpc606_5 gpc198 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[41],stage1_6[62],stage1_5[113],stage1_4[182]}
   );
   gpc606_5 gpc199 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[42],stage1_6[63],stage1_5[114],stage1_4[183]}
   );
   gpc606_5 gpc200 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[43],stage1_6[64],stage1_5[115],stage1_4[184]}
   );
   gpc606_5 gpc201 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[44],stage1_6[65],stage1_5[116],stage1_4[185]}
   );
   gpc606_5 gpc202 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[45],stage1_6[66],stage1_5[117],stage1_4[186]}
   );
   gpc606_5 gpc203 (
      {stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[46],stage1_6[67],stage1_5[118],stage1_4[187]}
   );
   gpc606_5 gpc204 (
      {stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[47],stage1_6[68],stage1_5[119],stage1_4[188]}
   );
   gpc606_5 gpc205 (
      {stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[48],stage1_6[69],stage1_5[120],stage1_4[189]}
   );
   gpc606_5 gpc206 (
      {stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[49],stage1_6[70],stage1_5[121],stage1_4[190]}
   );
   gpc606_5 gpc207 (
      {stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[50],stage1_6[71],stage1_5[122],stage1_4[191]}
   );
   gpc606_5 gpc208 (
      {stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[51],stage1_6[72],stage1_5[123],stage1_4[192]}
   );
   gpc606_5 gpc209 (
      {stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[52],stage1_6[73],stage1_5[124],stage1_4[193]}
   );
   gpc606_5 gpc210 (
      {stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[53],stage1_6[74],stage1_5[125],stage1_4[194]}
   );
   gpc606_5 gpc211 (
      {stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[54],stage1_6[75],stage1_5[126],stage1_4[195]}
   );
   gpc606_5 gpc212 (
      {stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[55],stage1_6[76],stage1_5[127],stage1_4[196]}
   );
   gpc606_5 gpc213 (
      {stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[56],stage1_6[77],stage1_5[128],stage1_4[197]}
   );
   gpc606_5 gpc214 (
      {stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[57],stage1_6[78],stage1_5[129],stage1_4[198]}
   );
   gpc606_5 gpc215 (
      {stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[58],stage1_6[79],stage1_5[130],stage1_4[199]}
   );
   gpc606_5 gpc216 (
      {stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[59],stage1_6[80],stage1_5[131],stage1_4[200]}
   );
   gpc606_5 gpc217 (
      {stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[60],stage1_6[81],stage1_5[132],stage1_4[201]}
   );
   gpc606_5 gpc218 (
      {stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[61],stage1_6[82],stage1_5[133],stage1_4[202]}
   );
   gpc606_5 gpc219 (
      {stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[62],stage1_6[83],stage1_5[134],stage1_4[203]}
   );
   gpc606_5 gpc220 (
      {stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[63],stage1_6[84],stage1_5[135],stage1_4[204]}
   );
   gpc606_5 gpc221 (
      {stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[64],stage1_6[85],stage1_5[136],stage1_4[205]}
   );
   gpc606_5 gpc222 (
      {stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[65],stage1_6[86],stage1_5[137],stage1_4[206]}
   );
   gpc606_5 gpc223 (
      {stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[66],stage1_6[87],stage1_5[138],stage1_4[207]}
   );
   gpc606_5 gpc224 (
      {stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[67],stage1_6[88],stage1_5[139],stage1_4[208]}
   );
   gpc606_5 gpc225 (
      {stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[68],stage1_6[89],stage1_5[140],stage1_4[209]}
   );
   gpc606_5 gpc226 (
      {stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[69],stage1_6[90],stage1_5[141],stage1_4[210]}
   );
   gpc606_5 gpc227 (
      {stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[70],stage1_6[91],stage1_5[142],stage1_4[211]}
   );
   gpc606_5 gpc228 (
      {stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[71],stage1_6[92],stage1_5[143],stage1_4[212]}
   );
   gpc606_5 gpc229 (
      {stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[72],stage1_6[93],stage1_5[144],stage1_4[213]}
   );
   gpc606_5 gpc230 (
      {stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[73],stage1_6[94],stage1_5[145],stage1_4[214]}
   );
   gpc606_5 gpc231 (
      {stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[74],stage1_6[95],stage1_5[146],stage1_4[215]}
   );
   gpc606_5 gpc232 (
      {stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[75],stage1_6[96],stage1_5[147],stage1_4[216]}
   );
   gpc606_5 gpc233 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[76],stage1_6[97],stage1_5[148],stage1_4[217]}
   );
   gpc606_5 gpc234 (
      {stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[77],stage1_6[98],stage1_5[149],stage1_4[218]}
   );
   gpc606_5 gpc235 (
      {stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[78],stage1_6[99],stage1_5[150],stage1_4[219]}
   );
   gpc606_5 gpc236 (
      {stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[79],stage1_6[100],stage1_5[151],stage1_4[220]}
   );
   gpc606_5 gpc237 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[80],stage1_6[101],stage1_5[152],stage1_4[221]}
   );
   gpc606_5 gpc238 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[81],stage1_6[102],stage1_5[153],stage1_4[222]}
   );
   gpc606_5 gpc239 (
      {stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[82],stage1_6[103],stage1_5[154],stage1_4[223]}
   );
   gpc606_5 gpc240 (
      {stage0_4[479], stage0_4[480], stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[83],stage1_6[104],stage1_5[155],stage1_4[224]}
   );
   gpc606_5 gpc241 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[84],stage1_6[105],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[85],stage1_6[106],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[86],stage1_6[107],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[87],stage1_6[108],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[88],stage1_6[109],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[89],stage1_6[110],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[90],stage1_6[111],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[91],stage1_6[112],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[92],stage1_6[113],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[93],stage1_6[114],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[94],stage1_6[115],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[95],stage1_6[116],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[96],stage1_6[117],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[97],stage1_6[118],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[98],stage1_6[119],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[99],stage1_6[120],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[100],stage1_6[121],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[101],stage1_6[122],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[102],stage1_6[123],stage1_5[174]}
   );
   gpc606_5 gpc260 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[103],stage1_6[124],stage1_5[175]}
   );
   gpc606_5 gpc261 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[104],stage1_6[125],stage1_5[176]}
   );
   gpc606_5 gpc262 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[105],stage1_6[126],stage1_5[177]}
   );
   gpc606_5 gpc263 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[106],stage1_6[127],stage1_5[178]}
   );
   gpc606_5 gpc264 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[107],stage1_6[128],stage1_5[179]}
   );
   gpc606_5 gpc265 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[108],stage1_6[129],stage1_5[180]}
   );
   gpc606_5 gpc266 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[109],stage1_6[130],stage1_5[181]}
   );
   gpc606_5 gpc267 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[110],stage1_6[131],stage1_5[182]}
   );
   gpc606_5 gpc268 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[111],stage1_6[132],stage1_5[183]}
   );
   gpc606_5 gpc269 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[112],stage1_6[133],stage1_5[184]}
   );
   gpc606_5 gpc270 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[113],stage1_6[134],stage1_5[185]}
   );
   gpc606_5 gpc271 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[114],stage1_6[135],stage1_5[186]}
   );
   gpc606_5 gpc272 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[115],stage1_6[136],stage1_5[187]}
   );
   gpc606_5 gpc273 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[116],stage1_6[137],stage1_5[188]}
   );
   gpc606_5 gpc274 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[117],stage1_6[138],stage1_5[189]}
   );
   gpc606_5 gpc275 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[118],stage1_6[139],stage1_5[190]}
   );
   gpc606_5 gpc276 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[119],stage1_6[140],stage1_5[191]}
   );
   gpc606_5 gpc277 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[120],stage1_6[141],stage1_5[192]}
   );
   gpc606_5 gpc278 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[121],stage1_6[142],stage1_5[193]}
   );
   gpc606_5 gpc279 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[122],stage1_6[143],stage1_5[194]}
   );
   gpc606_5 gpc280 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[123],stage1_6[144],stage1_5[195]}
   );
   gpc606_5 gpc281 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[124],stage1_6[145],stage1_5[196]}
   );
   gpc606_5 gpc282 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[125],stage1_6[146],stage1_5[197]}
   );
   gpc606_5 gpc283 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[126],stage1_6[147],stage1_5[198]}
   );
   gpc606_5 gpc284 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[127],stage1_6[148],stage1_5[199]}
   );
   gpc606_5 gpc285 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[128],stage1_6[149],stage1_5[200]}
   );
   gpc606_5 gpc286 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[129],stage1_6[150],stage1_5[201]}
   );
   gpc606_5 gpc287 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[130],stage1_6[151],stage1_5[202]}
   );
   gpc606_5 gpc288 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[131],stage1_6[152],stage1_5[203]}
   );
   gpc606_5 gpc289 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[132],stage1_6[153],stage1_5[204]}
   );
   gpc606_5 gpc290 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[133],stage1_6[154],stage1_5[205]}
   );
   gpc615_5 gpc291 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[105],stage1_7[134],stage1_6[155]}
   );
   gpc615_5 gpc292 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[106],stage1_7[135],stage1_6[156]}
   );
   gpc615_5 gpc293 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[107],stage1_7[136],stage1_6[157]}
   );
   gpc615_5 gpc294 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[108],stage1_7[137],stage1_6[158]}
   );
   gpc615_5 gpc295 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[109],stage1_7[138],stage1_6[159]}
   );
   gpc615_5 gpc296 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[110],stage1_7[139],stage1_6[160]}
   );
   gpc615_5 gpc297 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[111],stage1_7[140],stage1_6[161]}
   );
   gpc615_5 gpc298 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[112],stage1_7[141],stage1_6[162]}
   );
   gpc615_5 gpc299 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[113],stage1_7[142],stage1_6[163]}
   );
   gpc615_5 gpc300 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[114],stage1_7[143],stage1_6[164]}
   );
   gpc615_5 gpc301 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[115],stage1_7[144],stage1_6[165]}
   );
   gpc615_5 gpc302 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[116],stage1_7[145],stage1_6[166]}
   );
   gpc615_5 gpc303 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[117],stage1_7[146],stage1_6[167]}
   );
   gpc615_5 gpc304 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[118],stage1_7[147],stage1_6[168]}
   );
   gpc615_5 gpc305 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[119],stage1_7[148],stage1_6[169]}
   );
   gpc615_5 gpc306 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[120],stage1_7[149],stage1_6[170]}
   );
   gpc615_5 gpc307 (
      {stage0_7[316], stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320]},
      {stage0_8[96]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[16],stage1_9[66],stage1_8[121],stage1_7[150]}
   );
   gpc615_5 gpc308 (
      {stage0_7[321], stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325]},
      {stage0_8[97]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[17],stage1_9[67],stage1_8[122],stage1_7[151]}
   );
   gpc615_5 gpc309 (
      {stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330]},
      {stage0_8[98]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[18],stage1_9[68],stage1_8[123],stage1_7[152]}
   );
   gpc615_5 gpc310 (
      {stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage0_8[99]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[19],stage1_9[69],stage1_8[124],stage1_7[153]}
   );
   gpc615_5 gpc311 (
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340]},
      {stage0_8[100]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[20],stage1_9[70],stage1_8[125],stage1_7[154]}
   );
   gpc615_5 gpc312 (
      {stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345]},
      {stage0_8[101]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[21],stage1_9[71],stage1_8[126],stage1_7[155]}
   );
   gpc615_5 gpc313 (
      {stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350]},
      {stage0_8[102]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[22],stage1_9[72],stage1_8[127],stage1_7[156]}
   );
   gpc615_5 gpc314 (
      {stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355]},
      {stage0_8[103]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[23],stage1_9[73],stage1_8[128],stage1_7[157]}
   );
   gpc615_5 gpc315 (
      {stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360]},
      {stage0_8[104]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[24],stage1_9[74],stage1_8[129],stage1_7[158]}
   );
   gpc615_5 gpc316 (
      {stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage0_8[105]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[25],stage1_9[75],stage1_8[130],stage1_7[159]}
   );
   gpc615_5 gpc317 (
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_8[106]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[26],stage1_9[76],stage1_8[131],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375]},
      {stage0_8[107]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[27],stage1_9[77],stage1_8[132],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380]},
      {stage0_8[108]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[28],stage1_9[78],stage1_8[133],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385]},
      {stage0_8[109]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[29],stage1_9[79],stage1_8[134],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390]},
      {stage0_8[110]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[30],stage1_9[80],stage1_8[135],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage0_8[111]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[31],stage1_9[81],stage1_8[136],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_8[112]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[32],stage1_9[82],stage1_8[137],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405]},
      {stage0_8[113]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[33],stage1_9[83],stage1_8[138],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410]},
      {stage0_8[114]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[34],stage1_9[84],stage1_8[139],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415]},
      {stage0_8[115]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[35],stage1_9[85],stage1_8[140],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420]},
      {stage0_8[116]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[36],stage1_9[86],stage1_8[141],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage0_8[117]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[37],stage1_9[87],stage1_8[142],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_8[118]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[38],stage1_9[88],stage1_8[143],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435]},
      {stage0_8[119]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[39],stage1_9[89],stage1_8[144],stage1_7[173]}
   );
   gpc606_5 gpc331 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[24],stage1_10[40],stage1_9[90],stage1_8[145]}
   );
   gpc606_5 gpc332 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[25],stage1_10[41],stage1_9[91],stage1_8[146]}
   );
   gpc606_5 gpc333 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[26],stage1_10[42],stage1_9[92],stage1_8[147]}
   );
   gpc606_5 gpc334 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[27],stage1_10[43],stage1_9[93],stage1_8[148]}
   );
   gpc606_5 gpc335 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[28],stage1_10[44],stage1_9[94],stage1_8[149]}
   );
   gpc606_5 gpc336 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[29],stage1_10[45],stage1_9[95],stage1_8[150]}
   );
   gpc606_5 gpc337 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[30],stage1_10[46],stage1_9[96],stage1_8[151]}
   );
   gpc606_5 gpc338 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[31],stage1_10[47],stage1_9[97],stage1_8[152]}
   );
   gpc606_5 gpc339 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[32],stage1_10[48],stage1_9[98],stage1_8[153]}
   );
   gpc606_5 gpc340 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[33],stage1_10[49],stage1_9[99],stage1_8[154]}
   );
   gpc606_5 gpc341 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[34],stage1_10[50],stage1_9[100],stage1_8[155]}
   );
   gpc606_5 gpc342 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[35],stage1_10[51],stage1_9[101],stage1_8[156]}
   );
   gpc606_5 gpc343 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[36],stage1_10[52],stage1_9[102],stage1_8[157]}
   );
   gpc606_5 gpc344 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[37],stage1_10[53],stage1_9[103],stage1_8[158]}
   );
   gpc606_5 gpc345 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[38],stage1_10[54],stage1_9[104],stage1_8[159]}
   );
   gpc606_5 gpc346 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[39],stage1_10[55],stage1_9[105],stage1_8[160]}
   );
   gpc606_5 gpc347 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[40],stage1_10[56],stage1_9[106],stage1_8[161]}
   );
   gpc606_5 gpc348 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[41],stage1_10[57],stage1_9[107],stage1_8[162]}
   );
   gpc606_5 gpc349 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[42],stage1_10[58],stage1_9[108],stage1_8[163]}
   );
   gpc606_5 gpc350 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[43],stage1_10[59],stage1_9[109],stage1_8[164]}
   );
   gpc606_5 gpc351 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[44],stage1_10[60],stage1_9[110],stage1_8[165]}
   );
   gpc606_5 gpc352 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[45],stage1_10[61],stage1_9[111],stage1_8[166]}
   );
   gpc606_5 gpc353 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[46],stage1_10[62],stage1_9[112],stage1_8[167]}
   );
   gpc606_5 gpc354 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[47],stage1_10[63],stage1_9[113],stage1_8[168]}
   );
   gpc606_5 gpc355 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[48],stage1_10[64],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc356 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[49],stage1_10[65],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc357 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[50],stage1_10[66],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc358 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[51],stage1_10[67],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc359 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[52],stage1_10[68],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc360 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[53],stage1_10[69],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc361 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[54],stage1_10[70],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc362 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[55],stage1_10[71],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc363 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[56],stage1_10[72],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc364 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[57],stage1_10[73],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc365 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[58],stage1_10[74],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc366 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[59],stage1_10[75],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc367 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[60],stage1_10[76],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc368 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[61],stage1_10[77],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc369 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[62],stage1_10[78],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc370 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[63],stage1_10[79],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc371 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[64],stage1_10[80],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc372 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[65],stage1_10[81],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc373 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[66],stage1_10[82],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc374 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[67],stage1_10[83],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc375 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[68],stage1_10[84],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc376 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[69],stage1_10[85],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc377 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[70],stage1_10[86],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc378 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[71],stage1_10[87],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc379 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[72],stage1_10[88],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc380 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[73],stage1_10[89],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc381 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[74],stage1_10[90],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc382 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[75],stage1_10[91],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc383 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[76],stage1_10[92],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc384 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[77],stage1_10[93],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc385 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[78],stage1_10[94],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc386 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[79],stage1_10[95],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc387 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[80],stage1_10[96],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc388 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[81],stage1_10[97],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc389 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[82],stage1_10[98],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc390 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[83],stage1_10[99],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc391 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[84],stage1_10[100],stage1_9[150],stage1_8[205]}
   );
   gpc117_4 gpc392 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[366]},
      {stage0_11[0]},
      {stage1_12[61],stage1_11[85],stage1_10[101],stage1_9[151]}
   );
   gpc117_4 gpc393 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156], stage0_9[157]},
      {stage0_10[367]},
      {stage0_11[1]},
      {stage1_12[62],stage1_11[86],stage1_10[102],stage1_9[152]}
   );
   gpc117_4 gpc394 (
      {stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164]},
      {stage0_10[368]},
      {stage0_11[2]},
      {stage1_12[63],stage1_11[87],stage1_10[103],stage1_9[153]}
   );
   gpc117_4 gpc395 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171]},
      {stage0_10[369]},
      {stage0_11[3]},
      {stage1_12[64],stage1_11[88],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177]},
      {stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9]},
      {stage1_13[0],stage1_12[65],stage1_11[89],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183]},
      {stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15]},
      {stage1_13[1],stage1_12[66],stage1_11[90],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189]},
      {stage0_11[16], stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21]},
      {stage1_13[2],stage1_12[67],stage1_11[91],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage1_13[3],stage1_12[68],stage1_11[92],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201]},
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33]},
      {stage1_13[4],stage1_12[69],stage1_11[93],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207]},
      {stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39]},
      {stage1_13[5],stage1_12[70],stage1_11[94],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213]},
      {stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45]},
      {stage1_13[6],stage1_12[71],stage1_11[95],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_11[46], stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51]},
      {stage1_13[7],stage1_12[72],stage1_11[96],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_11[52], stage0_11[53], stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57]},
      {stage1_13[8],stage1_12[73],stage1_11[97],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231]},
      {stage0_11[58], stage0_11[59], stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63]},
      {stage1_13[9],stage1_12[74],stage1_11[98],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237]},
      {stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69]},
      {stage1_13[10],stage1_12[75],stage1_11[99],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243]},
      {stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75]},
      {stage1_13[11],stage1_12[76],stage1_11[100],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249]},
      {stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81]},
      {stage1_13[12],stage1_12[77],stage1_11[101],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87]},
      {stage1_13[13],stage1_12[78],stage1_11[102],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261]},
      {stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93]},
      {stage1_13[14],stage1_12[79],stage1_11[103],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267]},
      {stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99]},
      {stage1_13[15],stage1_12[80],stage1_11[104],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273]},
      {stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105]},
      {stage1_13[16],stage1_12[81],stage1_11[105],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279]},
      {stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111]},
      {stage1_13[17],stage1_12[82],stage1_11[106],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117]},
      {stage1_13[18],stage1_12[83],stage1_11[107],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291]},
      {stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123]},
      {stage1_13[19],stage1_12[84],stage1_11[108],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297]},
      {stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage1_13[20],stage1_12[85],stage1_11[109],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303]},
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135]},
      {stage1_13[21],stage1_12[86],stage1_11[110],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309]},
      {stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141]},
      {stage1_13[22],stage1_12[87],stage1_11[111],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_11[142], stage0_11[143], stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147]},
      {stage1_13[23],stage1_12[88],stage1_11[112],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321]},
      {stage0_11[148], stage0_11[149], stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153]},
      {stage1_13[24],stage1_12[89],stage1_11[113],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327]},
      {stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage1_13[25],stage1_12[90],stage1_11[114],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333]},
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165]},
      {stage1_13[26],stage1_12[91],stage1_11[115],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339]},
      {stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171]},
      {stage1_13[27],stage1_12[92],stage1_11[116],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_11[172], stage0_11[173], stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177]},
      {stage1_13[28],stage1_12[93],stage1_11[117],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351]},
      {stage0_11[178], stage0_11[179], stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183]},
      {stage1_13[29],stage1_12[94],stage1_11[118],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357]},
      {stage0_11[184], stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage1_13[30],stage1_12[95],stage1_11[119],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363]},
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195]},
      {stage1_13[31],stage1_12[96],stage1_11[120],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369]},
      {stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201]},
      {stage1_13[32],stage1_12[97],stage1_11[121],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_11[202], stage0_11[203], stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207]},
      {stage1_13[33],stage1_12[98],stage1_11[122],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381]},
      {stage0_11[208], stage0_11[209], stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213]},
      {stage1_13[34],stage1_12[99],stage1_11[123],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387]},
      {stage0_11[214], stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage1_13[35],stage1_12[100],stage1_11[124],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393]},
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225]},
      {stage1_13[36],stage1_12[101],stage1_11[125],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399]},
      {stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231]},
      {stage1_13[37],stage1_12[102],stage1_11[126],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_11[232], stage0_11[233], stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237]},
      {stage1_13[38],stage1_12[103],stage1_11[127],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411]},
      {stage0_11[238], stage0_11[239], stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243]},
      {stage1_13[39],stage1_12[104],stage1_11[128],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417]},
      {stage0_11[244], stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage1_13[40],stage1_12[105],stage1_11[129],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc437 (
      {stage0_9[418], stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255]},
      {stage1_13[41],stage1_12[106],stage1_11[130],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc438 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429]},
      {stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261]},
      {stage1_13[42],stage1_12[107],stage1_11[131],stage1_10[147],stage1_9[197]}
   );
   gpc606_5 gpc439 (
      {stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_11[262], stage0_11[263], stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267]},
      {stage1_13[43],stage1_12[108],stage1_11[132],stage1_10[148],stage1_9[198]}
   );
   gpc606_5 gpc440 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441]},
      {stage0_11[268], stage0_11[269], stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273]},
      {stage1_13[44],stage1_12[109],stage1_11[133],stage1_10[149],stage1_9[199]}
   );
   gpc606_5 gpc441 (
      {stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447]},
      {stage0_11[274], stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage1_13[45],stage1_12[110],stage1_11[134],stage1_10[150],stage1_9[200]}
   );
   gpc606_5 gpc442 (
      {stage0_9[448], stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285]},
      {stage1_13[46],stage1_12[111],stage1_11[135],stage1_10[151],stage1_9[201]}
   );
   gpc606_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459]},
      {stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291]},
      {stage1_13[47],stage1_12[112],stage1_11[136],stage1_10[152],stage1_9[202]}
   );
   gpc606_5 gpc444 (
      {stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_11[292], stage0_11[293], stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297]},
      {stage1_13[48],stage1_12[113],stage1_11[137],stage1_10[153],stage1_9[203]}
   );
   gpc606_5 gpc445 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471]},
      {stage0_11[298], stage0_11[299], stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303]},
      {stage1_13[49],stage1_12[114],stage1_11[138],stage1_10[154],stage1_9[204]}
   );
   gpc606_5 gpc446 (
      {stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477]},
      {stage0_11[304], stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage1_13[50],stage1_12[115],stage1_11[139],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc447 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374]},
      {stage0_11[310]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[51],stage1_12[116],stage1_11[140],stage1_10[156]}
   );
   gpc615_5 gpc448 (
      {stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379]},
      {stage0_11[311]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[52],stage1_12[117],stage1_11[141],stage1_10[157]}
   );
   gpc615_5 gpc449 (
      {stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383], stage0_10[384]},
      {stage0_11[312]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[53],stage1_12[118],stage1_11[142],stage1_10[158]}
   );
   gpc615_5 gpc450 (
      {stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage0_11[313]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[54],stage1_12[119],stage1_11[143],stage1_10[159]}
   );
   gpc615_5 gpc451 (
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394]},
      {stage0_11[314]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[55],stage1_12[120],stage1_11[144],stage1_10[160]}
   );
   gpc615_5 gpc452 (
      {stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_11[315]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[56],stage1_12[121],stage1_11[145],stage1_10[161]}
   );
   gpc615_5 gpc453 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404]},
      {stage0_11[316]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[57],stage1_12[122],stage1_11[146],stage1_10[162]}
   );
   gpc615_5 gpc454 (
      {stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409]},
      {stage0_11[317]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[58],stage1_12[123],stage1_11[147],stage1_10[163]}
   );
   gpc615_5 gpc455 (
      {stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413], stage0_10[414]},
      {stage0_11[318]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[59],stage1_12[124],stage1_11[148],stage1_10[164]}
   );
   gpc615_5 gpc456 (
      {stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage0_11[319]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[60],stage1_12[125],stage1_11[149],stage1_10[165]}
   );
   gpc615_5 gpc457 (
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424]},
      {stage0_11[320]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[61],stage1_12[126],stage1_11[150],stage1_10[166]}
   );
   gpc615_5 gpc458 (
      {stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429]},
      {stage0_11[321]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[62],stage1_12[127],stage1_11[151],stage1_10[167]}
   );
   gpc615_5 gpc459 (
      {stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433], stage0_10[434]},
      {stage0_11[322]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[63],stage1_12[128],stage1_11[152],stage1_10[168]}
   );
   gpc615_5 gpc460 (
      {stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438], stage0_10[439]},
      {stage0_11[323]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[64],stage1_12[129],stage1_11[153],stage1_10[169]}
   );
   gpc615_5 gpc461 (
      {stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443], stage0_10[444]},
      {stage0_11[324]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[65],stage1_12[130],stage1_11[154],stage1_10[170]}
   );
   gpc615_5 gpc462 (
      {stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage0_11[325]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[66],stage1_12[131],stage1_11[155],stage1_10[171]}
   );
   gpc615_5 gpc463 (
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454]},
      {stage0_11[326]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[67],stage1_12[132],stage1_11[156],stage1_10[172]}
   );
   gpc615_5 gpc464 (
      {stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459]},
      {stage0_11[327]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[68],stage1_12[133],stage1_11[157],stage1_10[173]}
   );
   gpc615_5 gpc465 (
      {stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463], stage0_10[464]},
      {stage0_11[328]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[69],stage1_12[134],stage1_11[158],stage1_10[174]}
   );
   gpc615_5 gpc466 (
      {stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468], stage0_10[469]},
      {stage0_11[329]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[70],stage1_12[135],stage1_11[159],stage1_10[175]}
   );
   gpc615_5 gpc467 (
      {stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473], stage0_10[474]},
      {stage0_11[330]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[71],stage1_12[136],stage1_11[160],stage1_10[176]}
   );
   gpc615_5 gpc468 (
      {stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage0_12[126]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[21],stage1_13[72],stage1_12[137],stage1_11[161]}
   );
   gpc615_5 gpc469 (
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340]},
      {stage0_12[127]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[22],stage1_13[73],stage1_12[138],stage1_11[162]}
   );
   gpc615_5 gpc470 (
      {stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345]},
      {stage0_12[128]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[23],stage1_13[74],stage1_12[139],stage1_11[163]}
   );
   gpc615_5 gpc471 (
      {stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350]},
      {stage0_12[129]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[24],stage1_13[75],stage1_12[140],stage1_11[164]}
   );
   gpc615_5 gpc472 (
      {stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355]},
      {stage0_12[130]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[25],stage1_13[76],stage1_12[141],stage1_11[165]}
   );
   gpc615_5 gpc473 (
      {stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360]},
      {stage0_12[131]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[26],stage1_13[77],stage1_12[142],stage1_11[166]}
   );
   gpc615_5 gpc474 (
      {stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage0_12[132]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[27],stage1_13[78],stage1_12[143],stage1_11[167]}
   );
   gpc615_5 gpc475 (
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370]},
      {stage0_12[133]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[28],stage1_13[79],stage1_12[144],stage1_11[168]}
   );
   gpc615_5 gpc476 (
      {stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375]},
      {stage0_12[134]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[29],stage1_13[80],stage1_12[145],stage1_11[169]}
   );
   gpc615_5 gpc477 (
      {stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379], stage0_11[380]},
      {stage0_12[135]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[30],stage1_13[81],stage1_12[146],stage1_11[170]}
   );
   gpc615_5 gpc478 (
      {stage0_11[381], stage0_11[382], stage0_11[383], stage0_11[384], stage0_11[385]},
      {stage0_12[136]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[31],stage1_13[82],stage1_12[147],stage1_11[171]}
   );
   gpc615_5 gpc479 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[137]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[32],stage1_13[83],stage1_12[148],stage1_11[172]}
   );
   gpc615_5 gpc480 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[138]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[33],stage1_13[84],stage1_12[149],stage1_11[173]}
   );
   gpc615_5 gpc481 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[139]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[34],stage1_13[85],stage1_12[150],stage1_11[174]}
   );
   gpc615_5 gpc482 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[140]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[35],stage1_13[86],stage1_12[151],stage1_11[175]}
   );
   gpc615_5 gpc483 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[141]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[36],stage1_13[87],stage1_12[152],stage1_11[176]}
   );
   gpc615_5 gpc484 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[142]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[37],stage1_13[88],stage1_12[153],stage1_11[177]}
   );
   gpc615_5 gpc485 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[143]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[38],stage1_13[89],stage1_12[154],stage1_11[178]}
   );
   gpc615_5 gpc486 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[144]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[39],stage1_13[90],stage1_12[155],stage1_11[179]}
   );
   gpc615_5 gpc487 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[145]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[40],stage1_13[91],stage1_12[156],stage1_11[180]}
   );
   gpc615_5 gpc488 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[146]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[41],stage1_13[92],stage1_12[157],stage1_11[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[147]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[42],stage1_13[93],stage1_12[158],stage1_11[182]}
   );
   gpc615_5 gpc490 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[148]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[43],stage1_13[94],stage1_12[159],stage1_11[183]}
   );
   gpc615_5 gpc491 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[149]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[44],stage1_13[95],stage1_12[160],stage1_11[184]}
   );
   gpc606_5 gpc492 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[24],stage1_14[45],stage1_13[96],stage1_12[161]}
   );
   gpc606_5 gpc493 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[25],stage1_14[46],stage1_13[97],stage1_12[162]}
   );
   gpc606_5 gpc494 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[26],stage1_14[47],stage1_13[98],stage1_12[163]}
   );
   gpc606_5 gpc495 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[27],stage1_14[48],stage1_13[99],stage1_12[164]}
   );
   gpc606_5 gpc496 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[28],stage1_14[49],stage1_13[100],stage1_12[165]}
   );
   gpc606_5 gpc497 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[29],stage1_14[50],stage1_13[101],stage1_12[166]}
   );
   gpc606_5 gpc498 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[30],stage1_14[51],stage1_13[102],stage1_12[167]}
   );
   gpc606_5 gpc499 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[31],stage1_14[52],stage1_13[103],stage1_12[168]}
   );
   gpc606_5 gpc500 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[32],stage1_14[53],stage1_13[104],stage1_12[169]}
   );
   gpc606_5 gpc501 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[33],stage1_14[54],stage1_13[105],stage1_12[170]}
   );
   gpc606_5 gpc502 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[34],stage1_14[55],stage1_13[106],stage1_12[171]}
   );
   gpc606_5 gpc503 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[35],stage1_14[56],stage1_13[107],stage1_12[172]}
   );
   gpc606_5 gpc504 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[36],stage1_14[57],stage1_13[108],stage1_12[173]}
   );
   gpc606_5 gpc505 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[37],stage1_14[58],stage1_13[109],stage1_12[174]}
   );
   gpc606_5 gpc506 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[38],stage1_14[59],stage1_13[110],stage1_12[175]}
   );
   gpc606_5 gpc507 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[39],stage1_14[60],stage1_13[111],stage1_12[176]}
   );
   gpc606_5 gpc508 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[40],stage1_14[61],stage1_13[112],stage1_12[177]}
   );
   gpc606_5 gpc509 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[41],stage1_14[62],stage1_13[113],stage1_12[178]}
   );
   gpc606_5 gpc510 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[42],stage1_14[63],stage1_13[114],stage1_12[179]}
   );
   gpc606_5 gpc511 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[43],stage1_14[64],stage1_13[115],stage1_12[180]}
   );
   gpc606_5 gpc512 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[44],stage1_14[65],stage1_13[116],stage1_12[181]}
   );
   gpc606_5 gpc513 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[45],stage1_14[66],stage1_13[117],stage1_12[182]}
   );
   gpc606_5 gpc514 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[46],stage1_14[67],stage1_13[118],stage1_12[183]}
   );
   gpc606_5 gpc515 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[47],stage1_14[68],stage1_13[119],stage1_12[184]}
   );
   gpc606_5 gpc516 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[48],stage1_14[69],stage1_13[120],stage1_12[185]}
   );
   gpc606_5 gpc517 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[49],stage1_14[70],stage1_13[121],stage1_12[186]}
   );
   gpc606_5 gpc518 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[50],stage1_14[71],stage1_13[122],stage1_12[187]}
   );
   gpc606_5 gpc519 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[51],stage1_14[72],stage1_13[123],stage1_12[188]}
   );
   gpc606_5 gpc520 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[52],stage1_14[73],stage1_13[124],stage1_12[189]}
   );
   gpc606_5 gpc521 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[53],stage1_14[74],stage1_13[125],stage1_12[190]}
   );
   gpc606_5 gpc522 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[54],stage1_14[75],stage1_13[126],stage1_12[191]}
   );
   gpc606_5 gpc523 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[55],stage1_14[76],stage1_13[127],stage1_12[192]}
   );
   gpc606_5 gpc524 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[56],stage1_14[77],stage1_13[128],stage1_12[193]}
   );
   gpc606_5 gpc525 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[57],stage1_14[78],stage1_13[129],stage1_12[194]}
   );
   gpc606_5 gpc526 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[58],stage1_14[79],stage1_13[130],stage1_12[195]}
   );
   gpc606_5 gpc527 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[59],stage1_14[80],stage1_13[131],stage1_12[196]}
   );
   gpc606_5 gpc528 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[60],stage1_14[81],stage1_13[132],stage1_12[197]}
   );
   gpc606_5 gpc529 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[61],stage1_14[82],stage1_13[133],stage1_12[198]}
   );
   gpc606_5 gpc530 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[62],stage1_14[83],stage1_13[134],stage1_12[199]}
   );
   gpc606_5 gpc531 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[63],stage1_14[84],stage1_13[135],stage1_12[200]}
   );
   gpc606_5 gpc532 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[64],stage1_14[85],stage1_13[136],stage1_12[201]}
   );
   gpc606_5 gpc533 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[65],stage1_14[86],stage1_13[137],stage1_12[202]}
   );
   gpc606_5 gpc534 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[66],stage1_14[87],stage1_13[138],stage1_12[203]}
   );
   gpc606_5 gpc535 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[43],stage1_15[67],stage1_14[88],stage1_13[139]}
   );
   gpc606_5 gpc536 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[44],stage1_15[68],stage1_14[89],stage1_13[140]}
   );
   gpc606_5 gpc537 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[45],stage1_15[69],stage1_14[90],stage1_13[141]}
   );
   gpc606_5 gpc538 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[46],stage1_15[70],stage1_14[91],stage1_13[142]}
   );
   gpc606_5 gpc539 (
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[47],stage1_15[71],stage1_14[92],stage1_13[143]}
   );
   gpc606_5 gpc540 (
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[48],stage1_15[72],stage1_14[93],stage1_13[144]}
   );
   gpc606_5 gpc541 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[49],stage1_15[73],stage1_14[94],stage1_13[145]}
   );
   gpc606_5 gpc542 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[50],stage1_15[74],stage1_14[95],stage1_13[146]}
   );
   gpc606_5 gpc543 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[51],stage1_15[75],stage1_14[96],stage1_13[147]}
   );
   gpc606_5 gpc544 (
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[52],stage1_15[76],stage1_14[97],stage1_13[148]}
   );
   gpc606_5 gpc545 (
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[53],stage1_15[77],stage1_14[98],stage1_13[149]}
   );
   gpc606_5 gpc546 (
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[54],stage1_15[78],stage1_14[99],stage1_13[150]}
   );
   gpc606_5 gpc547 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[55],stage1_15[79],stage1_14[100],stage1_13[151]}
   );
   gpc606_5 gpc548 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[56],stage1_15[80],stage1_14[101],stage1_13[152]}
   );
   gpc606_5 gpc549 (
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[57],stage1_15[81],stage1_14[102],stage1_13[153]}
   );
   gpc606_5 gpc550 (
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[58],stage1_15[82],stage1_14[103],stage1_13[154]}
   );
   gpc606_5 gpc551 (
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[59],stage1_15[83],stage1_14[104],stage1_13[155]}
   );
   gpc606_5 gpc552 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[60],stage1_15[84],stage1_14[105],stage1_13[156]}
   );
   gpc606_5 gpc553 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[61],stage1_15[85],stage1_14[106],stage1_13[157]}
   );
   gpc606_5 gpc554 (
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[62],stage1_15[86],stage1_14[107],stage1_13[158]}
   );
   gpc606_5 gpc555 (
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[63],stage1_15[87],stage1_14[108],stage1_13[159]}
   );
   gpc606_5 gpc556 (
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[64],stage1_15[88],stage1_14[109],stage1_13[160]}
   );
   gpc606_5 gpc557 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[65],stage1_15[89],stage1_14[110],stage1_13[161]}
   );
   gpc606_5 gpc558 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[66],stage1_15[90],stage1_14[111],stage1_13[162]}
   );
   gpc606_5 gpc559 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[67],stage1_15[91],stage1_14[112],stage1_13[163]}
   );
   gpc606_5 gpc560 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[68],stage1_15[92],stage1_14[113],stage1_13[164]}
   );
   gpc606_5 gpc561 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[69],stage1_15[93],stage1_14[114],stage1_13[165]}
   );
   gpc606_5 gpc562 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[70],stage1_15[94],stage1_14[115],stage1_13[166]}
   );
   gpc606_5 gpc563 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[71],stage1_15[95],stage1_14[116],stage1_13[167]}
   );
   gpc606_5 gpc564 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[72],stage1_15[96],stage1_14[117],stage1_13[168]}
   );
   gpc606_5 gpc565 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[73],stage1_15[97],stage1_14[118],stage1_13[169]}
   );
   gpc606_5 gpc566 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[74],stage1_15[98],stage1_14[119],stage1_13[170]}
   );
   gpc606_5 gpc567 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[75],stage1_15[99],stage1_14[120],stage1_13[171]}
   );
   gpc606_5 gpc568 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[76],stage1_15[100],stage1_14[121],stage1_13[172]}
   );
   gpc606_5 gpc569 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[77],stage1_15[101],stage1_14[122],stage1_13[173]}
   );
   gpc606_5 gpc570 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[78],stage1_15[102],stage1_14[123],stage1_13[174]}
   );
   gpc606_5 gpc571 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[79],stage1_15[103],stage1_14[124],stage1_13[175]}
   );
   gpc606_5 gpc572 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[80],stage1_15[104],stage1_14[125],stage1_13[176]}
   );
   gpc606_5 gpc573 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[81],stage1_15[105],stage1_14[126],stage1_13[177]}
   );
   gpc606_5 gpc574 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[82],stage1_15[106],stage1_14[127],stage1_13[178]}
   );
   gpc606_5 gpc575 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[83],stage1_15[107],stage1_14[128],stage1_13[179]}
   );
   gpc606_5 gpc576 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[84],stage1_15[108],stage1_14[129],stage1_13[180]}
   );
   gpc606_5 gpc577 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[85],stage1_15[109],stage1_14[130],stage1_13[181]}
   );
   gpc606_5 gpc578 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[86],stage1_15[110],stage1_14[131],stage1_13[182]}
   );
   gpc606_5 gpc579 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[87],stage1_15[111],stage1_14[132],stage1_13[183]}
   );
   gpc606_5 gpc580 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[88],stage1_15[112],stage1_14[133],stage1_13[184]}
   );
   gpc606_5 gpc581 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[89],stage1_15[113],stage1_14[134],stage1_13[185]}
   );
   gpc606_5 gpc582 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[90],stage1_15[114],stage1_14[135],stage1_13[186]}
   );
   gpc606_5 gpc583 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[91],stage1_15[115],stage1_14[136],stage1_13[187]}
   );
   gpc606_5 gpc584 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[92],stage1_15[116],stage1_14[137],stage1_13[188]}
   );
   gpc606_5 gpc585 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[93],stage1_15[117],stage1_14[138],stage1_13[189]}
   );
   gpc606_5 gpc586 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[94],stage1_15[118],stage1_14[139],stage1_13[190]}
   );
   gpc615_5 gpc587 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[258]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[95],stage1_15[119],stage1_14[140],stage1_13[191]}
   );
   gpc615_5 gpc588 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[259]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[96],stage1_15[120],stage1_14[141],stage1_13[192]}
   );
   gpc615_5 gpc589 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[260]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[97],stage1_15[121],stage1_14[142],stage1_13[193]}
   );
   gpc615_5 gpc590 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[261]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[98],stage1_15[122],stage1_14[143],stage1_13[194]}
   );
   gpc606_5 gpc591 (
      {stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[56],stage1_16[99],stage1_15[123],stage1_14[144]}
   );
   gpc606_5 gpc592 (
      {stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[57],stage1_16[100],stage1_15[124],stage1_14[145]}
   );
   gpc606_5 gpc593 (
      {stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[58],stage1_16[101],stage1_15[125],stage1_14[146]}
   );
   gpc606_5 gpc594 (
      {stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[59],stage1_16[102],stage1_15[126],stage1_14[147]}
   );
   gpc606_5 gpc595 (
      {stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[60],stage1_16[103],stage1_15[127],stage1_14[148]}
   );
   gpc606_5 gpc596 (
      {stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[61],stage1_16[104],stage1_15[128],stage1_14[149]}
   );
   gpc606_5 gpc597 (
      {stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[62],stage1_16[105],stage1_15[129],stage1_14[150]}
   );
   gpc615_5 gpc598 (
      {stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307], stage0_14[308]},
      {stage0_15[336]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[63],stage1_16[106],stage1_15[130],stage1_14[151]}
   );
   gpc615_5 gpc599 (
      {stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage0_15[337]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[64],stage1_16[107],stage1_15[131],stage1_14[152]}
   );
   gpc615_5 gpc600 (
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318]},
      {stage0_15[338]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[65],stage1_16[108],stage1_15[132],stage1_14[153]}
   );
   gpc615_5 gpc601 (
      {stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_15[339]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[66],stage1_16[109],stage1_15[133],stage1_14[154]}
   );
   gpc615_5 gpc602 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328]},
      {stage0_15[340]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[67],stage1_16[110],stage1_15[134],stage1_14[155]}
   );
   gpc615_5 gpc603 (
      {stage0_14[329], stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333]},
      {stage0_15[341]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[68],stage1_16[111],stage1_15[135],stage1_14[156]}
   );
   gpc615_5 gpc604 (
      {stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337], stage0_14[338]},
      {stage0_15[342]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[69],stage1_16[112],stage1_15[136],stage1_14[157]}
   );
   gpc615_5 gpc605 (
      {stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage0_15[343]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[70],stage1_16[113],stage1_15[137],stage1_14[158]}
   );
   gpc615_5 gpc606 (
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348]},
      {stage0_15[344]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[71],stage1_16[114],stage1_15[138],stage1_14[159]}
   );
   gpc615_5 gpc607 (
      {stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_16[96]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[16],stage1_17[72],stage1_16[115],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354]},
      {stage0_16[97]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[17],stage1_17[73],stage1_16[116],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage0_16[98]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[18],stage1_17[74],stage1_16[117],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364]},
      {stage0_16[99]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[19],stage1_17[75],stage1_16[118],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369]},
      {stage0_16[100]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[20],stage1_17[76],stage1_16[119],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374]},
      {stage0_16[101]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[21],stage1_17[77],stage1_16[120],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379]},
      {stage0_16[102]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[22],stage1_17[78],stage1_16[121],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384]},
      {stage0_16[103]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[23],stage1_17[79],stage1_16[122],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage0_16[104]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[24],stage1_17[80],stage1_16[123],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394]},
      {stage0_16[105]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[25],stage1_17[81],stage1_16[124],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399]},
      {stage0_16[106]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[26],stage1_17[82],stage1_16[125],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404]},
      {stage0_16[107]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[27],stage1_17[83],stage1_16[126],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409]},
      {stage0_16[108]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[28],stage1_17[84],stage1_16[127],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414]},
      {stage0_16[109]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[29],stage1_17[85],stage1_16[128],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage0_16[110]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[30],stage1_17[86],stage1_16[129],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424]},
      {stage0_16[111]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[31],stage1_17[87],stage1_16[130],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429]},
      {stage0_16[112]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[32],stage1_17[88],stage1_16[131],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434]},
      {stage0_16[113]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[33],stage1_17[89],stage1_16[132],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439]},
      {stage0_16[114]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[34],stage1_17[90],stage1_16[133],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444]},
      {stage0_16[115]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[35],stage1_17[91],stage1_16[134],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage0_16[116]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[36],stage1_17[92],stage1_16[135],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454]},
      {stage0_16[117]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[37],stage1_17[93],stage1_16[136],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459]},
      {stage0_16[118]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[38],stage1_17[94],stage1_16[137],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463], stage0_15[464]},
      {stage0_16[119]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[39],stage1_17[95],stage1_16[138],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468], stage0_15[469]},
      {stage0_16[120]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[40],stage1_17[96],stage1_16[139],stage1_15[163]}
   );
   gpc615_5 gpc632 (
      {stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473], stage0_15[474]},
      {stage0_16[121]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[41],stage1_17[97],stage1_16[140],stage1_15[164]}
   );
   gpc615_5 gpc633 (
      {stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage0_16[122]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[42],stage1_17[98],stage1_16[141],stage1_15[165]}
   );
   gpc606_5 gpc634 (
      {stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127], stage0_16[128]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[27],stage1_18[43],stage1_17[99],stage1_16[142]}
   );
   gpc606_5 gpc635 (
      {stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133], stage0_16[134]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[28],stage1_18[44],stage1_17[100],stage1_16[143]}
   );
   gpc606_5 gpc636 (
      {stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139], stage0_16[140]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[29],stage1_18[45],stage1_17[101],stage1_16[144]}
   );
   gpc606_5 gpc637 (
      {stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145], stage0_16[146]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[30],stage1_18[46],stage1_17[102],stage1_16[145]}
   );
   gpc606_5 gpc638 (
      {stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[31],stage1_18[47],stage1_17[103],stage1_16[146]}
   );
   gpc606_5 gpc639 (
      {stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[32],stage1_18[48],stage1_17[104],stage1_16[147]}
   );
   gpc606_5 gpc640 (
      {stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[33],stage1_18[49],stage1_17[105],stage1_16[148]}
   );
   gpc606_5 gpc641 (
      {stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[34],stage1_18[50],stage1_17[106],stage1_16[149]}
   );
   gpc606_5 gpc642 (
      {stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[35],stage1_18[51],stage1_17[107],stage1_16[150]}
   );
   gpc606_5 gpc643 (
      {stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[36],stage1_18[52],stage1_17[108],stage1_16[151]}
   );
   gpc606_5 gpc644 (
      {stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[37],stage1_18[53],stage1_17[109],stage1_16[152]}
   );
   gpc606_5 gpc645 (
      {stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[38],stage1_18[54],stage1_17[110],stage1_16[153]}
   );
   gpc606_5 gpc646 (
      {stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[39],stage1_18[55],stage1_17[111],stage1_16[154]}
   );
   gpc606_5 gpc647 (
      {stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[40],stage1_18[56],stage1_17[112],stage1_16[155]}
   );
   gpc606_5 gpc648 (
      {stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[41],stage1_18[57],stage1_17[113],stage1_16[156]}
   );
   gpc606_5 gpc649 (
      {stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[42],stage1_18[58],stage1_17[114],stage1_16[157]}
   );
   gpc606_5 gpc650 (
      {stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[43],stage1_18[59],stage1_17[115],stage1_16[158]}
   );
   gpc606_5 gpc651 (
      {stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[44],stage1_18[60],stage1_17[116],stage1_16[159]}
   );
   gpc606_5 gpc652 (
      {stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[45],stage1_18[61],stage1_17[117],stage1_16[160]}
   );
   gpc606_5 gpc653 (
      {stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[46],stage1_18[62],stage1_17[118],stage1_16[161]}
   );
   gpc606_5 gpc654 (
      {stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[47],stage1_18[63],stage1_17[119],stage1_16[162]}
   );
   gpc606_5 gpc655 (
      {stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[48],stage1_18[64],stage1_17[120],stage1_16[163]}
   );
   gpc606_5 gpc656 (
      {stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259], stage0_16[260]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[49],stage1_18[65],stage1_17[121],stage1_16[164]}
   );
   gpc606_5 gpc657 (
      {stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265], stage0_16[266]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[50],stage1_18[66],stage1_17[122],stage1_16[165]}
   );
   gpc606_5 gpc658 (
      {stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271], stage0_16[272]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[51],stage1_18[67],stage1_17[123],stage1_16[166]}
   );
   gpc606_5 gpc659 (
      {stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277], stage0_16[278]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[52],stage1_18[68],stage1_17[124],stage1_16[167]}
   );
   gpc606_5 gpc660 (
      {stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283], stage0_16[284]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[53],stage1_18[69],stage1_17[125],stage1_16[168]}
   );
   gpc606_5 gpc661 (
      {stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289], stage0_16[290]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[54],stage1_18[70],stage1_17[126],stage1_16[169]}
   );
   gpc606_5 gpc662 (
      {stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295], stage0_16[296]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[55],stage1_18[71],stage1_17[127],stage1_16[170]}
   );
   gpc606_5 gpc663 (
      {stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301], stage0_16[302]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[56],stage1_18[72],stage1_17[128],stage1_16[171]}
   );
   gpc606_5 gpc664 (
      {stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307], stage0_16[308]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[57],stage1_18[73],stage1_17[129],stage1_16[172]}
   );
   gpc606_5 gpc665 (
      {stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313], stage0_16[314]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[58],stage1_18[74],stage1_17[130],stage1_16[173]}
   );
   gpc606_5 gpc666 (
      {stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319], stage0_16[320]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[59],stage1_18[75],stage1_17[131],stage1_16[174]}
   );
   gpc606_5 gpc667 (
      {stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325], stage0_16[326]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[60],stage1_18[76],stage1_17[132],stage1_16[175]}
   );
   gpc606_5 gpc668 (
      {stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331], stage0_16[332]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[61],stage1_18[77],stage1_17[133],stage1_16[176]}
   );
   gpc606_5 gpc669 (
      {stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337], stage0_16[338]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[62],stage1_18[78],stage1_17[134],stage1_16[177]}
   );
   gpc606_5 gpc670 (
      {stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343], stage0_16[344]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[63],stage1_18[79],stage1_17[135],stage1_16[178]}
   );
   gpc606_5 gpc671 (
      {stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349], stage0_16[350]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[64],stage1_18[80],stage1_17[136],stage1_16[179]}
   );
   gpc606_5 gpc672 (
      {stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355], stage0_16[356]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[65],stage1_18[81],stage1_17[137],stage1_16[180]}
   );
   gpc606_5 gpc673 (
      {stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361], stage0_16[362]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[66],stage1_18[82],stage1_17[138],stage1_16[181]}
   );
   gpc606_5 gpc674 (
      {stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367], stage0_16[368]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[67],stage1_18[83],stage1_17[139],stage1_16[182]}
   );
   gpc606_5 gpc675 (
      {stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373], stage0_16[374]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[68],stage1_18[84],stage1_17[140],stage1_16[183]}
   );
   gpc606_5 gpc676 (
      {stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379], stage0_16[380]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[69],stage1_18[85],stage1_17[141],stage1_16[184]}
   );
   gpc606_5 gpc677 (
      {stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385], stage0_16[386]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[70],stage1_18[86],stage1_17[142],stage1_16[185]}
   );
   gpc606_5 gpc678 (
      {stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391], stage0_16[392]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[71],stage1_18[87],stage1_17[143],stage1_16[186]}
   );
   gpc606_5 gpc679 (
      {stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397], stage0_16[398]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[72],stage1_18[88],stage1_17[144],stage1_16[187]}
   );
   gpc606_5 gpc680 (
      {stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403], stage0_16[404]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[73],stage1_18[89],stage1_17[145],stage1_16[188]}
   );
   gpc606_5 gpc681 (
      {stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409], stage0_16[410]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[74],stage1_18[90],stage1_17[146],stage1_16[189]}
   );
   gpc606_5 gpc682 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[48],stage1_19[75],stage1_18[91],stage1_17[147]}
   );
   gpc606_5 gpc683 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[49],stage1_19[76],stage1_18[92],stage1_17[148]}
   );
   gpc606_5 gpc684 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[50],stage1_19[77],stage1_18[93],stage1_17[149]}
   );
   gpc606_5 gpc685 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[51],stage1_19[78],stage1_18[94],stage1_17[150]}
   );
   gpc606_5 gpc686 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[52],stage1_19[79],stage1_18[95],stage1_17[151]}
   );
   gpc606_5 gpc687 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[53],stage1_19[80],stage1_18[96],stage1_17[152]}
   );
   gpc606_5 gpc688 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[54],stage1_19[81],stage1_18[97],stage1_17[153]}
   );
   gpc606_5 gpc689 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[55],stage1_19[82],stage1_18[98],stage1_17[154]}
   );
   gpc606_5 gpc690 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[56],stage1_19[83],stage1_18[99],stage1_17[155]}
   );
   gpc606_5 gpc691 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[57],stage1_19[84],stage1_18[100],stage1_17[156]}
   );
   gpc606_5 gpc692 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[58],stage1_19[85],stage1_18[101],stage1_17[157]}
   );
   gpc606_5 gpc693 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[59],stage1_19[86],stage1_18[102],stage1_17[158]}
   );
   gpc606_5 gpc694 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[60],stage1_19[87],stage1_18[103],stage1_17[159]}
   );
   gpc606_5 gpc695 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[61],stage1_19[88],stage1_18[104],stage1_17[160]}
   );
   gpc606_5 gpc696 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[62],stage1_19[89],stage1_18[105],stage1_17[161]}
   );
   gpc606_5 gpc697 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[63],stage1_19[90],stage1_18[106],stage1_17[162]}
   );
   gpc606_5 gpc698 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[64],stage1_19[91],stage1_18[107],stage1_17[163]}
   );
   gpc606_5 gpc699 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[65],stage1_19[92],stage1_18[108],stage1_17[164]}
   );
   gpc606_5 gpc700 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[66],stage1_19[93],stage1_18[109],stage1_17[165]}
   );
   gpc606_5 gpc701 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[67],stage1_19[94],stage1_18[110],stage1_17[166]}
   );
   gpc606_5 gpc702 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[68],stage1_19[95],stage1_18[111],stage1_17[167]}
   );
   gpc606_5 gpc703 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[69],stage1_19[96],stage1_18[112],stage1_17[168]}
   );
   gpc606_5 gpc704 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[70],stage1_19[97],stage1_18[113],stage1_17[169]}
   );
   gpc606_5 gpc705 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[71],stage1_19[98],stage1_18[114],stage1_17[170]}
   );
   gpc606_5 gpc706 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[72],stage1_19[99],stage1_18[115],stage1_17[171]}
   );
   gpc606_5 gpc707 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[73],stage1_19[100],stage1_18[116],stage1_17[172]}
   );
   gpc606_5 gpc708 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[74],stage1_19[101],stage1_18[117],stage1_17[173]}
   );
   gpc606_5 gpc709 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[75],stage1_19[102],stage1_18[118],stage1_17[174]}
   );
   gpc606_5 gpc710 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[76],stage1_19[103],stage1_18[119],stage1_17[175]}
   );
   gpc606_5 gpc711 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[77],stage1_19[104],stage1_18[120],stage1_17[176]}
   );
   gpc606_5 gpc712 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[78],stage1_19[105],stage1_18[121],stage1_17[177]}
   );
   gpc606_5 gpc713 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[79],stage1_19[106],stage1_18[122],stage1_17[178]}
   );
   gpc606_5 gpc714 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[80],stage1_19[107],stage1_18[123],stage1_17[179]}
   );
   gpc606_5 gpc715 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[81],stage1_19[108],stage1_18[124],stage1_17[180]}
   );
   gpc606_5 gpc716 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[82],stage1_19[109],stage1_18[125],stage1_17[181]}
   );
   gpc606_5 gpc717 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[83],stage1_19[110],stage1_18[126],stage1_17[182]}
   );
   gpc606_5 gpc718 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[84],stage1_19[111],stage1_18[127],stage1_17[183]}
   );
   gpc606_5 gpc719 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[85],stage1_19[112],stage1_18[128],stage1_17[184]}
   );
   gpc606_5 gpc720 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[86],stage1_19[113],stage1_18[129],stage1_17[185]}
   );
   gpc606_5 gpc721 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[87],stage1_19[114],stage1_18[130],stage1_17[186]}
   );
   gpc606_5 gpc722 (
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[40],stage1_20[88],stage1_19[115],stage1_18[131]}
   );
   gpc606_5 gpc723 (
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[41],stage1_20[89],stage1_19[116],stage1_18[132]}
   );
   gpc606_5 gpc724 (
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[42],stage1_20[90],stage1_19[117],stage1_18[133]}
   );
   gpc606_5 gpc725 (
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[43],stage1_20[91],stage1_19[118],stage1_18[134]}
   );
   gpc615_5 gpc726 (
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316]},
      {stage0_19[240]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[44],stage1_20[92],stage1_19[119],stage1_18[135]}
   );
   gpc615_5 gpc727 (
      {stage0_18[317], stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321]},
      {stage0_19[241]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[45],stage1_20[93],stage1_19[120],stage1_18[136]}
   );
   gpc615_5 gpc728 (
      {stage0_18[322], stage0_18[323], stage0_18[324], stage0_18[325], stage0_18[326]},
      {stage0_19[242]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[46],stage1_20[94],stage1_19[121],stage1_18[137]}
   );
   gpc615_5 gpc729 (
      {stage0_18[327], stage0_18[328], stage0_18[329], stage0_18[330], stage0_18[331]},
      {stage0_19[243]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[47],stage1_20[95],stage1_19[122],stage1_18[138]}
   );
   gpc615_5 gpc730 (
      {stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335], stage0_18[336]},
      {stage0_19[244]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[48],stage1_20[96],stage1_19[123],stage1_18[139]}
   );
   gpc615_5 gpc731 (
      {stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage0_19[245]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[49],stage1_20[97],stage1_19[124],stage1_18[140]}
   );
   gpc615_5 gpc732 (
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346]},
      {stage0_19[246]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[50],stage1_20[98],stage1_19[125],stage1_18[141]}
   );
   gpc615_5 gpc733 (
      {stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351]},
      {stage0_19[247]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[51],stage1_20[99],stage1_19[126],stage1_18[142]}
   );
   gpc615_5 gpc734 (
      {stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355], stage0_18[356]},
      {stage0_19[248]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[52],stage1_20[100],stage1_19[127],stage1_18[143]}
   );
   gpc615_5 gpc735 (
      {stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360], stage0_18[361]},
      {stage0_19[249]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[53],stage1_20[101],stage1_19[128],stage1_18[144]}
   );
   gpc615_5 gpc736 (
      {stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365], stage0_18[366]},
      {stage0_19[250]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[54],stage1_20[102],stage1_19[129],stage1_18[145]}
   );
   gpc615_5 gpc737 (
      {stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage0_19[251]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[55],stage1_20[103],stage1_19[130],stage1_18[146]}
   );
   gpc615_5 gpc738 (
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376]},
      {stage0_19[252]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[56],stage1_20[104],stage1_19[131],stage1_18[147]}
   );
   gpc615_5 gpc739 (
      {stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381]},
      {stage0_19[253]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[57],stage1_20[105],stage1_19[132],stage1_18[148]}
   );
   gpc615_5 gpc740 (
      {stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385], stage0_18[386]},
      {stage0_19[254]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[58],stage1_20[106],stage1_19[133],stage1_18[149]}
   );
   gpc615_5 gpc741 (
      {stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390], stage0_18[391]},
      {stage0_19[255]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[59],stage1_20[107],stage1_19[134],stage1_18[150]}
   );
   gpc615_5 gpc742 (
      {stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395], stage0_18[396]},
      {stage0_19[256]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[60],stage1_20[108],stage1_19[135],stage1_18[151]}
   );
   gpc615_5 gpc743 (
      {stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage0_19[257]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[61],stage1_20[109],stage1_19[136],stage1_18[152]}
   );
   gpc615_5 gpc744 (
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406]},
      {stage0_19[258]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[62],stage1_20[110],stage1_19[137],stage1_18[153]}
   );
   gpc615_5 gpc745 (
      {stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411]},
      {stage0_19[259]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[63],stage1_20[111],stage1_19[138],stage1_18[154]}
   );
   gpc615_5 gpc746 (
      {stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415], stage0_18[416]},
      {stage0_19[260]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[64],stage1_20[112],stage1_19[139],stage1_18[155]}
   );
   gpc615_5 gpc747 (
      {stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420], stage0_18[421]},
      {stage0_19[261]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[65],stage1_20[113],stage1_19[140],stage1_18[156]}
   );
   gpc615_5 gpc748 (
      {stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425], stage0_18[426]},
      {stage0_19[262]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[66],stage1_20[114],stage1_19[141],stage1_18[157]}
   );
   gpc615_5 gpc749 (
      {stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430], stage0_18[431]},
      {stage0_19[263]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[67],stage1_20[115],stage1_19[142],stage1_18[158]}
   );
   gpc615_5 gpc750 (
      {stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435], stage0_18[436]},
      {stage0_19[264]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[68],stage1_20[116],stage1_19[143],stage1_18[159]}
   );
   gpc615_5 gpc751 (
      {stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440], stage0_18[441]},
      {stage0_19[265]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[69],stage1_20[117],stage1_19[144],stage1_18[160]}
   );
   gpc615_5 gpc752 (
      {stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445], stage0_18[446]},
      {stage0_19[266]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[70],stage1_20[118],stage1_19[145],stage1_18[161]}
   );
   gpc606_5 gpc753 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271], stage0_19[272]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[31],stage1_21[71],stage1_20[119],stage1_19[146]}
   );
   gpc606_5 gpc754 (
      {stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276], stage0_19[277], stage0_19[278]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[32],stage1_21[72],stage1_20[120],stage1_19[147]}
   );
   gpc606_5 gpc755 (
      {stage0_19[279], stage0_19[280], stage0_19[281], stage0_19[282], stage0_19[283], stage0_19[284]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[33],stage1_21[73],stage1_20[121],stage1_19[148]}
   );
   gpc606_5 gpc756 (
      {stage0_19[285], stage0_19[286], stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[34],stage1_21[74],stage1_20[122],stage1_19[149]}
   );
   gpc606_5 gpc757 (
      {stage0_19[291], stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[35],stage1_21[75],stage1_20[123],stage1_19[150]}
   );
   gpc615_5 gpc758 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[186]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[36],stage1_21[76],stage1_20[124],stage1_19[151]}
   );
   gpc615_5 gpc759 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[187]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[37],stage1_21[77],stage1_20[125],stage1_19[152]}
   );
   gpc615_5 gpc760 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[188]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[38],stage1_21[78],stage1_20[126],stage1_19[153]}
   );
   gpc615_5 gpc761 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[189]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[39],stage1_21[79],stage1_20[127],stage1_19[154]}
   );
   gpc615_5 gpc762 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[190]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[40],stage1_21[80],stage1_20[128],stage1_19[155]}
   );
   gpc615_5 gpc763 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[191]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[41],stage1_21[81],stage1_20[129],stage1_19[156]}
   );
   gpc615_5 gpc764 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[192]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[42],stage1_21[82],stage1_20[130],stage1_19[157]}
   );
   gpc615_5 gpc765 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[193]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[43],stage1_21[83],stage1_20[131],stage1_19[158]}
   );
   gpc615_5 gpc766 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[194]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[44],stage1_21[84],stage1_20[132],stage1_19[159]}
   );
   gpc615_5 gpc767 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[195]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[45],stage1_21[85],stage1_20[133],stage1_19[160]}
   );
   gpc606_5 gpc768 (
      {stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[15],stage1_22[46],stage1_21[86],stage1_20[134]}
   );
   gpc606_5 gpc769 (
      {stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[16],stage1_22[47],stage1_21[87],stage1_20[135]}
   );
   gpc606_5 gpc770 (
      {stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[17],stage1_22[48],stage1_21[88],stage1_20[136]}
   );
   gpc606_5 gpc771 (
      {stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[18],stage1_22[49],stage1_21[89],stage1_20[137]}
   );
   gpc606_5 gpc772 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[19],stage1_22[50],stage1_21[90],stage1_20[138]}
   );
   gpc606_5 gpc773 (
      {stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[20],stage1_22[51],stage1_21[91],stage1_20[139]}
   );
   gpc606_5 gpc774 (
      {stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[21],stage1_22[52],stage1_21[92],stage1_20[140]}
   );
   gpc606_5 gpc775 (
      {stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[22],stage1_22[53],stage1_21[93],stage1_20[141]}
   );
   gpc606_5 gpc776 (
      {stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[23],stage1_22[54],stage1_21[94],stage1_20[142]}
   );
   gpc606_5 gpc777 (
      {stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[24],stage1_22[55],stage1_21[95],stage1_20[143]}
   );
   gpc606_5 gpc778 (
      {stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[25],stage1_22[56],stage1_21[96],stage1_20[144]}
   );
   gpc606_5 gpc779 (
      {stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[26],stage1_22[57],stage1_21[97],stage1_20[145]}
   );
   gpc606_5 gpc780 (
      {stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[27],stage1_22[58],stage1_21[98],stage1_20[146]}
   );
   gpc606_5 gpc781 (
      {stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[28],stage1_22[59],stage1_21[99],stage1_20[147]}
   );
   gpc606_5 gpc782 (
      {stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[29],stage1_22[60],stage1_21[100],stage1_20[148]}
   );
   gpc606_5 gpc783 (
      {stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[30],stage1_22[61],stage1_21[101],stage1_20[149]}
   );
   gpc606_5 gpc784 (
      {stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[31],stage1_22[62],stage1_21[102],stage1_20[150]}
   );
   gpc606_5 gpc785 (
      {stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[32],stage1_22[63],stage1_21[103],stage1_20[151]}
   );
   gpc606_5 gpc786 (
      {stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[33],stage1_22[64],stage1_21[104],stage1_20[152]}
   );
   gpc606_5 gpc787 (
      {stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[34],stage1_22[65],stage1_21[105],stage1_20[153]}
   );
   gpc606_5 gpc788 (
      {stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[35],stage1_22[66],stage1_21[106],stage1_20[154]}
   );
   gpc606_5 gpc789 (
      {stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[36],stage1_22[67],stage1_21[107],stage1_20[155]}
   );
   gpc606_5 gpc790 (
      {stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[37],stage1_22[68],stage1_21[108],stage1_20[156]}
   );
   gpc606_5 gpc791 (
      {stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[38],stage1_22[69],stage1_21[109],stage1_20[157]}
   );
   gpc606_5 gpc792 (
      {stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[39],stage1_22[70],stage1_21[110],stage1_20[158]}
   );
   gpc606_5 gpc793 (
      {stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[40],stage1_22[71],stage1_21[111],stage1_20[159]}
   );
   gpc606_5 gpc794 (
      {stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[41],stage1_22[72],stage1_21[112],stage1_20[160]}
   );
   gpc606_5 gpc795 (
      {stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[42],stage1_22[73],stage1_21[113],stage1_20[161]}
   );
   gpc606_5 gpc796 (
      {stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[43],stage1_22[74],stage1_21[114],stage1_20[162]}
   );
   gpc606_5 gpc797 (
      {stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[44],stage1_22[75],stage1_21[115],stage1_20[163]}
   );
   gpc606_5 gpc798 (
      {stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[45],stage1_22[76],stage1_21[116],stage1_20[164]}
   );
   gpc606_5 gpc799 (
      {stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[46],stage1_22[77],stage1_21[117],stage1_20[165]}
   );
   gpc606_5 gpc800 (
      {stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[47],stage1_22[78],stage1_21[118],stage1_20[166]}
   );
   gpc606_5 gpc801 (
      {stage0_20[394], stage0_20[395], stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[48],stage1_22[79],stage1_21[119],stage1_20[167]}
   );
   gpc606_5 gpc802 (
      {stage0_20[400], stage0_20[401], stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[49],stage1_22[80],stage1_21[120],stage1_20[168]}
   );
   gpc606_5 gpc803 (
      {stage0_20[406], stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[50],stage1_22[81],stage1_21[121],stage1_20[169]}
   );
   gpc606_5 gpc804 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[51],stage1_22[82],stage1_21[122],stage1_20[170]}
   );
   gpc606_5 gpc805 (
      {stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[52],stage1_22[83],stage1_21[123],stage1_20[171]}
   );
   gpc606_5 gpc806 (
      {stage0_20[424], stage0_20[425], stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[53],stage1_22[84],stage1_21[124],stage1_20[172]}
   );
   gpc606_5 gpc807 (
      {stage0_20[430], stage0_20[431], stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[54],stage1_22[85],stage1_21[125],stage1_20[173]}
   );
   gpc606_5 gpc808 (
      {stage0_20[436], stage0_20[437], stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[55],stage1_22[86],stage1_21[126],stage1_20[174]}
   );
   gpc606_5 gpc809 (
      {stage0_20[442], stage0_20[443], stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[56],stage1_22[87],stage1_21[127],stage1_20[175]}
   );
   gpc606_5 gpc810 (
      {stage0_20[448], stage0_20[449], stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[57],stage1_22[88],stage1_21[128],stage1_20[176]}
   );
   gpc606_5 gpc811 (
      {stage0_20[454], stage0_20[455], stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[58],stage1_22[89],stage1_21[129],stage1_20[177]}
   );
   gpc606_5 gpc812 (
      {stage0_20[460], stage0_20[461], stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[59],stage1_22[90],stage1_21[130],stage1_20[178]}
   );
   gpc606_5 gpc813 (
      {stage0_20[466], stage0_20[467], stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[60],stage1_22[91],stage1_21[131],stage1_20[179]}
   );
   gpc606_5 gpc814 (
      {stage0_20[472], stage0_20[473], stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[61],stage1_22[92],stage1_21[132],stage1_20[180]}
   );
   gpc606_5 gpc815 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[47],stage1_23[62],stage1_22[93],stage1_21[133]}
   );
   gpc606_5 gpc816 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[48],stage1_23[63],stage1_22[94],stage1_21[134]}
   );
   gpc606_5 gpc817 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[49],stage1_23[64],stage1_22[95],stage1_21[135]}
   );
   gpc606_5 gpc818 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[50],stage1_23[65],stage1_22[96],stage1_21[136]}
   );
   gpc606_5 gpc819 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[51],stage1_23[66],stage1_22[97],stage1_21[137]}
   );
   gpc606_5 gpc820 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[52],stage1_23[67],stage1_22[98],stage1_21[138]}
   );
   gpc606_5 gpc821 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[53],stage1_23[68],stage1_22[99],stage1_21[139]}
   );
   gpc606_5 gpc822 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[54],stage1_23[69],stage1_22[100],stage1_21[140]}
   );
   gpc606_5 gpc823 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[55],stage1_23[70],stage1_22[101],stage1_21[141]}
   );
   gpc606_5 gpc824 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[56],stage1_23[71],stage1_22[102],stage1_21[142]}
   );
   gpc606_5 gpc825 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[57],stage1_23[72],stage1_22[103],stage1_21[143]}
   );
   gpc606_5 gpc826 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[58],stage1_23[73],stage1_22[104],stage1_21[144]}
   );
   gpc606_5 gpc827 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[59],stage1_23[74],stage1_22[105],stage1_21[145]}
   );
   gpc606_5 gpc828 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[60],stage1_23[75],stage1_22[106],stage1_21[146]}
   );
   gpc606_5 gpc829 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[61],stage1_23[76],stage1_22[107],stage1_21[147]}
   );
   gpc606_5 gpc830 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[62],stage1_23[77],stage1_22[108],stage1_21[148]}
   );
   gpc606_5 gpc831 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[63],stage1_23[78],stage1_22[109],stage1_21[149]}
   );
   gpc606_5 gpc832 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[64],stage1_23[79],stage1_22[110],stage1_21[150]}
   );
   gpc606_5 gpc833 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[65],stage1_23[80],stage1_22[111],stage1_21[151]}
   );
   gpc606_5 gpc834 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[66],stage1_23[81],stage1_22[112],stage1_21[152]}
   );
   gpc606_5 gpc835 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[67],stage1_23[82],stage1_22[113],stage1_21[153]}
   );
   gpc606_5 gpc836 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[68],stage1_23[83],stage1_22[114],stage1_21[154]}
   );
   gpc606_5 gpc837 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[69],stage1_23[84],stage1_22[115],stage1_21[155]}
   );
   gpc606_5 gpc838 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[70],stage1_23[85],stage1_22[116],stage1_21[156]}
   );
   gpc606_5 gpc839 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[71],stage1_23[86],stage1_22[117],stage1_21[157]}
   );
   gpc606_5 gpc840 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[72],stage1_23[87],stage1_22[118],stage1_21[158]}
   );
   gpc606_5 gpc841 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[73],stage1_23[88],stage1_22[119],stage1_21[159]}
   );
   gpc606_5 gpc842 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[74],stage1_23[89],stage1_22[120],stage1_21[160]}
   );
   gpc606_5 gpc843 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[75],stage1_23[90],stage1_22[121],stage1_21[161]}
   );
   gpc606_5 gpc844 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[76],stage1_23[91],stage1_22[122],stage1_21[162]}
   );
   gpc606_5 gpc845 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[77],stage1_23[92],stage1_22[123],stage1_21[163]}
   );
   gpc606_5 gpc846 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[78],stage1_23[93],stage1_22[124],stage1_21[164]}
   );
   gpc606_5 gpc847 (
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[79],stage1_23[94],stage1_22[125],stage1_21[165]}
   );
   gpc606_5 gpc848 (
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[80],stage1_23[95],stage1_22[126],stage1_21[166]}
   );
   gpc606_5 gpc849 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[81],stage1_23[96],stage1_22[127],stage1_21[167]}
   );
   gpc606_5 gpc850 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[82],stage1_23[97],stage1_22[128],stage1_21[168]}
   );
   gpc606_5 gpc851 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[83],stage1_23[98],stage1_22[129],stage1_21[169]}
   );
   gpc606_5 gpc852 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[84],stage1_23[99],stage1_22[130],stage1_21[170]}
   );
   gpc606_5 gpc853 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[85],stage1_23[100],stage1_22[131],stage1_21[171]}
   );
   gpc606_5 gpc854 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[86],stage1_23[101],stage1_22[132],stage1_21[172]}
   );
   gpc606_5 gpc855 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[87],stage1_23[102],stage1_22[133],stage1_21[173]}
   );
   gpc606_5 gpc856 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[88],stage1_23[103],stage1_22[134],stage1_21[174]}
   );
   gpc606_5 gpc857 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[89],stage1_23[104],stage1_22[135],stage1_21[175]}
   );
   gpc606_5 gpc858 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[90],stage1_23[105],stage1_22[136],stage1_21[176]}
   );
   gpc606_5 gpc859 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[91],stage1_23[106],stage1_22[137],stage1_21[177]}
   );
   gpc606_5 gpc860 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[92],stage1_23[107],stage1_22[138],stage1_21[178]}
   );
   gpc606_5 gpc861 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[93],stage1_23[108],stage1_22[139],stage1_21[179]}
   );
   gpc606_5 gpc862 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[94],stage1_23[109],stage1_22[140],stage1_21[180]}
   );
   gpc606_5 gpc863 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[95],stage1_23[110],stage1_22[141],stage1_21[181]}
   );
   gpc606_5 gpc864 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[96],stage1_23[111],stage1_22[142],stage1_21[182]}
   );
   gpc606_5 gpc865 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[97],stage1_23[112],stage1_22[143],stage1_21[183]}
   );
   gpc606_5 gpc866 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[98],stage1_23[113],stage1_22[144],stage1_21[184]}
   );
   gpc606_5 gpc867 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[99],stage1_23[114],stage1_22[145],stage1_21[185]}
   );
   gpc606_5 gpc868 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[100],stage1_23[115],stage1_22[146],stage1_21[186]}
   );
   gpc606_5 gpc869 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[101],stage1_23[116],stage1_22[147],stage1_21[187]}
   );
   gpc606_5 gpc870 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[102],stage1_23[117],stage1_22[148],stage1_21[188]}
   );
   gpc606_5 gpc871 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[103],stage1_23[118],stage1_22[149],stage1_21[189]}
   );
   gpc606_5 gpc872 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[104],stage1_23[119],stage1_22[150],stage1_21[190]}
   );
   gpc606_5 gpc873 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[105],stage1_23[120],stage1_22[151],stage1_21[191]}
   );
   gpc606_5 gpc874 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[106],stage1_23[121],stage1_22[152],stage1_21[192]}
   );
   gpc606_5 gpc875 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[107],stage1_23[122],stage1_22[153],stage1_21[193]}
   );
   gpc606_5 gpc876 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[108],stage1_23[123],stage1_22[154],stage1_21[194]}
   );
   gpc606_5 gpc877 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[109],stage1_23[124],stage1_22[155],stage1_21[195]}
   );
   gpc606_5 gpc878 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[110],stage1_23[125],stage1_22[156],stage1_21[196]}
   );
   gpc606_5 gpc879 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[111],stage1_23[126],stage1_22[157],stage1_21[197]}
   );
   gpc606_5 gpc880 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[112],stage1_23[127],stage1_22[158],stage1_21[198]}
   );
   gpc615_5 gpc881 (
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286]},
      {stage0_23[396]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[66],stage1_24[113],stage1_23[128],stage1_22[159]}
   );
   gpc615_5 gpc882 (
      {stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291]},
      {stage0_23[397]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[67],stage1_24[114],stage1_23[129],stage1_22[160]}
   );
   gpc615_5 gpc883 (
      {stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage0_23[398]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[68],stage1_24[115],stage1_23[130],stage1_22[161]}
   );
   gpc615_5 gpc884 (
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301]},
      {stage0_23[399]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[69],stage1_24[116],stage1_23[131],stage1_22[162]}
   );
   gpc615_5 gpc885 (
      {stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306]},
      {stage0_23[400]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[70],stage1_24[117],stage1_23[132],stage1_22[163]}
   );
   gpc615_5 gpc886 (
      {stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage0_23[401]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[71],stage1_24[118],stage1_23[133],stage1_22[164]}
   );
   gpc615_5 gpc887 (
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316]},
      {stage0_23[402]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[72],stage1_24[119],stage1_23[134],stage1_22[165]}
   );
   gpc615_5 gpc888 (
      {stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321]},
      {stage0_23[403]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[73],stage1_24[120],stage1_23[135],stage1_22[166]}
   );
   gpc615_5 gpc889 (
      {stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage0_23[404]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[74],stage1_24[121],stage1_23[136],stage1_22[167]}
   );
   gpc615_5 gpc890 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331]},
      {stage0_23[405]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[75],stage1_24[122],stage1_23[137],stage1_22[168]}
   );
   gpc615_5 gpc891 (
      {stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336]},
      {stage0_23[406]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[76],stage1_24[123],stage1_23[138],stage1_22[169]}
   );
   gpc615_5 gpc892 (
      {stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage0_23[407]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[77],stage1_24[124],stage1_23[139],stage1_22[170]}
   );
   gpc615_5 gpc893 (
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346]},
      {stage0_23[408]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[78],stage1_24[125],stage1_23[140],stage1_22[171]}
   );
   gpc615_5 gpc894 (
      {stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351]},
      {stage0_23[409]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[79],stage1_24[126],stage1_23[141],stage1_22[172]}
   );
   gpc615_5 gpc895 (
      {stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_23[410]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[80],stage1_24[127],stage1_23[142],stage1_22[173]}
   );
   gpc615_5 gpc896 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361]},
      {stage0_23[411]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[81],stage1_24[128],stage1_23[143],stage1_22[174]}
   );
   gpc615_5 gpc897 (
      {stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366]},
      {stage0_23[412]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[82],stage1_24[129],stage1_23[144],stage1_22[175]}
   );
   gpc615_5 gpc898 (
      {stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage0_23[413]},
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage1_26[17],stage1_25[83],stage1_24[130],stage1_23[145],stage1_22[176]}
   );
   gpc615_5 gpc899 (
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376]},
      {stage0_23[414]},
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage1_26[18],stage1_25[84],stage1_24[131],stage1_23[146],stage1_22[177]}
   );
   gpc615_5 gpc900 (
      {stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381]},
      {stage0_23[415]},
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage1_26[19],stage1_25[85],stage1_24[132],stage1_23[147],stage1_22[178]}
   );
   gpc615_5 gpc901 (
      {stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_23[416]},
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage1_26[20],stage1_25[86],stage1_24[133],stage1_23[148],stage1_22[179]}
   );
   gpc615_5 gpc902 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[417]},
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage1_26[21],stage1_25[87],stage1_24[134],stage1_23[149],stage1_22[180]}
   );
   gpc615_5 gpc903 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[418]},
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage1_26[22],stage1_25[88],stage1_24[135],stage1_23[150],stage1_22[181]}
   );
   gpc615_5 gpc904 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[419]},
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage1_26[23],stage1_25[89],stage1_24[136],stage1_23[151],stage1_22[182]}
   );
   gpc615_5 gpc905 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[420]},
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage1_26[24],stage1_25[90],stage1_24[137],stage1_23[152],stage1_22[183]}
   );
   gpc615_5 gpc906 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[421]},
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage1_26[25],stage1_25[91],stage1_24[138],stage1_23[153],stage1_22[184]}
   );
   gpc615_5 gpc907 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[422]},
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage1_26[26],stage1_25[92],stage1_24[139],stage1_23[154],stage1_22[185]}
   );
   gpc615_5 gpc908 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[423]},
      {stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167]},
      {stage1_26[27],stage1_25[93],stage1_24[140],stage1_23[155],stage1_22[186]}
   );
   gpc615_5 gpc909 (
      {stage0_23[424], stage0_23[425], stage0_23[426], stage0_23[427], stage0_23[428]},
      {stage0_24[168]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[28],stage1_25[94],stage1_24[141],stage1_23[156]}
   );
   gpc615_5 gpc910 (
      {stage0_23[429], stage0_23[430], stage0_23[431], stage0_23[432], stage0_23[433]},
      {stage0_24[169]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[29],stage1_25[95],stage1_24[142],stage1_23[157]}
   );
   gpc615_5 gpc911 (
      {stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437], stage0_23[438]},
      {stage0_24[170]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[30],stage1_25[96],stage1_24[143],stage1_23[158]}
   );
   gpc615_5 gpc912 (
      {stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage0_24[171]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[31],stage1_25[97],stage1_24[144],stage1_23[159]}
   );
   gpc615_5 gpc913 (
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448]},
      {stage0_24[172]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[32],stage1_25[98],stage1_24[145],stage1_23[160]}
   );
   gpc615_5 gpc914 (
      {stage0_23[449], stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453]},
      {stage0_24[173]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[33],stage1_25[99],stage1_24[146],stage1_23[161]}
   );
   gpc615_5 gpc915 (
      {stage0_23[454], stage0_23[455], stage0_23[456], stage0_23[457], stage0_23[458]},
      {stage0_24[174]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[34],stage1_25[100],stage1_24[147],stage1_23[162]}
   );
   gpc615_5 gpc916 (
      {stage0_23[459], stage0_23[460], stage0_23[461], stage0_23[462], stage0_23[463]},
      {stage0_24[175]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[35],stage1_25[101],stage1_24[148],stage1_23[163]}
   );
   gpc615_5 gpc917 (
      {stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467], stage0_23[468]},
      {stage0_24[176]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[36],stage1_25[102],stage1_24[149],stage1_23[164]}
   );
   gpc615_5 gpc918 (
      {stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage0_24[177]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[37],stage1_25[103],stage1_24[150],stage1_23[165]}
   );
   gpc606_5 gpc919 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[38],stage1_25[104],stage1_24[151]}
   );
   gpc606_5 gpc920 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[39],stage1_25[105],stage1_24[152]}
   );
   gpc606_5 gpc921 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[40],stage1_25[106],stage1_24[153]}
   );
   gpc615_5 gpc922 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200]},
      {stage0_25[60]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[41],stage1_25[107],stage1_24[154]}
   );
   gpc615_5 gpc923 (
      {stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205]},
      {stage0_25[61]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[42],stage1_25[108],stage1_24[155]}
   );
   gpc615_5 gpc924 (
      {stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_25[62]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[43],stage1_25[109],stage1_24[156]}
   );
   gpc615_5 gpc925 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215]},
      {stage0_25[63]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[44],stage1_25[110],stage1_24[157]}
   );
   gpc615_5 gpc926 (
      {stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_25[64]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[45],stage1_25[111],stage1_24[158]}
   );
   gpc615_5 gpc927 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_25[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[46],stage1_25[112],stage1_24[159]}
   );
   gpc615_5 gpc928 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230]},
      {stage0_25[66]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[47],stage1_25[113],stage1_24[160]}
   );
   gpc615_5 gpc929 (
      {stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235]},
      {stage0_25[67]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[48],stage1_25[114],stage1_24[161]}
   );
   gpc615_5 gpc930 (
      {stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_25[68]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[49],stage1_25[115],stage1_24[162]}
   );
   gpc615_5 gpc931 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245]},
      {stage0_25[69]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[22],stage1_26[50],stage1_25[116],stage1_24[163]}
   );
   gpc615_5 gpc932 (
      {stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_25[70]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[23],stage1_26[51],stage1_25[117],stage1_24[164]}
   );
   gpc615_5 gpc933 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_25[71]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[24],stage1_26[52],stage1_25[118],stage1_24[165]}
   );
   gpc615_5 gpc934 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260]},
      {stage0_25[72]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[25],stage1_26[53],stage1_25[119],stage1_24[166]}
   );
   gpc615_5 gpc935 (
      {stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265]},
      {stage0_25[73]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[26],stage1_26[54],stage1_25[120],stage1_24[167]}
   );
   gpc615_5 gpc936 (
      {stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_25[74]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[27],stage1_26[55],stage1_25[121],stage1_24[168]}
   );
   gpc615_5 gpc937 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275]},
      {stage0_25[75]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[28],stage1_26[56],stage1_25[122],stage1_24[169]}
   );
   gpc615_5 gpc938 (
      {stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_25[76]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[29],stage1_26[57],stage1_25[123],stage1_24[170]}
   );
   gpc615_5 gpc939 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_25[77]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[30],stage1_26[58],stage1_25[124],stage1_24[171]}
   );
   gpc615_5 gpc940 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290]},
      {stage0_25[78]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[31],stage1_26[59],stage1_25[125],stage1_24[172]}
   );
   gpc615_5 gpc941 (
      {stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295]},
      {stage0_25[79]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[32],stage1_26[60],stage1_25[126],stage1_24[173]}
   );
   gpc615_5 gpc942 (
      {stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_25[80]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[33],stage1_26[61],stage1_25[127],stage1_24[174]}
   );
   gpc615_5 gpc943 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305]},
      {stage0_25[81]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[34],stage1_26[62],stage1_25[128],stage1_24[175]}
   );
   gpc615_5 gpc944 (
      {stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_25[82]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[35],stage1_26[63],stage1_25[129],stage1_24[176]}
   );
   gpc615_5 gpc945 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_25[83]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[36],stage1_26[64],stage1_25[130],stage1_24[177]}
   );
   gpc615_5 gpc946 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320]},
      {stage0_25[84]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[37],stage1_26[65],stage1_25[131],stage1_24[178]}
   );
   gpc615_5 gpc947 (
      {stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325]},
      {stage0_25[85]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[38],stage1_26[66],stage1_25[132],stage1_24[179]}
   );
   gpc615_5 gpc948 (
      {stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_25[86]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[39],stage1_26[67],stage1_25[133],stage1_24[180]}
   );
   gpc615_5 gpc949 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335]},
      {stage0_25[87]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[40],stage1_26[68],stage1_25[134],stage1_24[181]}
   );
   gpc615_5 gpc950 (
      {stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_25[88]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[41],stage1_26[69],stage1_25[135],stage1_24[182]}
   );
   gpc615_5 gpc951 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_25[89]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[42],stage1_26[70],stage1_25[136],stage1_24[183]}
   );
   gpc615_5 gpc952 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350]},
      {stage0_25[90]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[43],stage1_26[71],stage1_25[137],stage1_24[184]}
   );
   gpc615_5 gpc953 (
      {stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355]},
      {stage0_25[91]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[44],stage1_26[72],stage1_25[138],stage1_24[185]}
   );
   gpc615_5 gpc954 (
      {stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_25[92]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[45],stage1_26[73],stage1_25[139],stage1_24[186]}
   );
   gpc615_5 gpc955 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365]},
      {stage0_25[93]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[46],stage1_26[74],stage1_25[140],stage1_24[187]}
   );
   gpc615_5 gpc956 (
      {stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_25[94]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[47],stage1_26[75],stage1_25[141],stage1_24[188]}
   );
   gpc615_5 gpc957 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375]},
      {stage0_25[95]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[48],stage1_26[76],stage1_25[142],stage1_24[189]}
   );
   gpc615_5 gpc958 (
      {stage0_24[376], stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380]},
      {stage0_25[96]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[49],stage1_26[77],stage1_25[143],stage1_24[190]}
   );
   gpc615_5 gpc959 (
      {stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385]},
      {stage0_25[97]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[50],stage1_26[78],stage1_25[144],stage1_24[191]}
   );
   gpc615_5 gpc960 (
      {stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_25[98]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[51],stage1_26[79],stage1_25[145],stage1_24[192]}
   );
   gpc615_5 gpc961 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395]},
      {stage0_25[99]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[52],stage1_26[80],stage1_25[146],stage1_24[193]}
   );
   gpc615_5 gpc962 (
      {stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_25[100]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[53],stage1_26[81],stage1_25[147],stage1_24[194]}
   );
   gpc615_5 gpc963 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405]},
      {stage0_25[101]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[54],stage1_26[82],stage1_25[148],stage1_24[195]}
   );
   gpc615_5 gpc964 (
      {stage0_24[406], stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410]},
      {stage0_25[102]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[55],stage1_26[83],stage1_25[149],stage1_24[196]}
   );
   gpc615_5 gpc965 (
      {stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415]},
      {stage0_25[103]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[56],stage1_26[84],stage1_25[150],stage1_24[197]}
   );
   gpc615_5 gpc966 (
      {stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_25[104]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[57],stage1_26[85],stage1_25[151],stage1_24[198]}
   );
   gpc615_5 gpc967 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425]},
      {stage0_25[105]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[58],stage1_26[86],stage1_25[152],stage1_24[199]}
   );
   gpc615_5 gpc968 (
      {stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_25[106]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[59],stage1_26[87],stage1_25[153],stage1_24[200]}
   );
   gpc615_5 gpc969 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435]},
      {stage0_25[107]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[60],stage1_26[88],stage1_25[154],stage1_24[201]}
   );
   gpc615_5 gpc970 (
      {stage0_24[436], stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440]},
      {stage0_25[108]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[61],stage1_26[89],stage1_25[155],stage1_24[202]}
   );
   gpc615_5 gpc971 (
      {stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445]},
      {stage0_25[109]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[62],stage1_26[90],stage1_25[156],stage1_24[203]}
   );
   gpc615_5 gpc972 (
      {stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_25[110]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[63],stage1_26[91],stage1_25[157],stage1_24[204]}
   );
   gpc615_5 gpc973 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455]},
      {stage0_25[111]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[64],stage1_26[92],stage1_25[158],stage1_24[205]}
   );
   gpc615_5 gpc974 (
      {stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_25[112]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[65],stage1_26[93],stage1_25[159],stage1_24[206]}
   );
   gpc615_5 gpc975 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465]},
      {stage0_25[113]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[66],stage1_26[94],stage1_25[160],stage1_24[207]}
   );
   gpc615_5 gpc976 (
      {stage0_24[466], stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470]},
      {stage0_25[114]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[67],stage1_26[95],stage1_25[161],stage1_24[208]}
   );
   gpc615_5 gpc977 (
      {stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475]},
      {stage0_25[115]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[68],stage1_26[96],stage1_25[162],stage1_24[209]}
   );
   gpc615_5 gpc978 (
      {stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_25[116]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[69],stage1_26[97],stage1_25[163],stage1_24[210]}
   );
   gpc615_5 gpc979 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485]},
      {stage0_25[117]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[70],stage1_26[98],stage1_25[164],stage1_24[211]}
   );
   gpc606_5 gpc980 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[61],stage1_27[71],stage1_26[99],stage1_25[165]}
   );
   gpc606_5 gpc981 (
      {stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[62],stage1_27[72],stage1_26[100],stage1_25[166]}
   );
   gpc606_5 gpc982 (
      {stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[63],stage1_27[73],stage1_26[101],stage1_25[167]}
   );
   gpc606_5 gpc983 (
      {stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[64],stage1_27[74],stage1_26[102],stage1_25[168]}
   );
   gpc606_5 gpc984 (
      {stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[65],stage1_27[75],stage1_26[103],stage1_25[169]}
   );
   gpc606_5 gpc985 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[66],stage1_27[76],stage1_26[104],stage1_25[170]}
   );
   gpc606_5 gpc986 (
      {stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[67],stage1_27[77],stage1_26[105],stage1_25[171]}
   );
   gpc606_5 gpc987 (
      {stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[68],stage1_27[78],stage1_26[106],stage1_25[172]}
   );
   gpc606_5 gpc988 (
      {stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[69],stage1_27[79],stage1_26[107],stage1_25[173]}
   );
   gpc606_5 gpc989 (
      {stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[70],stage1_27[80],stage1_26[108],stage1_25[174]}
   );
   gpc606_5 gpc990 (
      {stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[71],stage1_27[81],stage1_26[109],stage1_25[175]}
   );
   gpc606_5 gpc991 (
      {stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[72],stage1_27[82],stage1_26[110],stage1_25[176]}
   );
   gpc606_5 gpc992 (
      {stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[73],stage1_27[83],stage1_26[111],stage1_25[177]}
   );
   gpc606_5 gpc993 (
      {stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[74],stage1_27[84],stage1_26[112],stage1_25[178]}
   );
   gpc606_5 gpc994 (
      {stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[75],stage1_27[85],stage1_26[113],stage1_25[179]}
   );
   gpc606_5 gpc995 (
      {stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[76],stage1_27[86],stage1_26[114],stage1_25[180]}
   );
   gpc606_5 gpc996 (
      {stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[77],stage1_27[87],stage1_26[115],stage1_25[181]}
   );
   gpc606_5 gpc997 (
      {stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[78],stage1_27[88],stage1_26[116],stage1_25[182]}
   );
   gpc615_5 gpc998 (
      {stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229], stage0_25[230]},
      {stage0_26[366]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[79],stage1_27[89],stage1_26[117],stage1_25[183]}
   );
   gpc615_5 gpc999 (
      {stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_26[367]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[80],stage1_27[90],stage1_26[118],stage1_25[184]}
   );
   gpc615_5 gpc1000 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240]},
      {stage0_26[368]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[81],stage1_27[91],stage1_26[119],stage1_25[185]}
   );
   gpc615_5 gpc1001 (
      {stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_26[369]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[82],stage1_27[92],stage1_26[120],stage1_25[186]}
   );
   gpc615_5 gpc1002 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[370]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[83],stage1_27[93],stage1_26[121],stage1_25[187]}
   );
   gpc615_5 gpc1003 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[371]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[84],stage1_27[94],stage1_26[122],stage1_25[188]}
   );
   gpc615_5 gpc1004 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[372]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[85],stage1_27[95],stage1_26[123],stage1_25[189]}
   );
   gpc615_5 gpc1005 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[373]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[86],stage1_27[96],stage1_26[124],stage1_25[190]}
   );
   gpc615_5 gpc1006 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[374]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[87],stage1_27[97],stage1_26[125],stage1_25[191]}
   );
   gpc615_5 gpc1007 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[375]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[88],stage1_27[98],stage1_26[126],stage1_25[192]}
   );
   gpc615_5 gpc1008 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[376]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[89],stage1_27[99],stage1_26[127],stage1_25[193]}
   );
   gpc615_5 gpc1009 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[377]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[90],stage1_27[100],stage1_26[128],stage1_25[194]}
   );
   gpc615_5 gpc1010 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[378]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[91],stage1_27[101],stage1_26[129],stage1_25[195]}
   );
   gpc615_5 gpc1011 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[379]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[92],stage1_27[102],stage1_26[130],stage1_25[196]}
   );
   gpc615_5 gpc1012 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[380]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[93],stage1_27[103],stage1_26[131],stage1_25[197]}
   );
   gpc615_5 gpc1013 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[381]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[94],stage1_27[104],stage1_26[132],stage1_25[198]}
   );
   gpc615_5 gpc1014 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[382]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[95],stage1_27[105],stage1_26[133],stage1_25[199]}
   );
   gpc615_5 gpc1015 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[383]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[96],stage1_27[106],stage1_26[134],stage1_25[200]}
   );
   gpc615_5 gpc1016 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[384]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[97],stage1_27[107],stage1_26[135],stage1_25[201]}
   );
   gpc615_5 gpc1017 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[385]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[98],stage1_27[108],stage1_26[136],stage1_25[202]}
   );
   gpc615_5 gpc1018 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[386]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[99],stage1_27[109],stage1_26[137],stage1_25[203]}
   );
   gpc615_5 gpc1019 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[387]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[100],stage1_27[110],stage1_26[138],stage1_25[204]}
   );
   gpc615_5 gpc1020 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[388]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[101],stage1_27[111],stage1_26[139],stage1_25[205]}
   );
   gpc615_5 gpc1021 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[389]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[102],stage1_27[112],stage1_26[140],stage1_25[206]}
   );
   gpc615_5 gpc1022 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[390]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[103],stage1_27[113],stage1_26[141],stage1_25[207]}
   );
   gpc615_5 gpc1023 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[391]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[104],stage1_27[114],stage1_26[142],stage1_25[208]}
   );
   gpc615_5 gpc1024 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[392]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[105],stage1_27[115],stage1_26[143],stage1_25[209]}
   );
   gpc615_5 gpc1025 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[393]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[106],stage1_27[116],stage1_26[144],stage1_25[210]}
   );
   gpc615_5 gpc1026 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[394]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[107],stage1_27[117],stage1_26[145],stage1_25[211]}
   );
   gpc615_5 gpc1027 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[395]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[108],stage1_27[118],stage1_26[146],stage1_25[212]}
   );
   gpc615_5 gpc1028 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[396]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[109],stage1_27[119],stage1_26[147],stage1_25[213]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[397]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[110],stage1_27[120],stage1_26[148],stage1_25[214]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[398]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[111],stage1_27[121],stage1_26[149],stage1_25[215]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[399]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[112],stage1_27[122],stage1_26[150],stage1_25[216]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[400]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[113],stage1_27[123],stage1_26[151],stage1_25[217]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[401]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[114],stage1_27[124],stage1_26[152],stage1_25[218]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[402]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[115],stage1_27[125],stage1_26[153],stage1_25[219]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[403]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[116],stage1_27[126],stage1_26[154],stage1_25[220]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[404]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[117],stage1_27[127],stage1_26[155],stage1_25[221]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[405]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[118],stage1_27[128],stage1_26[156],stage1_25[222]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[406]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[119],stage1_27[129],stage1_26[157],stage1_25[223]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[407]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[120],stage1_27[130],stage1_26[158],stage1_25[224]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[408]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[121],stage1_27[131],stage1_26[159],stage1_25[225]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[409]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[122],stage1_27[132],stage1_26[160],stage1_25[226]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[410]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[123],stage1_27[133],stage1_26[161],stage1_25[227]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[411]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[124],stage1_27[134],stage1_26[162],stage1_25[228]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[412]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[125],stage1_27[135],stage1_26[163],stage1_25[229]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[413]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[126],stage1_27[136],stage1_26[164],stage1_25[230]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[414]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[127],stage1_27[137],stage1_26[165],stage1_25[231]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[415]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[128],stage1_27[138],stage1_26[166],stage1_25[232]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[416]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[129],stage1_27[139],stage1_26[167],stage1_25[233]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[417]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[130],stage1_27[140],stage1_26[168],stage1_25[234]}
   );
   gpc606_5 gpc1050 (
      {stage0_26[418], stage0_26[419], stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[70],stage1_28[131],stage1_27[141],stage1_26[169]}
   );
   gpc606_5 gpc1051 (
      {stage0_26[424], stage0_26[425], stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[71],stage1_28[132],stage1_27[142],stage1_26[170]}
   );
   gpc615_5 gpc1052 (
      {stage0_26[430], stage0_26[431], stage0_26[432], stage0_26[433], stage0_26[434]},
      {stage0_27[420]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[72],stage1_28[133],stage1_27[143],stage1_26[171]}
   );
   gpc615_5 gpc1053 (
      {stage0_26[435], stage0_26[436], stage0_26[437], stage0_26[438], stage0_26[439]},
      {stage0_27[421]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[73],stage1_28[134],stage1_27[144],stage1_26[172]}
   );
   gpc615_5 gpc1054 (
      {stage0_26[440], stage0_26[441], stage0_26[442], stage0_26[443], stage0_26[444]},
      {stage0_27[422]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[74],stage1_28[135],stage1_27[145],stage1_26[173]}
   );
   gpc606_5 gpc1055 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427], stage0_27[428]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[75],stage1_28[136],stage1_27[146]}
   );
   gpc606_5 gpc1056 (
      {stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432], stage0_27[433], stage0_27[434]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[76],stage1_28[137],stage1_27[147]}
   );
   gpc606_5 gpc1057 (
      {stage0_27[435], stage0_27[436], stage0_27[437], stage0_27[438], stage0_27[439], stage0_27[440]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[77],stage1_28[138],stage1_27[148]}
   );
   gpc606_5 gpc1058 (
      {stage0_27[441], stage0_27[442], stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[78],stage1_28[139],stage1_27[149]}
   );
   gpc606_5 gpc1059 (
      {stage0_27[447], stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[79],stage1_28[140],stage1_27[150]}
   );
   gpc606_5 gpc1060 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457], stage0_27[458]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[80],stage1_28[141],stage1_27[151]}
   );
   gpc606_5 gpc1061 (
      {stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462], stage0_27[463], stage0_27[464]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[81],stage1_28[142],stage1_27[152]}
   );
   gpc606_5 gpc1062 (
      {stage0_27[465], stage0_27[466], stage0_27[467], stage0_27[468], stage0_27[469], stage0_27[470]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[82],stage1_28[143],stage1_27[153]}
   );
   gpc606_5 gpc1063 (
      {stage0_27[471], stage0_27[472], stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[83],stage1_28[144],stage1_27[154]}
   );
   gpc606_5 gpc1064 (
      {stage0_27[477], stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[84],stage1_28[145],stage1_27[155]}
   );
   gpc606_5 gpc1065 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[10],stage1_30[15],stage1_29[85],stage1_28[146]}
   );
   gpc606_5 gpc1066 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[11],stage1_30[16],stage1_29[86],stage1_28[147]}
   );
   gpc606_5 gpc1067 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[12],stage1_30[17],stage1_29[87],stage1_28[148]}
   );
   gpc606_5 gpc1068 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[13],stage1_30[18],stage1_29[88],stage1_28[149]}
   );
   gpc606_5 gpc1069 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[14],stage1_30[19],stage1_29[89],stage1_28[150]}
   );
   gpc606_5 gpc1070 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[15],stage1_30[20],stage1_29[90],stage1_28[151]}
   );
   gpc606_5 gpc1071 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[16],stage1_30[21],stage1_29[91],stage1_28[152]}
   );
   gpc606_5 gpc1072 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[17],stage1_30[22],stage1_29[92],stage1_28[153]}
   );
   gpc606_5 gpc1073 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[18],stage1_30[23],stage1_29[93],stage1_28[154]}
   );
   gpc606_5 gpc1074 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[19],stage1_30[24],stage1_29[94],stage1_28[155]}
   );
   gpc606_5 gpc1075 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[20],stage1_30[25],stage1_29[95],stage1_28[156]}
   );
   gpc606_5 gpc1076 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[21],stage1_30[26],stage1_29[96],stage1_28[157]}
   );
   gpc606_5 gpc1077 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[22],stage1_30[27],stage1_29[97],stage1_28[158]}
   );
   gpc606_5 gpc1078 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[23],stage1_30[28],stage1_29[98],stage1_28[159]}
   );
   gpc606_5 gpc1079 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[24],stage1_30[29],stage1_29[99],stage1_28[160]}
   );
   gpc606_5 gpc1080 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[25],stage1_30[30],stage1_29[100],stage1_28[161]}
   );
   gpc606_5 gpc1081 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[26],stage1_30[31],stage1_29[101],stage1_28[162]}
   );
   gpc606_5 gpc1082 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[27],stage1_30[32],stage1_29[102],stage1_28[163]}
   );
   gpc606_5 gpc1083 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[28],stage1_30[33],stage1_29[103],stage1_28[164]}
   );
   gpc606_5 gpc1084 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[29],stage1_30[34],stage1_29[104],stage1_28[165]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[30],stage1_30[35],stage1_29[105],stage1_28[166]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[31],stage1_30[36],stage1_29[106],stage1_28[167]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[32],stage1_30[37],stage1_29[107],stage1_28[168]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[33],stage1_30[38],stage1_29[108],stage1_28[169]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[34],stage1_30[39],stage1_29[109],stage1_28[170]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[35],stage1_30[40],stage1_29[110],stage1_28[171]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[36],stage1_30[41],stage1_29[111],stage1_28[172]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[37],stage1_30[42],stage1_29[112],stage1_28[173]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[38],stage1_30[43],stage1_29[113],stage1_28[174]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[39],stage1_30[44],stage1_29[114],stage1_28[175]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[40],stage1_30[45],stage1_29[115],stage1_28[176]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[41],stage1_30[46],stage1_29[116],stage1_28[177]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[42],stage1_30[47],stage1_29[117],stage1_28[178]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[43],stage1_30[48],stage1_29[118],stage1_28[179]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[44],stage1_30[49],stage1_29[119],stage1_28[180]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[240], stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[45],stage1_30[50],stage1_29[120],stage1_28[181]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[246], stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[46],stage1_30[51],stage1_29[121],stage1_28[182]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[252], stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[47],stage1_30[52],stage1_29[122],stage1_28[183]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[258], stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[48],stage1_30[53],stage1_29[123],stage1_28[184]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[264], stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[49],stage1_30[54],stage1_29[124],stage1_28[185]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[270], stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[50],stage1_30[55],stage1_29[125],stage1_28[186]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[276], stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[51],stage1_30[56],stage1_29[126],stage1_28[187]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[282], stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[52],stage1_30[57],stage1_29[127],stage1_28[188]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[288], stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[53],stage1_30[58],stage1_29[128],stage1_28[189]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[294], stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[54],stage1_30[59],stage1_29[129],stage1_28[190]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[300], stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[55],stage1_30[60],stage1_29[130],stage1_28[191]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[56],stage1_30[61],stage1_29[131],stage1_28[192]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[57],stage1_30[62],stage1_29[132],stage1_28[193]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[318], stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[58],stage1_30[63],stage1_29[133],stage1_28[194]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[324], stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[59],stage1_30[64],stage1_29[134],stage1_28[195]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[330], stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[60],stage1_30[65],stage1_29[135],stage1_28[196]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[61],stage1_30[66],stage1_29[136],stage1_28[197]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[62],stage1_30[67],stage1_29[137],stage1_28[198]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[348], stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[63],stage1_30[68],stage1_29[138],stage1_28[199]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[354], stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[64],stage1_30[69],stage1_29[139],stage1_28[200]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[360], stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[65],stage1_30[70],stage1_29[140],stage1_28[201]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[66],stage1_30[71],stage1_29[141],stage1_28[202]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[67],stage1_30[72],stage1_29[142],stage1_28[203]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[378], stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[68],stage1_30[73],stage1_29[143],stage1_28[204]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[384], stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[69],stage1_30[74],stage1_29[144],stage1_28[205]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[390], stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[70],stage1_30[75],stage1_29[145],stage1_28[206]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[71],stage1_30[76],stage1_29[146],stage1_28[207]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[72],stage1_30[77],stage1_29[147],stage1_28[208]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[408], stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[73],stage1_30[78],stage1_29[148],stage1_28[209]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[414], stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[74],stage1_30[79],stage1_29[149],stage1_28[210]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[420], stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[75],stage1_30[80],stage1_29[150],stage1_28[211]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[76],stage1_30[81],stage1_29[151],stage1_28[212]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[77],stage1_30[82],stage1_29[152],stage1_28[213]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[438], stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[78],stage1_30[83],stage1_29[153],stage1_28[214]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[444], stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[79],stage1_30[84],stage1_29[154],stage1_28[215]}
   );
   gpc606_5 gpc1135 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[70],stage1_31[80],stage1_30[85],stage1_29[155]}
   );
   gpc606_5 gpc1136 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[71],stage1_31[81],stage1_30[86],stage1_29[156]}
   );
   gpc606_5 gpc1137 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[72],stage1_31[82],stage1_30[87],stage1_29[157]}
   );
   gpc606_5 gpc1138 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[73],stage1_31[83],stage1_30[88],stage1_29[158]}
   );
   gpc606_5 gpc1139 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[74],stage1_31[84],stage1_30[89],stage1_29[159]}
   );
   gpc606_5 gpc1140 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[75],stage1_31[85],stage1_30[90],stage1_29[160]}
   );
   gpc606_5 gpc1141 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[76],stage1_31[86],stage1_30[91],stage1_29[161]}
   );
   gpc606_5 gpc1142 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[77],stage1_31[87],stage1_30[92],stage1_29[162]}
   );
   gpc606_5 gpc1143 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[78],stage1_31[88],stage1_30[93],stage1_29[163]}
   );
   gpc606_5 gpc1144 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[79],stage1_31[89],stage1_30[94],stage1_29[164]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[80],stage1_31[90],stage1_30[95],stage1_29[165]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[81],stage1_31[91],stage1_30[96],stage1_29[166]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[82],stage1_31[92],stage1_30[97],stage1_29[167]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[83],stage1_31[93],stage1_30[98],stage1_29[168]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[84],stage1_31[94],stage1_30[99],stage1_29[169]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[85],stage1_31[95],stage1_30[100],stage1_29[170]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[86],stage1_31[96],stage1_30[101],stage1_29[171]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[87],stage1_31[97],stage1_30[102],stage1_29[172]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[88],stage1_31[98],stage1_30[103],stage1_29[173]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[89],stage1_31[99],stage1_30[104],stage1_29[174]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[90],stage1_31[100],stage1_30[105],stage1_29[175]}
   );
   gpc615_5 gpc1156 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_30[420]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[91],stage1_31[101],stage1_30[106],stage1_29[176]}
   );
   gpc615_5 gpc1157 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195]},
      {stage0_30[421]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[92],stage1_31[102],stage1_30[107],stage1_29[177]}
   );
   gpc615_5 gpc1158 (
      {stage0_29[196], stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200]},
      {stage0_30[422]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[93],stage1_31[103],stage1_30[108],stage1_29[178]}
   );
   gpc615_5 gpc1159 (
      {stage0_29[201], stage0_29[202], stage0_29[203], stage0_29[204], stage0_29[205]},
      {stage0_30[423]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[94],stage1_31[104],stage1_30[109],stage1_29[179]}
   );
   gpc615_5 gpc1160 (
      {stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209], stage0_29[210]},
      {stage0_30[424]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[95],stage1_31[105],stage1_30[110],stage1_29[180]}
   );
   gpc615_5 gpc1161 (
      {stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_30[425]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[96],stage1_31[106],stage1_30[111],stage1_29[181]}
   );
   gpc615_5 gpc1162 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_30[426]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[97],stage1_31[107],stage1_30[112],stage1_29[182]}
   );
   gpc615_5 gpc1163 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225]},
      {stage0_30[427]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[98],stage1_31[108],stage1_30[113],stage1_29[183]}
   );
   gpc615_5 gpc1164 (
      {stage0_29[226], stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230]},
      {stage0_30[428]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[99],stage1_31[109],stage1_30[114],stage1_29[184]}
   );
   gpc615_5 gpc1165 (
      {stage0_29[231], stage0_29[232], stage0_29[233], stage0_29[234], stage0_29[235]},
      {stage0_30[429]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[100],stage1_31[110],stage1_30[115],stage1_29[185]}
   );
   gpc615_5 gpc1166 (
      {stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239], stage0_29[240]},
      {stage0_30[430]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[101],stage1_31[111],stage1_30[116],stage1_29[186]}
   );
   gpc615_5 gpc1167 (
      {stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_30[431]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[102],stage1_31[112],stage1_30[117],stage1_29[187]}
   );
   gpc615_5 gpc1168 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_30[432]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[103],stage1_31[113],stage1_30[118],stage1_29[188]}
   );
   gpc615_5 gpc1169 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255]},
      {stage0_30[433]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[104],stage1_31[114],stage1_30[119],stage1_29[189]}
   );
   gpc615_5 gpc1170 (
      {stage0_29[256], stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260]},
      {stage0_30[434]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[105],stage1_31[115],stage1_30[120],stage1_29[190]}
   );
   gpc615_5 gpc1171 (
      {stage0_29[261], stage0_29[262], stage0_29[263], stage0_29[264], stage0_29[265]},
      {stage0_30[435]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[106],stage1_31[116],stage1_30[121],stage1_29[191]}
   );
   gpc615_5 gpc1172 (
      {stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269], stage0_29[270]},
      {stage0_30[436]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[107],stage1_31[117],stage1_30[122],stage1_29[192]}
   );
   gpc615_5 gpc1173 (
      {stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_30[437]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[108],stage1_31[118],stage1_30[123],stage1_29[193]}
   );
   gpc615_5 gpc1174 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_30[438]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[109],stage1_31[119],stage1_30[124],stage1_29[194]}
   );
   gpc615_5 gpc1175 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285]},
      {stage0_30[439]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[110],stage1_31[120],stage1_30[125],stage1_29[195]}
   );
   gpc615_5 gpc1176 (
      {stage0_29[286], stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290]},
      {stage0_30[440]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[111],stage1_31[121],stage1_30[126],stage1_29[196]}
   );
   gpc615_5 gpc1177 (
      {stage0_29[291], stage0_29[292], stage0_29[293], stage0_29[294], stage0_29[295]},
      {stage0_30[441]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[112],stage1_31[122],stage1_30[127],stage1_29[197]}
   );
   gpc615_5 gpc1178 (
      {stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299], stage0_29[300]},
      {stage0_30[442]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[113],stage1_31[123],stage1_30[128],stage1_29[198]}
   );
   gpc615_5 gpc1179 (
      {stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_30[443]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[114],stage1_31[124],stage1_30[129],stage1_29[199]}
   );
   gpc615_5 gpc1180 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_30[444]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[115],stage1_31[125],stage1_30[130],stage1_29[200]}
   );
   gpc615_5 gpc1181 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315]},
      {stage0_30[445]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[116],stage1_31[126],stage1_30[131],stage1_29[201]}
   );
   gpc615_5 gpc1182 (
      {stage0_29[316], stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320]},
      {stage0_30[446]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[117],stage1_31[127],stage1_30[132],stage1_29[202]}
   );
   gpc615_5 gpc1183 (
      {stage0_29[321], stage0_29[322], stage0_29[323], stage0_29[324], stage0_29[325]},
      {stage0_30[447]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[118],stage1_31[128],stage1_30[133],stage1_29[203]}
   );
   gpc615_5 gpc1184 (
      {stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329], stage0_29[330]},
      {stage0_30[448]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[119],stage1_31[129],stage1_30[134],stage1_29[204]}
   );
   gpc615_5 gpc1185 (
      {stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_30[449]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[120],stage1_31[130],stage1_30[135],stage1_29[205]}
   );
   gpc615_5 gpc1186 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_30[450]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[121],stage1_31[131],stage1_30[136],stage1_29[206]}
   );
   gpc615_5 gpc1187 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345]},
      {stage0_30[451]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[122],stage1_31[132],stage1_30[137],stage1_29[207]}
   );
   gpc615_5 gpc1188 (
      {stage0_29[346], stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350]},
      {stage0_30[452]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[123],stage1_31[133],stage1_30[138],stage1_29[208]}
   );
   gpc615_5 gpc1189 (
      {stage0_29[351], stage0_29[352], stage0_29[353], stage0_29[354], stage0_29[355]},
      {stage0_30[453]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[124],stage1_31[134],stage1_30[139],stage1_29[209]}
   );
   gpc615_5 gpc1190 (
      {stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359], stage0_29[360]},
      {stage0_30[454]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[125],stage1_31[135],stage1_30[140],stage1_29[210]}
   );
   gpc615_5 gpc1191 (
      {stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_30[455]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[126],stage1_31[136],stage1_30[141],stage1_29[211]}
   );
   gpc615_5 gpc1192 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_30[456]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[127],stage1_31[137],stage1_30[142],stage1_29[212]}
   );
   gpc615_5 gpc1193 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375]},
      {stage0_30[457]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[128],stage1_31[138],stage1_30[143],stage1_29[213]}
   );
   gpc615_5 gpc1194 (
      {stage0_29[376], stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380]},
      {stage0_30[458]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[129],stage1_31[139],stage1_30[144],stage1_29[214]}
   );
   gpc615_5 gpc1195 (
      {stage0_29[381], stage0_29[382], stage0_29[383], stage0_29[384], stage0_29[385]},
      {stage0_30[459]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[130],stage1_31[140],stage1_30[145],stage1_29[215]}
   );
   gpc615_5 gpc1196 (
      {stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389], stage0_29[390]},
      {stage0_30[460]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[131],stage1_31[141],stage1_30[146],stage1_29[216]}
   );
   gpc615_5 gpc1197 (
      {stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_30[461]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[132],stage1_31[142],stage1_30[147],stage1_29[217]}
   );
   gpc615_5 gpc1198 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_30[462]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[133],stage1_31[143],stage1_30[148],stage1_29[218]}
   );
   gpc615_5 gpc1199 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405]},
      {stage0_30[463]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[134],stage1_31[144],stage1_30[149],stage1_29[219]}
   );
   gpc615_5 gpc1200 (
      {stage0_29[406], stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410]},
      {stage0_30[464]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[135],stage1_31[145],stage1_30[150],stage1_29[220]}
   );
   gpc615_5 gpc1201 (
      {stage0_29[411], stage0_29[412], stage0_29[413], stage0_29[414], stage0_29[415]},
      {stage0_30[465]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[136],stage1_31[146],stage1_30[151],stage1_29[221]}
   );
   gpc615_5 gpc1202 (
      {stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419], stage0_29[420]},
      {stage0_30[466]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[137],stage1_31[147],stage1_30[152],stage1_29[222]}
   );
   gpc615_5 gpc1203 (
      {stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_30[467]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[138],stage1_31[148],stage1_30[153],stage1_29[223]}
   );
   gpc615_5 gpc1204 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_30[468]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[139],stage1_31[149],stage1_30[154],stage1_29[224]}
   );
   gpc615_5 gpc1205 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435]},
      {stage0_30[469]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[140],stage1_31[150],stage1_30[155],stage1_29[225]}
   );
   gpc615_5 gpc1206 (
      {stage0_29[436], stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440]},
      {stage0_30[470]},
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430], stage0_31[431]},
      {stage1_33[71],stage1_32[141],stage1_31[151],stage1_30[156],stage1_29[226]}
   );
   gpc615_5 gpc1207 (
      {stage0_29[441], stage0_29[442], stage0_29[443], stage0_29[444], stage0_29[445]},
      {stage0_30[471]},
      {stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437]},
      {stage1_33[72],stage1_32[142],stage1_31[152],stage1_30[157],stage1_29[227]}
   );
   gpc615_5 gpc1208 (
      {stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449], stage0_29[450]},
      {stage0_30[472]},
      {stage0_31[438], stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage1_33[73],stage1_32[143],stage1_31[153],stage1_30[158],stage1_29[228]}
   );
   gpc615_5 gpc1209 (
      {stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_30[473]},
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449]},
      {stage1_33[74],stage1_32[144],stage1_31[154],stage1_30[159],stage1_29[229]}
   );
   gpc615_5 gpc1210 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_30[474]},
      {stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage1_33[75],stage1_32[145],stage1_31[155],stage1_30[160],stage1_29[230]}
   );
   gpc615_5 gpc1211 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465]},
      {stage0_30[475]},
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460], stage0_31[461]},
      {stage1_33[76],stage1_32[146],stage1_31[156],stage1_30[161],stage1_29[231]}
   );
   gpc615_5 gpc1212 (
      {stage0_29[466], stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470]},
      {stage0_30[476]},
      {stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467]},
      {stage1_33[77],stage1_32[147],stage1_31[157],stage1_30[162],stage1_29[232]}
   );
   gpc615_5 gpc1213 (
      {stage0_29[471], stage0_29[472], stage0_29[473], stage0_29[474], stage0_29[475]},
      {stage0_30[477]},
      {stage0_31[468], stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage1_33[78],stage1_32[148],stage1_31[158],stage1_30[163],stage1_29[233]}
   );
   gpc615_5 gpc1214 (
      {stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479], stage0_29[480]},
      {stage0_30[478]},
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478], stage0_31[479]},
      {stage1_33[79],stage1_32[149],stage1_31[159],stage1_30[164],stage1_29[234]}
   );
   gpc615_5 gpc1215 (
      {stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_30[479]},
      {stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483], stage0_31[484], stage0_31[485]},
      {stage1_33[80],stage1_32[150],stage1_31[160],stage1_30[165],stage1_29[235]}
   );
   gpc1_1 gpc1216 (
      {stage0_0[444]},
      {stage1_0[85]}
   );
   gpc1_1 gpc1217 (
      {stage0_0[445]},
      {stage1_0[86]}
   );
   gpc1_1 gpc1218 (
      {stage0_0[446]},
      {stage1_0[87]}
   );
   gpc1_1 gpc1219 (
      {stage0_0[447]},
      {stage1_0[88]}
   );
   gpc1_1 gpc1220 (
      {stage0_0[448]},
      {stage1_0[89]}
   );
   gpc1_1 gpc1221 (
      {stage0_0[449]},
      {stage1_0[90]}
   );
   gpc1_1 gpc1222 (
      {stage0_0[450]},
      {stage1_0[91]}
   );
   gpc1_1 gpc1223 (
      {stage0_0[451]},
      {stage1_0[92]}
   );
   gpc1_1 gpc1224 (
      {stage0_0[452]},
      {stage1_0[93]}
   );
   gpc1_1 gpc1225 (
      {stage0_0[453]},
      {stage1_0[94]}
   );
   gpc1_1 gpc1226 (
      {stage0_0[454]},
      {stage1_0[95]}
   );
   gpc1_1 gpc1227 (
      {stage0_0[455]},
      {stage1_0[96]}
   );
   gpc1_1 gpc1228 (
      {stage0_0[456]},
      {stage1_0[97]}
   );
   gpc1_1 gpc1229 (
      {stage0_0[457]},
      {stage1_0[98]}
   );
   gpc1_1 gpc1230 (
      {stage0_0[458]},
      {stage1_0[99]}
   );
   gpc1_1 gpc1231 (
      {stage0_0[459]},
      {stage1_0[100]}
   );
   gpc1_1 gpc1232 (
      {stage0_0[460]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1233 (
      {stage0_0[461]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1234 (
      {stage0_0[462]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1235 (
      {stage0_0[463]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1236 (
      {stage0_0[464]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1237 (
      {stage0_0[465]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1238 (
      {stage0_0[466]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1239 (
      {stage0_0[467]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1240 (
      {stage0_0[468]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1241 (
      {stage0_0[469]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1242 (
      {stage0_0[470]},
      {stage1_0[111]}
   );
   gpc1_1 gpc1243 (
      {stage0_0[471]},
      {stage1_0[112]}
   );
   gpc1_1 gpc1244 (
      {stage0_0[472]},
      {stage1_0[113]}
   );
   gpc1_1 gpc1245 (
      {stage0_0[473]},
      {stage1_0[114]}
   );
   gpc1_1 gpc1246 (
      {stage0_0[474]},
      {stage1_0[115]}
   );
   gpc1_1 gpc1247 (
      {stage0_0[475]},
      {stage1_0[116]}
   );
   gpc1_1 gpc1248 (
      {stage0_0[476]},
      {stage1_0[117]}
   );
   gpc1_1 gpc1249 (
      {stage0_0[477]},
      {stage1_0[118]}
   );
   gpc1_1 gpc1250 (
      {stage0_0[478]},
      {stage1_0[119]}
   );
   gpc1_1 gpc1251 (
      {stage0_0[479]},
      {stage1_0[120]}
   );
   gpc1_1 gpc1252 (
      {stage0_0[480]},
      {stage1_0[121]}
   );
   gpc1_1 gpc1253 (
      {stage0_0[481]},
      {stage1_0[122]}
   );
   gpc1_1 gpc1254 (
      {stage0_0[482]},
      {stage1_0[123]}
   );
   gpc1_1 gpc1255 (
      {stage0_0[483]},
      {stage1_0[124]}
   );
   gpc1_1 gpc1256 (
      {stage0_0[484]},
      {stage1_0[125]}
   );
   gpc1_1 gpc1257 (
      {stage0_0[485]},
      {stage1_0[126]}
   );
   gpc1_1 gpc1258 (
      {stage0_1[484]},
      {stage1_1[136]}
   );
   gpc1_1 gpc1259 (
      {stage0_1[485]},
      {stage1_1[137]}
   );
   gpc1_1 gpc1260 (
      {stage0_2[415]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1261 (
      {stage0_2[416]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1262 (
      {stage0_2[417]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1263 (
      {stage0_2[418]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1264 (
      {stage0_2[419]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1265 (
      {stage0_2[420]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1266 (
      {stage0_2[421]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1267 (
      {stage0_2[422]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1268 (
      {stage0_2[423]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1269 (
      {stage0_2[424]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1270 (
      {stage0_2[425]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1271 (
      {stage0_2[426]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1272 (
      {stage0_2[427]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1273 (
      {stage0_2[428]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1274 (
      {stage0_2[429]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1275 (
      {stage0_2[430]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1276 (
      {stage0_2[431]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1277 (
      {stage0_2[432]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1278 (
      {stage0_2[433]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1279 (
      {stage0_2[434]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1280 (
      {stage0_2[435]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1281 (
      {stage0_2[436]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1282 (
      {stage0_2[437]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1283 (
      {stage0_2[438]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1284 (
      {stage0_2[439]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1285 (
      {stage0_2[440]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1286 (
      {stage0_2[441]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1287 (
      {stage0_2[442]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1288 (
      {stage0_2[443]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1289 (
      {stage0_2[444]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1290 (
      {stage0_2[445]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1291 (
      {stage0_2[446]},
      {stage1_2[188]}
   );
   gpc1_1 gpc1292 (
      {stage0_2[447]},
      {stage1_2[189]}
   );
   gpc1_1 gpc1293 (
      {stage0_2[448]},
      {stage1_2[190]}
   );
   gpc1_1 gpc1294 (
      {stage0_2[449]},
      {stage1_2[191]}
   );
   gpc1_1 gpc1295 (
      {stage0_2[450]},
      {stage1_2[192]}
   );
   gpc1_1 gpc1296 (
      {stage0_2[451]},
      {stage1_2[193]}
   );
   gpc1_1 gpc1297 (
      {stage0_2[452]},
      {stage1_2[194]}
   );
   gpc1_1 gpc1298 (
      {stage0_2[453]},
      {stage1_2[195]}
   );
   gpc1_1 gpc1299 (
      {stage0_2[454]},
      {stage1_2[196]}
   );
   gpc1_1 gpc1300 (
      {stage0_2[455]},
      {stage1_2[197]}
   );
   gpc1_1 gpc1301 (
      {stage0_2[456]},
      {stage1_2[198]}
   );
   gpc1_1 gpc1302 (
      {stage0_2[457]},
      {stage1_2[199]}
   );
   gpc1_1 gpc1303 (
      {stage0_2[458]},
      {stage1_2[200]}
   );
   gpc1_1 gpc1304 (
      {stage0_2[459]},
      {stage1_2[201]}
   );
   gpc1_1 gpc1305 (
      {stage0_2[460]},
      {stage1_2[202]}
   );
   gpc1_1 gpc1306 (
      {stage0_2[461]},
      {stage1_2[203]}
   );
   gpc1_1 gpc1307 (
      {stage0_2[462]},
      {stage1_2[204]}
   );
   gpc1_1 gpc1308 (
      {stage0_2[463]},
      {stage1_2[205]}
   );
   gpc1_1 gpc1309 (
      {stage0_2[464]},
      {stage1_2[206]}
   );
   gpc1_1 gpc1310 (
      {stage0_2[465]},
      {stage1_2[207]}
   );
   gpc1_1 gpc1311 (
      {stage0_2[466]},
      {stage1_2[208]}
   );
   gpc1_1 gpc1312 (
      {stage0_2[467]},
      {stage1_2[209]}
   );
   gpc1_1 gpc1313 (
      {stage0_2[468]},
      {stage1_2[210]}
   );
   gpc1_1 gpc1314 (
      {stage0_2[469]},
      {stage1_2[211]}
   );
   gpc1_1 gpc1315 (
      {stage0_2[470]},
      {stage1_2[212]}
   );
   gpc1_1 gpc1316 (
      {stage0_2[471]},
      {stage1_2[213]}
   );
   gpc1_1 gpc1317 (
      {stage0_2[472]},
      {stage1_2[214]}
   );
   gpc1_1 gpc1318 (
      {stage0_2[473]},
      {stage1_2[215]}
   );
   gpc1_1 gpc1319 (
      {stage0_2[474]},
      {stage1_2[216]}
   );
   gpc1_1 gpc1320 (
      {stage0_2[475]},
      {stage1_2[217]}
   );
   gpc1_1 gpc1321 (
      {stage0_2[476]},
      {stage1_2[218]}
   );
   gpc1_1 gpc1322 (
      {stage0_2[477]},
      {stage1_2[219]}
   );
   gpc1_1 gpc1323 (
      {stage0_2[478]},
      {stage1_2[220]}
   );
   gpc1_1 gpc1324 (
      {stage0_2[479]},
      {stage1_2[221]}
   );
   gpc1_1 gpc1325 (
      {stage0_2[480]},
      {stage1_2[222]}
   );
   gpc1_1 gpc1326 (
      {stage0_2[481]},
      {stage1_2[223]}
   );
   gpc1_1 gpc1327 (
      {stage0_2[482]},
      {stage1_2[224]}
   );
   gpc1_1 gpc1328 (
      {stage0_2[483]},
      {stage1_2[225]}
   );
   gpc1_1 gpc1329 (
      {stage0_2[484]},
      {stage1_2[226]}
   );
   gpc1_1 gpc1330 (
      {stage0_2[485]},
      {stage1_2[227]}
   );
   gpc1_1 gpc1331 (
      {stage0_3[484]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1332 (
      {stage0_3[485]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1333 (
      {stage0_4[485]},
      {stage1_4[225]}
   );
   gpc1_1 gpc1334 (
      {stage0_5[474]},
      {stage1_5[206]}
   );
   gpc1_1 gpc1335 (
      {stage0_5[475]},
      {stage1_5[207]}
   );
   gpc1_1 gpc1336 (
      {stage0_5[476]},
      {stage1_5[208]}
   );
   gpc1_1 gpc1337 (
      {stage0_5[477]},
      {stage1_5[209]}
   );
   gpc1_1 gpc1338 (
      {stage0_5[478]},
      {stage1_5[210]}
   );
   gpc1_1 gpc1339 (
      {stage0_5[479]},
      {stage1_5[211]}
   );
   gpc1_1 gpc1340 (
      {stage0_5[480]},
      {stage1_5[212]}
   );
   gpc1_1 gpc1341 (
      {stage0_5[481]},
      {stage1_5[213]}
   );
   gpc1_1 gpc1342 (
      {stage0_5[482]},
      {stage1_5[214]}
   );
   gpc1_1 gpc1343 (
      {stage0_5[483]},
      {stage1_5[215]}
   );
   gpc1_1 gpc1344 (
      {stage0_5[484]},
      {stage1_5[216]}
   );
   gpc1_1 gpc1345 (
      {stage0_5[485]},
      {stage1_5[217]}
   );
   gpc1_1 gpc1346 (
      {stage0_6[410]},
      {stage1_6[171]}
   );
   gpc1_1 gpc1347 (
      {stage0_6[411]},
      {stage1_6[172]}
   );
   gpc1_1 gpc1348 (
      {stage0_6[412]},
      {stage1_6[173]}
   );
   gpc1_1 gpc1349 (
      {stage0_6[413]},
      {stage1_6[174]}
   );
   gpc1_1 gpc1350 (
      {stage0_6[414]},
      {stage1_6[175]}
   );
   gpc1_1 gpc1351 (
      {stage0_6[415]},
      {stage1_6[176]}
   );
   gpc1_1 gpc1352 (
      {stage0_6[416]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1353 (
      {stage0_6[417]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1354 (
      {stage0_6[418]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1355 (
      {stage0_6[419]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1356 (
      {stage0_6[420]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1357 (
      {stage0_6[421]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1358 (
      {stage0_6[422]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1359 (
      {stage0_6[423]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1360 (
      {stage0_6[424]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1361 (
      {stage0_6[425]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1362 (
      {stage0_6[426]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1363 (
      {stage0_6[427]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1364 (
      {stage0_6[428]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1365 (
      {stage0_6[429]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1366 (
      {stage0_6[430]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1367 (
      {stage0_6[431]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1368 (
      {stage0_6[432]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1369 (
      {stage0_6[433]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1370 (
      {stage0_6[434]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1371 (
      {stage0_6[435]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1372 (
      {stage0_6[436]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1373 (
      {stage0_6[437]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1374 (
      {stage0_6[438]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1375 (
      {stage0_6[439]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1376 (
      {stage0_6[440]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1377 (
      {stage0_6[441]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1378 (
      {stage0_6[442]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1379 (
      {stage0_6[443]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1380 (
      {stage0_6[444]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1381 (
      {stage0_6[445]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1382 (
      {stage0_6[446]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1383 (
      {stage0_6[447]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1384 (
      {stage0_6[448]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1385 (
      {stage0_6[449]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1386 (
      {stage0_6[450]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1387 (
      {stage0_6[451]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1388 (
      {stage0_6[452]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1389 (
      {stage0_6[453]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1390 (
      {stage0_6[454]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1391 (
      {stage0_6[455]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1392 (
      {stage0_6[456]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1393 (
      {stage0_6[457]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1394 (
      {stage0_6[458]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1395 (
      {stage0_6[459]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1396 (
      {stage0_6[460]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1397 (
      {stage0_6[461]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1398 (
      {stage0_6[462]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1399 (
      {stage0_6[463]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1400 (
      {stage0_6[464]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1401 (
      {stage0_6[465]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1402 (
      {stage0_6[466]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1403 (
      {stage0_6[467]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1404 (
      {stage0_6[468]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1405 (
      {stage0_6[469]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1406 (
      {stage0_6[470]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1407 (
      {stage0_6[471]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1408 (
      {stage0_6[472]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1409 (
      {stage0_6[473]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1410 (
      {stage0_6[474]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1411 (
      {stage0_6[475]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1412 (
      {stage0_6[476]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1413 (
      {stage0_6[477]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1414 (
      {stage0_6[478]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1415 (
      {stage0_6[479]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1416 (
      {stage0_6[480]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1417 (
      {stage0_6[481]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1418 (
      {stage0_6[482]},
      {stage1_6[243]}
   );
   gpc1_1 gpc1419 (
      {stage0_6[483]},
      {stage1_6[244]}
   );
   gpc1_1 gpc1420 (
      {stage0_6[484]},
      {stage1_6[245]}
   );
   gpc1_1 gpc1421 (
      {stage0_6[485]},
      {stage1_6[246]}
   );
   gpc1_1 gpc1422 (
      {stage0_7[436]},
      {stage1_7[174]}
   );
   gpc1_1 gpc1423 (
      {stage0_7[437]},
      {stage1_7[175]}
   );
   gpc1_1 gpc1424 (
      {stage0_7[438]},
      {stage1_7[176]}
   );
   gpc1_1 gpc1425 (
      {stage0_7[439]},
      {stage1_7[177]}
   );
   gpc1_1 gpc1426 (
      {stage0_7[440]},
      {stage1_7[178]}
   );
   gpc1_1 gpc1427 (
      {stage0_7[441]},
      {stage1_7[179]}
   );
   gpc1_1 gpc1428 (
      {stage0_7[442]},
      {stage1_7[180]}
   );
   gpc1_1 gpc1429 (
      {stage0_7[443]},
      {stage1_7[181]}
   );
   gpc1_1 gpc1430 (
      {stage0_7[444]},
      {stage1_7[182]}
   );
   gpc1_1 gpc1431 (
      {stage0_7[445]},
      {stage1_7[183]}
   );
   gpc1_1 gpc1432 (
      {stage0_7[446]},
      {stage1_7[184]}
   );
   gpc1_1 gpc1433 (
      {stage0_7[447]},
      {stage1_7[185]}
   );
   gpc1_1 gpc1434 (
      {stage0_7[448]},
      {stage1_7[186]}
   );
   gpc1_1 gpc1435 (
      {stage0_7[449]},
      {stage1_7[187]}
   );
   gpc1_1 gpc1436 (
      {stage0_7[450]},
      {stage1_7[188]}
   );
   gpc1_1 gpc1437 (
      {stage0_7[451]},
      {stage1_7[189]}
   );
   gpc1_1 gpc1438 (
      {stage0_7[452]},
      {stage1_7[190]}
   );
   gpc1_1 gpc1439 (
      {stage0_7[453]},
      {stage1_7[191]}
   );
   gpc1_1 gpc1440 (
      {stage0_7[454]},
      {stage1_7[192]}
   );
   gpc1_1 gpc1441 (
      {stage0_7[455]},
      {stage1_7[193]}
   );
   gpc1_1 gpc1442 (
      {stage0_7[456]},
      {stage1_7[194]}
   );
   gpc1_1 gpc1443 (
      {stage0_7[457]},
      {stage1_7[195]}
   );
   gpc1_1 gpc1444 (
      {stage0_7[458]},
      {stage1_7[196]}
   );
   gpc1_1 gpc1445 (
      {stage0_7[459]},
      {stage1_7[197]}
   );
   gpc1_1 gpc1446 (
      {stage0_7[460]},
      {stage1_7[198]}
   );
   gpc1_1 gpc1447 (
      {stage0_7[461]},
      {stage1_7[199]}
   );
   gpc1_1 gpc1448 (
      {stage0_7[462]},
      {stage1_7[200]}
   );
   gpc1_1 gpc1449 (
      {stage0_7[463]},
      {stage1_7[201]}
   );
   gpc1_1 gpc1450 (
      {stage0_7[464]},
      {stage1_7[202]}
   );
   gpc1_1 gpc1451 (
      {stage0_7[465]},
      {stage1_7[203]}
   );
   gpc1_1 gpc1452 (
      {stage0_7[466]},
      {stage1_7[204]}
   );
   gpc1_1 gpc1453 (
      {stage0_7[467]},
      {stage1_7[205]}
   );
   gpc1_1 gpc1454 (
      {stage0_7[468]},
      {stage1_7[206]}
   );
   gpc1_1 gpc1455 (
      {stage0_7[469]},
      {stage1_7[207]}
   );
   gpc1_1 gpc1456 (
      {stage0_7[470]},
      {stage1_7[208]}
   );
   gpc1_1 gpc1457 (
      {stage0_7[471]},
      {stage1_7[209]}
   );
   gpc1_1 gpc1458 (
      {stage0_7[472]},
      {stage1_7[210]}
   );
   gpc1_1 gpc1459 (
      {stage0_7[473]},
      {stage1_7[211]}
   );
   gpc1_1 gpc1460 (
      {stage0_7[474]},
      {stage1_7[212]}
   );
   gpc1_1 gpc1461 (
      {stage0_7[475]},
      {stage1_7[213]}
   );
   gpc1_1 gpc1462 (
      {stage0_7[476]},
      {stage1_7[214]}
   );
   gpc1_1 gpc1463 (
      {stage0_7[477]},
      {stage1_7[215]}
   );
   gpc1_1 gpc1464 (
      {stage0_7[478]},
      {stage1_7[216]}
   );
   gpc1_1 gpc1465 (
      {stage0_7[479]},
      {stage1_7[217]}
   );
   gpc1_1 gpc1466 (
      {stage0_7[480]},
      {stage1_7[218]}
   );
   gpc1_1 gpc1467 (
      {stage0_7[481]},
      {stage1_7[219]}
   );
   gpc1_1 gpc1468 (
      {stage0_7[482]},
      {stage1_7[220]}
   );
   gpc1_1 gpc1469 (
      {stage0_7[483]},
      {stage1_7[221]}
   );
   gpc1_1 gpc1470 (
      {stage0_7[484]},
      {stage1_7[222]}
   );
   gpc1_1 gpc1471 (
      {stage0_7[485]},
      {stage1_7[223]}
   );
   gpc1_1 gpc1472 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc1473 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc1474 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc1475 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1476 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1477 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1478 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc1479 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc1480 (
      {stage0_10[475]},
      {stage1_10[177]}
   );
   gpc1_1 gpc1481 (
      {stage0_10[476]},
      {stage1_10[178]}
   );
   gpc1_1 gpc1482 (
      {stage0_10[477]},
      {stage1_10[179]}
   );
   gpc1_1 gpc1483 (
      {stage0_10[478]},
      {stage1_10[180]}
   );
   gpc1_1 gpc1484 (
      {stage0_10[479]},
      {stage1_10[181]}
   );
   gpc1_1 gpc1485 (
      {stage0_10[480]},
      {stage1_10[182]}
   );
   gpc1_1 gpc1486 (
      {stage0_10[481]},
      {stage1_10[183]}
   );
   gpc1_1 gpc1487 (
      {stage0_10[482]},
      {stage1_10[184]}
   );
   gpc1_1 gpc1488 (
      {stage0_10[483]},
      {stage1_10[185]}
   );
   gpc1_1 gpc1489 (
      {stage0_10[484]},
      {stage1_10[186]}
   );
   gpc1_1 gpc1490 (
      {stage0_10[485]},
      {stage1_10[187]}
   );
   gpc1_1 gpc1491 (
      {stage0_11[451]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1492 (
      {stage0_11[452]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1493 (
      {stage0_11[453]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1494 (
      {stage0_11[454]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1495 (
      {stage0_11[455]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1496 (
      {stage0_11[456]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1497 (
      {stage0_11[457]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1498 (
      {stage0_11[458]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1499 (
      {stage0_11[459]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1500 (
      {stage0_11[460]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1501 (
      {stage0_11[461]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1502 (
      {stage0_11[462]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1503 (
      {stage0_11[463]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1504 (
      {stage0_11[464]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1505 (
      {stage0_11[465]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1506 (
      {stage0_11[466]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1507 (
      {stage0_11[467]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1508 (
      {stage0_11[468]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1509 (
      {stage0_11[469]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1510 (
      {stage0_11[470]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1511 (
      {stage0_11[471]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1512 (
      {stage0_11[472]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1513 (
      {stage0_11[473]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1514 (
      {stage0_11[474]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1515 (
      {stage0_11[475]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1516 (
      {stage0_11[476]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1517 (
      {stage0_11[477]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1518 (
      {stage0_11[478]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1519 (
      {stage0_11[479]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1520 (
      {stage0_11[480]},
      {stage1_11[214]}
   );
   gpc1_1 gpc1521 (
      {stage0_11[481]},
      {stage1_11[215]}
   );
   gpc1_1 gpc1522 (
      {stage0_11[482]},
      {stage1_11[216]}
   );
   gpc1_1 gpc1523 (
      {stage0_11[483]},
      {stage1_11[217]}
   );
   gpc1_1 gpc1524 (
      {stage0_11[484]},
      {stage1_11[218]}
   );
   gpc1_1 gpc1525 (
      {stage0_11[485]},
      {stage1_11[219]}
   );
   gpc1_1 gpc1526 (
      {stage0_12[408]},
      {stage1_12[204]}
   );
   gpc1_1 gpc1527 (
      {stage0_12[409]},
      {stage1_12[205]}
   );
   gpc1_1 gpc1528 (
      {stage0_12[410]},
      {stage1_12[206]}
   );
   gpc1_1 gpc1529 (
      {stage0_12[411]},
      {stage1_12[207]}
   );
   gpc1_1 gpc1530 (
      {stage0_12[412]},
      {stage1_12[208]}
   );
   gpc1_1 gpc1531 (
      {stage0_12[413]},
      {stage1_12[209]}
   );
   gpc1_1 gpc1532 (
      {stage0_12[414]},
      {stage1_12[210]}
   );
   gpc1_1 gpc1533 (
      {stage0_12[415]},
      {stage1_12[211]}
   );
   gpc1_1 gpc1534 (
      {stage0_12[416]},
      {stage1_12[212]}
   );
   gpc1_1 gpc1535 (
      {stage0_12[417]},
      {stage1_12[213]}
   );
   gpc1_1 gpc1536 (
      {stage0_12[418]},
      {stage1_12[214]}
   );
   gpc1_1 gpc1537 (
      {stage0_12[419]},
      {stage1_12[215]}
   );
   gpc1_1 gpc1538 (
      {stage0_12[420]},
      {stage1_12[216]}
   );
   gpc1_1 gpc1539 (
      {stage0_12[421]},
      {stage1_12[217]}
   );
   gpc1_1 gpc1540 (
      {stage0_12[422]},
      {stage1_12[218]}
   );
   gpc1_1 gpc1541 (
      {stage0_12[423]},
      {stage1_12[219]}
   );
   gpc1_1 gpc1542 (
      {stage0_12[424]},
      {stage1_12[220]}
   );
   gpc1_1 gpc1543 (
      {stage0_12[425]},
      {stage1_12[221]}
   );
   gpc1_1 gpc1544 (
      {stage0_12[426]},
      {stage1_12[222]}
   );
   gpc1_1 gpc1545 (
      {stage0_12[427]},
      {stage1_12[223]}
   );
   gpc1_1 gpc1546 (
      {stage0_12[428]},
      {stage1_12[224]}
   );
   gpc1_1 gpc1547 (
      {stage0_12[429]},
      {stage1_12[225]}
   );
   gpc1_1 gpc1548 (
      {stage0_12[430]},
      {stage1_12[226]}
   );
   gpc1_1 gpc1549 (
      {stage0_12[431]},
      {stage1_12[227]}
   );
   gpc1_1 gpc1550 (
      {stage0_12[432]},
      {stage1_12[228]}
   );
   gpc1_1 gpc1551 (
      {stage0_12[433]},
      {stage1_12[229]}
   );
   gpc1_1 gpc1552 (
      {stage0_12[434]},
      {stage1_12[230]}
   );
   gpc1_1 gpc1553 (
      {stage0_12[435]},
      {stage1_12[231]}
   );
   gpc1_1 gpc1554 (
      {stage0_12[436]},
      {stage1_12[232]}
   );
   gpc1_1 gpc1555 (
      {stage0_12[437]},
      {stage1_12[233]}
   );
   gpc1_1 gpc1556 (
      {stage0_12[438]},
      {stage1_12[234]}
   );
   gpc1_1 gpc1557 (
      {stage0_12[439]},
      {stage1_12[235]}
   );
   gpc1_1 gpc1558 (
      {stage0_12[440]},
      {stage1_12[236]}
   );
   gpc1_1 gpc1559 (
      {stage0_12[441]},
      {stage1_12[237]}
   );
   gpc1_1 gpc1560 (
      {stage0_12[442]},
      {stage1_12[238]}
   );
   gpc1_1 gpc1561 (
      {stage0_12[443]},
      {stage1_12[239]}
   );
   gpc1_1 gpc1562 (
      {stage0_12[444]},
      {stage1_12[240]}
   );
   gpc1_1 gpc1563 (
      {stage0_12[445]},
      {stage1_12[241]}
   );
   gpc1_1 gpc1564 (
      {stage0_12[446]},
      {stage1_12[242]}
   );
   gpc1_1 gpc1565 (
      {stage0_12[447]},
      {stage1_12[243]}
   );
   gpc1_1 gpc1566 (
      {stage0_12[448]},
      {stage1_12[244]}
   );
   gpc1_1 gpc1567 (
      {stage0_12[449]},
      {stage1_12[245]}
   );
   gpc1_1 gpc1568 (
      {stage0_12[450]},
      {stage1_12[246]}
   );
   gpc1_1 gpc1569 (
      {stage0_12[451]},
      {stage1_12[247]}
   );
   gpc1_1 gpc1570 (
      {stage0_12[452]},
      {stage1_12[248]}
   );
   gpc1_1 gpc1571 (
      {stage0_12[453]},
      {stage1_12[249]}
   );
   gpc1_1 gpc1572 (
      {stage0_12[454]},
      {stage1_12[250]}
   );
   gpc1_1 gpc1573 (
      {stage0_12[455]},
      {stage1_12[251]}
   );
   gpc1_1 gpc1574 (
      {stage0_12[456]},
      {stage1_12[252]}
   );
   gpc1_1 gpc1575 (
      {stage0_12[457]},
      {stage1_12[253]}
   );
   gpc1_1 gpc1576 (
      {stage0_12[458]},
      {stage1_12[254]}
   );
   gpc1_1 gpc1577 (
      {stage0_12[459]},
      {stage1_12[255]}
   );
   gpc1_1 gpc1578 (
      {stage0_12[460]},
      {stage1_12[256]}
   );
   gpc1_1 gpc1579 (
      {stage0_12[461]},
      {stage1_12[257]}
   );
   gpc1_1 gpc1580 (
      {stage0_12[462]},
      {stage1_12[258]}
   );
   gpc1_1 gpc1581 (
      {stage0_12[463]},
      {stage1_12[259]}
   );
   gpc1_1 gpc1582 (
      {stage0_12[464]},
      {stage1_12[260]}
   );
   gpc1_1 gpc1583 (
      {stage0_12[465]},
      {stage1_12[261]}
   );
   gpc1_1 gpc1584 (
      {stage0_12[466]},
      {stage1_12[262]}
   );
   gpc1_1 gpc1585 (
      {stage0_12[467]},
      {stage1_12[263]}
   );
   gpc1_1 gpc1586 (
      {stage0_12[468]},
      {stage1_12[264]}
   );
   gpc1_1 gpc1587 (
      {stage0_12[469]},
      {stage1_12[265]}
   );
   gpc1_1 gpc1588 (
      {stage0_12[470]},
      {stage1_12[266]}
   );
   gpc1_1 gpc1589 (
      {stage0_12[471]},
      {stage1_12[267]}
   );
   gpc1_1 gpc1590 (
      {stage0_12[472]},
      {stage1_12[268]}
   );
   gpc1_1 gpc1591 (
      {stage0_12[473]},
      {stage1_12[269]}
   );
   gpc1_1 gpc1592 (
      {stage0_12[474]},
      {stage1_12[270]}
   );
   gpc1_1 gpc1593 (
      {stage0_12[475]},
      {stage1_12[271]}
   );
   gpc1_1 gpc1594 (
      {stage0_12[476]},
      {stage1_12[272]}
   );
   gpc1_1 gpc1595 (
      {stage0_12[477]},
      {stage1_12[273]}
   );
   gpc1_1 gpc1596 (
      {stage0_12[478]},
      {stage1_12[274]}
   );
   gpc1_1 gpc1597 (
      {stage0_12[479]},
      {stage1_12[275]}
   );
   gpc1_1 gpc1598 (
      {stage0_12[480]},
      {stage1_12[276]}
   );
   gpc1_1 gpc1599 (
      {stage0_12[481]},
      {stage1_12[277]}
   );
   gpc1_1 gpc1600 (
      {stage0_12[482]},
      {stage1_12[278]}
   );
   gpc1_1 gpc1601 (
      {stage0_12[483]},
      {stage1_12[279]}
   );
   gpc1_1 gpc1602 (
      {stage0_12[484]},
      {stage1_12[280]}
   );
   gpc1_1 gpc1603 (
      {stage0_12[485]},
      {stage1_12[281]}
   );
   gpc1_1 gpc1604 (
      {stage0_13[476]},
      {stage1_13[195]}
   );
   gpc1_1 gpc1605 (
      {stage0_13[477]},
      {stage1_13[196]}
   );
   gpc1_1 gpc1606 (
      {stage0_13[478]},
      {stage1_13[197]}
   );
   gpc1_1 gpc1607 (
      {stage0_13[479]},
      {stage1_13[198]}
   );
   gpc1_1 gpc1608 (
      {stage0_13[480]},
      {stage1_13[199]}
   );
   gpc1_1 gpc1609 (
      {stage0_13[481]},
      {stage1_13[200]}
   );
   gpc1_1 gpc1610 (
      {stage0_13[482]},
      {stage1_13[201]}
   );
   gpc1_1 gpc1611 (
      {stage0_13[483]},
      {stage1_13[202]}
   );
   gpc1_1 gpc1612 (
      {stage0_13[484]},
      {stage1_13[203]}
   );
   gpc1_1 gpc1613 (
      {stage0_13[485]},
      {stage1_13[204]}
   );
   gpc1_1 gpc1614 (
      {stage0_14[349]},
      {stage1_14[160]}
   );
   gpc1_1 gpc1615 (
      {stage0_14[350]},
      {stage1_14[161]}
   );
   gpc1_1 gpc1616 (
      {stage0_14[351]},
      {stage1_14[162]}
   );
   gpc1_1 gpc1617 (
      {stage0_14[352]},
      {stage1_14[163]}
   );
   gpc1_1 gpc1618 (
      {stage0_14[353]},
      {stage1_14[164]}
   );
   gpc1_1 gpc1619 (
      {stage0_14[354]},
      {stage1_14[165]}
   );
   gpc1_1 gpc1620 (
      {stage0_14[355]},
      {stage1_14[166]}
   );
   gpc1_1 gpc1621 (
      {stage0_14[356]},
      {stage1_14[167]}
   );
   gpc1_1 gpc1622 (
      {stage0_14[357]},
      {stage1_14[168]}
   );
   gpc1_1 gpc1623 (
      {stage0_14[358]},
      {stage1_14[169]}
   );
   gpc1_1 gpc1624 (
      {stage0_14[359]},
      {stage1_14[170]}
   );
   gpc1_1 gpc1625 (
      {stage0_14[360]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1626 (
      {stage0_14[361]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1627 (
      {stage0_14[362]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1628 (
      {stage0_14[363]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1629 (
      {stage0_14[364]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1630 (
      {stage0_14[365]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1631 (
      {stage0_14[366]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1632 (
      {stage0_14[367]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1633 (
      {stage0_14[368]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1634 (
      {stage0_14[369]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1635 (
      {stage0_14[370]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1636 (
      {stage0_14[371]},
      {stage1_14[182]}
   );
   gpc1_1 gpc1637 (
      {stage0_14[372]},
      {stage1_14[183]}
   );
   gpc1_1 gpc1638 (
      {stage0_14[373]},
      {stage1_14[184]}
   );
   gpc1_1 gpc1639 (
      {stage0_14[374]},
      {stage1_14[185]}
   );
   gpc1_1 gpc1640 (
      {stage0_14[375]},
      {stage1_14[186]}
   );
   gpc1_1 gpc1641 (
      {stage0_14[376]},
      {stage1_14[187]}
   );
   gpc1_1 gpc1642 (
      {stage0_14[377]},
      {stage1_14[188]}
   );
   gpc1_1 gpc1643 (
      {stage0_14[378]},
      {stage1_14[189]}
   );
   gpc1_1 gpc1644 (
      {stage0_14[379]},
      {stage1_14[190]}
   );
   gpc1_1 gpc1645 (
      {stage0_14[380]},
      {stage1_14[191]}
   );
   gpc1_1 gpc1646 (
      {stage0_14[381]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1647 (
      {stage0_14[382]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1648 (
      {stage0_14[383]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1649 (
      {stage0_14[384]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1650 (
      {stage0_14[385]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1651 (
      {stage0_14[386]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1652 (
      {stage0_14[387]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1653 (
      {stage0_14[388]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1654 (
      {stage0_14[389]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1655 (
      {stage0_14[390]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1656 (
      {stage0_14[391]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1657 (
      {stage0_14[392]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1658 (
      {stage0_14[393]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1659 (
      {stage0_14[394]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1660 (
      {stage0_14[395]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1661 (
      {stage0_14[396]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1662 (
      {stage0_14[397]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1663 (
      {stage0_14[398]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1664 (
      {stage0_14[399]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1665 (
      {stage0_14[400]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1666 (
      {stage0_14[401]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1667 (
      {stage0_14[402]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1668 (
      {stage0_14[403]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1669 (
      {stage0_14[404]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1670 (
      {stage0_14[405]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1671 (
      {stage0_14[406]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1672 (
      {stage0_14[407]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1673 (
      {stage0_14[408]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1674 (
      {stage0_14[409]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1675 (
      {stage0_14[410]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1676 (
      {stage0_14[411]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1677 (
      {stage0_14[412]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1678 (
      {stage0_14[413]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1679 (
      {stage0_14[414]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1680 (
      {stage0_14[415]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1681 (
      {stage0_14[416]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1682 (
      {stage0_14[417]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1683 (
      {stage0_14[418]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1684 (
      {stage0_14[419]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1685 (
      {stage0_14[420]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1686 (
      {stage0_14[421]},
      {stage1_14[232]}
   );
   gpc1_1 gpc1687 (
      {stage0_14[422]},
      {stage1_14[233]}
   );
   gpc1_1 gpc1688 (
      {stage0_14[423]},
      {stage1_14[234]}
   );
   gpc1_1 gpc1689 (
      {stage0_14[424]},
      {stage1_14[235]}
   );
   gpc1_1 gpc1690 (
      {stage0_14[425]},
      {stage1_14[236]}
   );
   gpc1_1 gpc1691 (
      {stage0_14[426]},
      {stage1_14[237]}
   );
   gpc1_1 gpc1692 (
      {stage0_14[427]},
      {stage1_14[238]}
   );
   gpc1_1 gpc1693 (
      {stage0_14[428]},
      {stage1_14[239]}
   );
   gpc1_1 gpc1694 (
      {stage0_14[429]},
      {stage1_14[240]}
   );
   gpc1_1 gpc1695 (
      {stage0_14[430]},
      {stage1_14[241]}
   );
   gpc1_1 gpc1696 (
      {stage0_14[431]},
      {stage1_14[242]}
   );
   gpc1_1 gpc1697 (
      {stage0_14[432]},
      {stage1_14[243]}
   );
   gpc1_1 gpc1698 (
      {stage0_14[433]},
      {stage1_14[244]}
   );
   gpc1_1 gpc1699 (
      {stage0_14[434]},
      {stage1_14[245]}
   );
   gpc1_1 gpc1700 (
      {stage0_14[435]},
      {stage1_14[246]}
   );
   gpc1_1 gpc1701 (
      {stage0_14[436]},
      {stage1_14[247]}
   );
   gpc1_1 gpc1702 (
      {stage0_14[437]},
      {stage1_14[248]}
   );
   gpc1_1 gpc1703 (
      {stage0_14[438]},
      {stage1_14[249]}
   );
   gpc1_1 gpc1704 (
      {stage0_14[439]},
      {stage1_14[250]}
   );
   gpc1_1 gpc1705 (
      {stage0_14[440]},
      {stage1_14[251]}
   );
   gpc1_1 gpc1706 (
      {stage0_14[441]},
      {stage1_14[252]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[442]},
      {stage1_14[253]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[443]},
      {stage1_14[254]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[444]},
      {stage1_14[255]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[445]},
      {stage1_14[256]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[446]},
      {stage1_14[257]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[447]},
      {stage1_14[258]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[448]},
      {stage1_14[259]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[449]},
      {stage1_14[260]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[450]},
      {stage1_14[261]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[451]},
      {stage1_14[262]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[452]},
      {stage1_14[263]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[453]},
      {stage1_14[264]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[454]},
      {stage1_14[265]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[455]},
      {stage1_14[266]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[456]},
      {stage1_14[267]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[457]},
      {stage1_14[268]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[458]},
      {stage1_14[269]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[459]},
      {stage1_14[270]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[460]},
      {stage1_14[271]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[461]},
      {stage1_14[272]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[462]},
      {stage1_14[273]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[463]},
      {stage1_14[274]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[464]},
      {stage1_14[275]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[465]},
      {stage1_14[276]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[466]},
      {stage1_14[277]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[467]},
      {stage1_14[278]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[468]},
      {stage1_14[279]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[469]},
      {stage1_14[280]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[470]},
      {stage1_14[281]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[471]},
      {stage1_14[282]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[472]},
      {stage1_14[283]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[473]},
      {stage1_14[284]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[474]},
      {stage1_14[285]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[475]},
      {stage1_14[286]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[476]},
      {stage1_14[287]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[477]},
      {stage1_14[288]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[478]},
      {stage1_14[289]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[479]},
      {stage1_14[290]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[480]},
      {stage1_14[291]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[481]},
      {stage1_14[292]}
   );
   gpc1_1 gpc1747 (
      {stage0_14[482]},
      {stage1_14[293]}
   );
   gpc1_1 gpc1748 (
      {stage0_14[483]},
      {stage1_14[294]}
   );
   gpc1_1 gpc1749 (
      {stage0_14[484]},
      {stage1_14[295]}
   );
   gpc1_1 gpc1750 (
      {stage0_14[485]},
      {stage1_14[296]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[480]},
      {stage1_15[166]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[481]},
      {stage1_15[167]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[482]},
      {stage1_15[168]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[483]},
      {stage1_15[169]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[484]},
      {stage1_15[170]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[485]},
      {stage1_15[171]}
   );
   gpc1_1 gpc1757 (
      {stage0_16[411]},
      {stage1_16[190]}
   );
   gpc1_1 gpc1758 (
      {stage0_16[412]},
      {stage1_16[191]}
   );
   gpc1_1 gpc1759 (
      {stage0_16[413]},
      {stage1_16[192]}
   );
   gpc1_1 gpc1760 (
      {stage0_16[414]},
      {stage1_16[193]}
   );
   gpc1_1 gpc1761 (
      {stage0_16[415]},
      {stage1_16[194]}
   );
   gpc1_1 gpc1762 (
      {stage0_16[416]},
      {stage1_16[195]}
   );
   gpc1_1 gpc1763 (
      {stage0_16[417]},
      {stage1_16[196]}
   );
   gpc1_1 gpc1764 (
      {stage0_16[418]},
      {stage1_16[197]}
   );
   gpc1_1 gpc1765 (
      {stage0_16[419]},
      {stage1_16[198]}
   );
   gpc1_1 gpc1766 (
      {stage0_16[420]},
      {stage1_16[199]}
   );
   gpc1_1 gpc1767 (
      {stage0_16[421]},
      {stage1_16[200]}
   );
   gpc1_1 gpc1768 (
      {stage0_16[422]},
      {stage1_16[201]}
   );
   gpc1_1 gpc1769 (
      {stage0_16[423]},
      {stage1_16[202]}
   );
   gpc1_1 gpc1770 (
      {stage0_16[424]},
      {stage1_16[203]}
   );
   gpc1_1 gpc1771 (
      {stage0_16[425]},
      {stage1_16[204]}
   );
   gpc1_1 gpc1772 (
      {stage0_16[426]},
      {stage1_16[205]}
   );
   gpc1_1 gpc1773 (
      {stage0_16[427]},
      {stage1_16[206]}
   );
   gpc1_1 gpc1774 (
      {stage0_16[428]},
      {stage1_16[207]}
   );
   gpc1_1 gpc1775 (
      {stage0_16[429]},
      {stage1_16[208]}
   );
   gpc1_1 gpc1776 (
      {stage0_16[430]},
      {stage1_16[209]}
   );
   gpc1_1 gpc1777 (
      {stage0_16[431]},
      {stage1_16[210]}
   );
   gpc1_1 gpc1778 (
      {stage0_16[432]},
      {stage1_16[211]}
   );
   gpc1_1 gpc1779 (
      {stage0_16[433]},
      {stage1_16[212]}
   );
   gpc1_1 gpc1780 (
      {stage0_16[434]},
      {stage1_16[213]}
   );
   gpc1_1 gpc1781 (
      {stage0_16[435]},
      {stage1_16[214]}
   );
   gpc1_1 gpc1782 (
      {stage0_16[436]},
      {stage1_16[215]}
   );
   gpc1_1 gpc1783 (
      {stage0_16[437]},
      {stage1_16[216]}
   );
   gpc1_1 gpc1784 (
      {stage0_16[438]},
      {stage1_16[217]}
   );
   gpc1_1 gpc1785 (
      {stage0_16[439]},
      {stage1_16[218]}
   );
   gpc1_1 gpc1786 (
      {stage0_16[440]},
      {stage1_16[219]}
   );
   gpc1_1 gpc1787 (
      {stage0_16[441]},
      {stage1_16[220]}
   );
   gpc1_1 gpc1788 (
      {stage0_16[442]},
      {stage1_16[221]}
   );
   gpc1_1 gpc1789 (
      {stage0_16[443]},
      {stage1_16[222]}
   );
   gpc1_1 gpc1790 (
      {stage0_16[444]},
      {stage1_16[223]}
   );
   gpc1_1 gpc1791 (
      {stage0_16[445]},
      {stage1_16[224]}
   );
   gpc1_1 gpc1792 (
      {stage0_16[446]},
      {stage1_16[225]}
   );
   gpc1_1 gpc1793 (
      {stage0_16[447]},
      {stage1_16[226]}
   );
   gpc1_1 gpc1794 (
      {stage0_16[448]},
      {stage1_16[227]}
   );
   gpc1_1 gpc1795 (
      {stage0_16[449]},
      {stage1_16[228]}
   );
   gpc1_1 gpc1796 (
      {stage0_16[450]},
      {stage1_16[229]}
   );
   gpc1_1 gpc1797 (
      {stage0_16[451]},
      {stage1_16[230]}
   );
   gpc1_1 gpc1798 (
      {stage0_16[452]},
      {stage1_16[231]}
   );
   gpc1_1 gpc1799 (
      {stage0_16[453]},
      {stage1_16[232]}
   );
   gpc1_1 gpc1800 (
      {stage0_16[454]},
      {stage1_16[233]}
   );
   gpc1_1 gpc1801 (
      {stage0_16[455]},
      {stage1_16[234]}
   );
   gpc1_1 gpc1802 (
      {stage0_16[456]},
      {stage1_16[235]}
   );
   gpc1_1 gpc1803 (
      {stage0_16[457]},
      {stage1_16[236]}
   );
   gpc1_1 gpc1804 (
      {stage0_16[458]},
      {stage1_16[237]}
   );
   gpc1_1 gpc1805 (
      {stage0_16[459]},
      {stage1_16[238]}
   );
   gpc1_1 gpc1806 (
      {stage0_16[460]},
      {stage1_16[239]}
   );
   gpc1_1 gpc1807 (
      {stage0_16[461]},
      {stage1_16[240]}
   );
   gpc1_1 gpc1808 (
      {stage0_16[462]},
      {stage1_16[241]}
   );
   gpc1_1 gpc1809 (
      {stage0_16[463]},
      {stage1_16[242]}
   );
   gpc1_1 gpc1810 (
      {stage0_16[464]},
      {stage1_16[243]}
   );
   gpc1_1 gpc1811 (
      {stage0_16[465]},
      {stage1_16[244]}
   );
   gpc1_1 gpc1812 (
      {stage0_16[466]},
      {stage1_16[245]}
   );
   gpc1_1 gpc1813 (
      {stage0_16[467]},
      {stage1_16[246]}
   );
   gpc1_1 gpc1814 (
      {stage0_16[468]},
      {stage1_16[247]}
   );
   gpc1_1 gpc1815 (
      {stage0_16[469]},
      {stage1_16[248]}
   );
   gpc1_1 gpc1816 (
      {stage0_16[470]},
      {stage1_16[249]}
   );
   gpc1_1 gpc1817 (
      {stage0_16[471]},
      {stage1_16[250]}
   );
   gpc1_1 gpc1818 (
      {stage0_16[472]},
      {stage1_16[251]}
   );
   gpc1_1 gpc1819 (
      {stage0_16[473]},
      {stage1_16[252]}
   );
   gpc1_1 gpc1820 (
      {stage0_16[474]},
      {stage1_16[253]}
   );
   gpc1_1 gpc1821 (
      {stage0_16[475]},
      {stage1_16[254]}
   );
   gpc1_1 gpc1822 (
      {stage0_16[476]},
      {stage1_16[255]}
   );
   gpc1_1 gpc1823 (
      {stage0_16[477]},
      {stage1_16[256]}
   );
   gpc1_1 gpc1824 (
      {stage0_16[478]},
      {stage1_16[257]}
   );
   gpc1_1 gpc1825 (
      {stage0_16[479]},
      {stage1_16[258]}
   );
   gpc1_1 gpc1826 (
      {stage0_16[480]},
      {stage1_16[259]}
   );
   gpc1_1 gpc1827 (
      {stage0_16[481]},
      {stage1_16[260]}
   );
   gpc1_1 gpc1828 (
      {stage0_16[482]},
      {stage1_16[261]}
   );
   gpc1_1 gpc1829 (
      {stage0_16[483]},
      {stage1_16[262]}
   );
   gpc1_1 gpc1830 (
      {stage0_16[484]},
      {stage1_16[263]}
   );
   gpc1_1 gpc1831 (
      {stage0_16[485]},
      {stage1_16[264]}
   );
   gpc1_1 gpc1832 (
      {stage0_17[402]},
      {stage1_17[187]}
   );
   gpc1_1 gpc1833 (
      {stage0_17[403]},
      {stage1_17[188]}
   );
   gpc1_1 gpc1834 (
      {stage0_17[404]},
      {stage1_17[189]}
   );
   gpc1_1 gpc1835 (
      {stage0_17[405]},
      {stage1_17[190]}
   );
   gpc1_1 gpc1836 (
      {stage0_17[406]},
      {stage1_17[191]}
   );
   gpc1_1 gpc1837 (
      {stage0_17[407]},
      {stage1_17[192]}
   );
   gpc1_1 gpc1838 (
      {stage0_17[408]},
      {stage1_17[193]}
   );
   gpc1_1 gpc1839 (
      {stage0_17[409]},
      {stage1_17[194]}
   );
   gpc1_1 gpc1840 (
      {stage0_17[410]},
      {stage1_17[195]}
   );
   gpc1_1 gpc1841 (
      {stage0_17[411]},
      {stage1_17[196]}
   );
   gpc1_1 gpc1842 (
      {stage0_17[412]},
      {stage1_17[197]}
   );
   gpc1_1 gpc1843 (
      {stage0_17[413]},
      {stage1_17[198]}
   );
   gpc1_1 gpc1844 (
      {stage0_17[414]},
      {stage1_17[199]}
   );
   gpc1_1 gpc1845 (
      {stage0_17[415]},
      {stage1_17[200]}
   );
   gpc1_1 gpc1846 (
      {stage0_17[416]},
      {stage1_17[201]}
   );
   gpc1_1 gpc1847 (
      {stage0_17[417]},
      {stage1_17[202]}
   );
   gpc1_1 gpc1848 (
      {stage0_17[418]},
      {stage1_17[203]}
   );
   gpc1_1 gpc1849 (
      {stage0_17[419]},
      {stage1_17[204]}
   );
   gpc1_1 gpc1850 (
      {stage0_17[420]},
      {stage1_17[205]}
   );
   gpc1_1 gpc1851 (
      {stage0_17[421]},
      {stage1_17[206]}
   );
   gpc1_1 gpc1852 (
      {stage0_17[422]},
      {stage1_17[207]}
   );
   gpc1_1 gpc1853 (
      {stage0_17[423]},
      {stage1_17[208]}
   );
   gpc1_1 gpc1854 (
      {stage0_17[424]},
      {stage1_17[209]}
   );
   gpc1_1 gpc1855 (
      {stage0_17[425]},
      {stage1_17[210]}
   );
   gpc1_1 gpc1856 (
      {stage0_17[426]},
      {stage1_17[211]}
   );
   gpc1_1 gpc1857 (
      {stage0_17[427]},
      {stage1_17[212]}
   );
   gpc1_1 gpc1858 (
      {stage0_17[428]},
      {stage1_17[213]}
   );
   gpc1_1 gpc1859 (
      {stage0_17[429]},
      {stage1_17[214]}
   );
   gpc1_1 gpc1860 (
      {stage0_17[430]},
      {stage1_17[215]}
   );
   gpc1_1 gpc1861 (
      {stage0_17[431]},
      {stage1_17[216]}
   );
   gpc1_1 gpc1862 (
      {stage0_17[432]},
      {stage1_17[217]}
   );
   gpc1_1 gpc1863 (
      {stage0_17[433]},
      {stage1_17[218]}
   );
   gpc1_1 gpc1864 (
      {stage0_17[434]},
      {stage1_17[219]}
   );
   gpc1_1 gpc1865 (
      {stage0_17[435]},
      {stage1_17[220]}
   );
   gpc1_1 gpc1866 (
      {stage0_17[436]},
      {stage1_17[221]}
   );
   gpc1_1 gpc1867 (
      {stage0_17[437]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1868 (
      {stage0_17[438]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1869 (
      {stage0_17[439]},
      {stage1_17[224]}
   );
   gpc1_1 gpc1870 (
      {stage0_17[440]},
      {stage1_17[225]}
   );
   gpc1_1 gpc1871 (
      {stage0_17[441]},
      {stage1_17[226]}
   );
   gpc1_1 gpc1872 (
      {stage0_17[442]},
      {stage1_17[227]}
   );
   gpc1_1 gpc1873 (
      {stage0_17[443]},
      {stage1_17[228]}
   );
   gpc1_1 gpc1874 (
      {stage0_17[444]},
      {stage1_17[229]}
   );
   gpc1_1 gpc1875 (
      {stage0_17[445]},
      {stage1_17[230]}
   );
   gpc1_1 gpc1876 (
      {stage0_17[446]},
      {stage1_17[231]}
   );
   gpc1_1 gpc1877 (
      {stage0_17[447]},
      {stage1_17[232]}
   );
   gpc1_1 gpc1878 (
      {stage0_17[448]},
      {stage1_17[233]}
   );
   gpc1_1 gpc1879 (
      {stage0_17[449]},
      {stage1_17[234]}
   );
   gpc1_1 gpc1880 (
      {stage0_17[450]},
      {stage1_17[235]}
   );
   gpc1_1 gpc1881 (
      {stage0_17[451]},
      {stage1_17[236]}
   );
   gpc1_1 gpc1882 (
      {stage0_17[452]},
      {stage1_17[237]}
   );
   gpc1_1 gpc1883 (
      {stage0_17[453]},
      {stage1_17[238]}
   );
   gpc1_1 gpc1884 (
      {stage0_17[454]},
      {stage1_17[239]}
   );
   gpc1_1 gpc1885 (
      {stage0_17[455]},
      {stage1_17[240]}
   );
   gpc1_1 gpc1886 (
      {stage0_17[456]},
      {stage1_17[241]}
   );
   gpc1_1 gpc1887 (
      {stage0_17[457]},
      {stage1_17[242]}
   );
   gpc1_1 gpc1888 (
      {stage0_17[458]},
      {stage1_17[243]}
   );
   gpc1_1 gpc1889 (
      {stage0_17[459]},
      {stage1_17[244]}
   );
   gpc1_1 gpc1890 (
      {stage0_17[460]},
      {stage1_17[245]}
   );
   gpc1_1 gpc1891 (
      {stage0_17[461]},
      {stage1_17[246]}
   );
   gpc1_1 gpc1892 (
      {stage0_17[462]},
      {stage1_17[247]}
   );
   gpc1_1 gpc1893 (
      {stage0_17[463]},
      {stage1_17[248]}
   );
   gpc1_1 gpc1894 (
      {stage0_17[464]},
      {stage1_17[249]}
   );
   gpc1_1 gpc1895 (
      {stage0_17[465]},
      {stage1_17[250]}
   );
   gpc1_1 gpc1896 (
      {stage0_17[466]},
      {stage1_17[251]}
   );
   gpc1_1 gpc1897 (
      {stage0_17[467]},
      {stage1_17[252]}
   );
   gpc1_1 gpc1898 (
      {stage0_17[468]},
      {stage1_17[253]}
   );
   gpc1_1 gpc1899 (
      {stage0_17[469]},
      {stage1_17[254]}
   );
   gpc1_1 gpc1900 (
      {stage0_17[470]},
      {stage1_17[255]}
   );
   gpc1_1 gpc1901 (
      {stage0_17[471]},
      {stage1_17[256]}
   );
   gpc1_1 gpc1902 (
      {stage0_17[472]},
      {stage1_17[257]}
   );
   gpc1_1 gpc1903 (
      {stage0_17[473]},
      {stage1_17[258]}
   );
   gpc1_1 gpc1904 (
      {stage0_17[474]},
      {stage1_17[259]}
   );
   gpc1_1 gpc1905 (
      {stage0_17[475]},
      {stage1_17[260]}
   );
   gpc1_1 gpc1906 (
      {stage0_17[476]},
      {stage1_17[261]}
   );
   gpc1_1 gpc1907 (
      {stage0_17[477]},
      {stage1_17[262]}
   );
   gpc1_1 gpc1908 (
      {stage0_17[478]},
      {stage1_17[263]}
   );
   gpc1_1 gpc1909 (
      {stage0_17[479]},
      {stage1_17[264]}
   );
   gpc1_1 gpc1910 (
      {stage0_17[480]},
      {stage1_17[265]}
   );
   gpc1_1 gpc1911 (
      {stage0_17[481]},
      {stage1_17[266]}
   );
   gpc1_1 gpc1912 (
      {stage0_17[482]},
      {stage1_17[267]}
   );
   gpc1_1 gpc1913 (
      {stage0_17[483]},
      {stage1_17[268]}
   );
   gpc1_1 gpc1914 (
      {stage0_17[484]},
      {stage1_17[269]}
   );
   gpc1_1 gpc1915 (
      {stage0_17[485]},
      {stage1_17[270]}
   );
   gpc1_1 gpc1916 (
      {stage0_18[447]},
      {stage1_18[162]}
   );
   gpc1_1 gpc1917 (
      {stage0_18[448]},
      {stage1_18[163]}
   );
   gpc1_1 gpc1918 (
      {stage0_18[449]},
      {stage1_18[164]}
   );
   gpc1_1 gpc1919 (
      {stage0_18[450]},
      {stage1_18[165]}
   );
   gpc1_1 gpc1920 (
      {stage0_18[451]},
      {stage1_18[166]}
   );
   gpc1_1 gpc1921 (
      {stage0_18[452]},
      {stage1_18[167]}
   );
   gpc1_1 gpc1922 (
      {stage0_18[453]},
      {stage1_18[168]}
   );
   gpc1_1 gpc1923 (
      {stage0_18[454]},
      {stage1_18[169]}
   );
   gpc1_1 gpc1924 (
      {stage0_18[455]},
      {stage1_18[170]}
   );
   gpc1_1 gpc1925 (
      {stage0_18[456]},
      {stage1_18[171]}
   );
   gpc1_1 gpc1926 (
      {stage0_18[457]},
      {stage1_18[172]}
   );
   gpc1_1 gpc1927 (
      {stage0_18[458]},
      {stage1_18[173]}
   );
   gpc1_1 gpc1928 (
      {stage0_18[459]},
      {stage1_18[174]}
   );
   gpc1_1 gpc1929 (
      {stage0_18[460]},
      {stage1_18[175]}
   );
   gpc1_1 gpc1930 (
      {stage0_18[461]},
      {stage1_18[176]}
   );
   gpc1_1 gpc1931 (
      {stage0_18[462]},
      {stage1_18[177]}
   );
   gpc1_1 gpc1932 (
      {stage0_18[463]},
      {stage1_18[178]}
   );
   gpc1_1 gpc1933 (
      {stage0_18[464]},
      {stage1_18[179]}
   );
   gpc1_1 gpc1934 (
      {stage0_18[465]},
      {stage1_18[180]}
   );
   gpc1_1 gpc1935 (
      {stage0_18[466]},
      {stage1_18[181]}
   );
   gpc1_1 gpc1936 (
      {stage0_18[467]},
      {stage1_18[182]}
   );
   gpc1_1 gpc1937 (
      {stage0_18[468]},
      {stage1_18[183]}
   );
   gpc1_1 gpc1938 (
      {stage0_18[469]},
      {stage1_18[184]}
   );
   gpc1_1 gpc1939 (
      {stage0_18[470]},
      {stage1_18[185]}
   );
   gpc1_1 gpc1940 (
      {stage0_18[471]},
      {stage1_18[186]}
   );
   gpc1_1 gpc1941 (
      {stage0_18[472]},
      {stage1_18[187]}
   );
   gpc1_1 gpc1942 (
      {stage0_18[473]},
      {stage1_18[188]}
   );
   gpc1_1 gpc1943 (
      {stage0_18[474]},
      {stage1_18[189]}
   );
   gpc1_1 gpc1944 (
      {stage0_18[475]},
      {stage1_18[190]}
   );
   gpc1_1 gpc1945 (
      {stage0_18[476]},
      {stage1_18[191]}
   );
   gpc1_1 gpc1946 (
      {stage0_18[477]},
      {stage1_18[192]}
   );
   gpc1_1 gpc1947 (
      {stage0_18[478]},
      {stage1_18[193]}
   );
   gpc1_1 gpc1948 (
      {stage0_18[479]},
      {stage1_18[194]}
   );
   gpc1_1 gpc1949 (
      {stage0_18[480]},
      {stage1_18[195]}
   );
   gpc1_1 gpc1950 (
      {stage0_18[481]},
      {stage1_18[196]}
   );
   gpc1_1 gpc1951 (
      {stage0_18[482]},
      {stage1_18[197]}
   );
   gpc1_1 gpc1952 (
      {stage0_18[483]},
      {stage1_18[198]}
   );
   gpc1_1 gpc1953 (
      {stage0_18[484]},
      {stage1_18[199]}
   );
   gpc1_1 gpc1954 (
      {stage0_18[485]},
      {stage1_18[200]}
   );
   gpc1_1 gpc1955 (
      {stage0_19[347]},
      {stage1_19[161]}
   );
   gpc1_1 gpc1956 (
      {stage0_19[348]},
      {stage1_19[162]}
   );
   gpc1_1 gpc1957 (
      {stage0_19[349]},
      {stage1_19[163]}
   );
   gpc1_1 gpc1958 (
      {stage0_19[350]},
      {stage1_19[164]}
   );
   gpc1_1 gpc1959 (
      {stage0_19[351]},
      {stage1_19[165]}
   );
   gpc1_1 gpc1960 (
      {stage0_19[352]},
      {stage1_19[166]}
   );
   gpc1_1 gpc1961 (
      {stage0_19[353]},
      {stage1_19[167]}
   );
   gpc1_1 gpc1962 (
      {stage0_19[354]},
      {stage1_19[168]}
   );
   gpc1_1 gpc1963 (
      {stage0_19[355]},
      {stage1_19[169]}
   );
   gpc1_1 gpc1964 (
      {stage0_19[356]},
      {stage1_19[170]}
   );
   gpc1_1 gpc1965 (
      {stage0_19[357]},
      {stage1_19[171]}
   );
   gpc1_1 gpc1966 (
      {stage0_19[358]},
      {stage1_19[172]}
   );
   gpc1_1 gpc1967 (
      {stage0_19[359]},
      {stage1_19[173]}
   );
   gpc1_1 gpc1968 (
      {stage0_19[360]},
      {stage1_19[174]}
   );
   gpc1_1 gpc1969 (
      {stage0_19[361]},
      {stage1_19[175]}
   );
   gpc1_1 gpc1970 (
      {stage0_19[362]},
      {stage1_19[176]}
   );
   gpc1_1 gpc1971 (
      {stage0_19[363]},
      {stage1_19[177]}
   );
   gpc1_1 gpc1972 (
      {stage0_19[364]},
      {stage1_19[178]}
   );
   gpc1_1 gpc1973 (
      {stage0_19[365]},
      {stage1_19[179]}
   );
   gpc1_1 gpc1974 (
      {stage0_19[366]},
      {stage1_19[180]}
   );
   gpc1_1 gpc1975 (
      {stage0_19[367]},
      {stage1_19[181]}
   );
   gpc1_1 gpc1976 (
      {stage0_19[368]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1977 (
      {stage0_19[369]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1978 (
      {stage0_19[370]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1979 (
      {stage0_19[371]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1980 (
      {stage0_19[372]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1981 (
      {stage0_19[373]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1982 (
      {stage0_19[374]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1983 (
      {stage0_19[375]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1984 (
      {stage0_19[376]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1985 (
      {stage0_19[377]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1986 (
      {stage0_19[378]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1987 (
      {stage0_19[379]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1988 (
      {stage0_19[380]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1989 (
      {stage0_19[381]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1990 (
      {stage0_19[382]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1991 (
      {stage0_19[383]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1992 (
      {stage0_19[384]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1993 (
      {stage0_19[385]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1994 (
      {stage0_19[386]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1995 (
      {stage0_19[387]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1996 (
      {stage0_19[388]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1997 (
      {stage0_19[389]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1998 (
      {stage0_19[390]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1999 (
      {stage0_19[391]},
      {stage1_19[205]}
   );
   gpc1_1 gpc2000 (
      {stage0_19[392]},
      {stage1_19[206]}
   );
   gpc1_1 gpc2001 (
      {stage0_19[393]},
      {stage1_19[207]}
   );
   gpc1_1 gpc2002 (
      {stage0_19[394]},
      {stage1_19[208]}
   );
   gpc1_1 gpc2003 (
      {stage0_19[395]},
      {stage1_19[209]}
   );
   gpc1_1 gpc2004 (
      {stage0_19[396]},
      {stage1_19[210]}
   );
   gpc1_1 gpc2005 (
      {stage0_19[397]},
      {stage1_19[211]}
   );
   gpc1_1 gpc2006 (
      {stage0_19[398]},
      {stage1_19[212]}
   );
   gpc1_1 gpc2007 (
      {stage0_19[399]},
      {stage1_19[213]}
   );
   gpc1_1 gpc2008 (
      {stage0_19[400]},
      {stage1_19[214]}
   );
   gpc1_1 gpc2009 (
      {stage0_19[401]},
      {stage1_19[215]}
   );
   gpc1_1 gpc2010 (
      {stage0_19[402]},
      {stage1_19[216]}
   );
   gpc1_1 gpc2011 (
      {stage0_19[403]},
      {stage1_19[217]}
   );
   gpc1_1 gpc2012 (
      {stage0_19[404]},
      {stage1_19[218]}
   );
   gpc1_1 gpc2013 (
      {stage0_19[405]},
      {stage1_19[219]}
   );
   gpc1_1 gpc2014 (
      {stage0_19[406]},
      {stage1_19[220]}
   );
   gpc1_1 gpc2015 (
      {stage0_19[407]},
      {stage1_19[221]}
   );
   gpc1_1 gpc2016 (
      {stage0_19[408]},
      {stage1_19[222]}
   );
   gpc1_1 gpc2017 (
      {stage0_19[409]},
      {stage1_19[223]}
   );
   gpc1_1 gpc2018 (
      {stage0_19[410]},
      {stage1_19[224]}
   );
   gpc1_1 gpc2019 (
      {stage0_19[411]},
      {stage1_19[225]}
   );
   gpc1_1 gpc2020 (
      {stage0_19[412]},
      {stage1_19[226]}
   );
   gpc1_1 gpc2021 (
      {stage0_19[413]},
      {stage1_19[227]}
   );
   gpc1_1 gpc2022 (
      {stage0_19[414]},
      {stage1_19[228]}
   );
   gpc1_1 gpc2023 (
      {stage0_19[415]},
      {stage1_19[229]}
   );
   gpc1_1 gpc2024 (
      {stage0_19[416]},
      {stage1_19[230]}
   );
   gpc1_1 gpc2025 (
      {stage0_19[417]},
      {stage1_19[231]}
   );
   gpc1_1 gpc2026 (
      {stage0_19[418]},
      {stage1_19[232]}
   );
   gpc1_1 gpc2027 (
      {stage0_19[419]},
      {stage1_19[233]}
   );
   gpc1_1 gpc2028 (
      {stage0_19[420]},
      {stage1_19[234]}
   );
   gpc1_1 gpc2029 (
      {stage0_19[421]},
      {stage1_19[235]}
   );
   gpc1_1 gpc2030 (
      {stage0_19[422]},
      {stage1_19[236]}
   );
   gpc1_1 gpc2031 (
      {stage0_19[423]},
      {stage1_19[237]}
   );
   gpc1_1 gpc2032 (
      {stage0_19[424]},
      {stage1_19[238]}
   );
   gpc1_1 gpc2033 (
      {stage0_19[425]},
      {stage1_19[239]}
   );
   gpc1_1 gpc2034 (
      {stage0_19[426]},
      {stage1_19[240]}
   );
   gpc1_1 gpc2035 (
      {stage0_19[427]},
      {stage1_19[241]}
   );
   gpc1_1 gpc2036 (
      {stage0_19[428]},
      {stage1_19[242]}
   );
   gpc1_1 gpc2037 (
      {stage0_19[429]},
      {stage1_19[243]}
   );
   gpc1_1 gpc2038 (
      {stage0_19[430]},
      {stage1_19[244]}
   );
   gpc1_1 gpc2039 (
      {stage0_19[431]},
      {stage1_19[245]}
   );
   gpc1_1 gpc2040 (
      {stage0_19[432]},
      {stage1_19[246]}
   );
   gpc1_1 gpc2041 (
      {stage0_19[433]},
      {stage1_19[247]}
   );
   gpc1_1 gpc2042 (
      {stage0_19[434]},
      {stage1_19[248]}
   );
   gpc1_1 gpc2043 (
      {stage0_19[435]},
      {stage1_19[249]}
   );
   gpc1_1 gpc2044 (
      {stage0_19[436]},
      {stage1_19[250]}
   );
   gpc1_1 gpc2045 (
      {stage0_19[437]},
      {stage1_19[251]}
   );
   gpc1_1 gpc2046 (
      {stage0_19[438]},
      {stage1_19[252]}
   );
   gpc1_1 gpc2047 (
      {stage0_19[439]},
      {stage1_19[253]}
   );
   gpc1_1 gpc2048 (
      {stage0_19[440]},
      {stage1_19[254]}
   );
   gpc1_1 gpc2049 (
      {stage0_19[441]},
      {stage1_19[255]}
   );
   gpc1_1 gpc2050 (
      {stage0_19[442]},
      {stage1_19[256]}
   );
   gpc1_1 gpc2051 (
      {stage0_19[443]},
      {stage1_19[257]}
   );
   gpc1_1 gpc2052 (
      {stage0_19[444]},
      {stage1_19[258]}
   );
   gpc1_1 gpc2053 (
      {stage0_19[445]},
      {stage1_19[259]}
   );
   gpc1_1 gpc2054 (
      {stage0_19[446]},
      {stage1_19[260]}
   );
   gpc1_1 gpc2055 (
      {stage0_19[447]},
      {stage1_19[261]}
   );
   gpc1_1 gpc2056 (
      {stage0_19[448]},
      {stage1_19[262]}
   );
   gpc1_1 gpc2057 (
      {stage0_19[449]},
      {stage1_19[263]}
   );
   gpc1_1 gpc2058 (
      {stage0_19[450]},
      {stage1_19[264]}
   );
   gpc1_1 gpc2059 (
      {stage0_19[451]},
      {stage1_19[265]}
   );
   gpc1_1 gpc2060 (
      {stage0_19[452]},
      {stage1_19[266]}
   );
   gpc1_1 gpc2061 (
      {stage0_19[453]},
      {stage1_19[267]}
   );
   gpc1_1 gpc2062 (
      {stage0_19[454]},
      {stage1_19[268]}
   );
   gpc1_1 gpc2063 (
      {stage0_19[455]},
      {stage1_19[269]}
   );
   gpc1_1 gpc2064 (
      {stage0_19[456]},
      {stage1_19[270]}
   );
   gpc1_1 gpc2065 (
      {stage0_19[457]},
      {stage1_19[271]}
   );
   gpc1_1 gpc2066 (
      {stage0_19[458]},
      {stage1_19[272]}
   );
   gpc1_1 gpc2067 (
      {stage0_19[459]},
      {stage1_19[273]}
   );
   gpc1_1 gpc2068 (
      {stage0_19[460]},
      {stage1_19[274]}
   );
   gpc1_1 gpc2069 (
      {stage0_19[461]},
      {stage1_19[275]}
   );
   gpc1_1 gpc2070 (
      {stage0_19[462]},
      {stage1_19[276]}
   );
   gpc1_1 gpc2071 (
      {stage0_19[463]},
      {stage1_19[277]}
   );
   gpc1_1 gpc2072 (
      {stage0_19[464]},
      {stage1_19[278]}
   );
   gpc1_1 gpc2073 (
      {stage0_19[465]},
      {stage1_19[279]}
   );
   gpc1_1 gpc2074 (
      {stage0_19[466]},
      {stage1_19[280]}
   );
   gpc1_1 gpc2075 (
      {stage0_19[467]},
      {stage1_19[281]}
   );
   gpc1_1 gpc2076 (
      {stage0_19[468]},
      {stage1_19[282]}
   );
   gpc1_1 gpc2077 (
      {stage0_19[469]},
      {stage1_19[283]}
   );
   gpc1_1 gpc2078 (
      {stage0_19[470]},
      {stage1_19[284]}
   );
   gpc1_1 gpc2079 (
      {stage0_19[471]},
      {stage1_19[285]}
   );
   gpc1_1 gpc2080 (
      {stage0_19[472]},
      {stage1_19[286]}
   );
   gpc1_1 gpc2081 (
      {stage0_19[473]},
      {stage1_19[287]}
   );
   gpc1_1 gpc2082 (
      {stage0_19[474]},
      {stage1_19[288]}
   );
   gpc1_1 gpc2083 (
      {stage0_19[475]},
      {stage1_19[289]}
   );
   gpc1_1 gpc2084 (
      {stage0_19[476]},
      {stage1_19[290]}
   );
   gpc1_1 gpc2085 (
      {stage0_19[477]},
      {stage1_19[291]}
   );
   gpc1_1 gpc2086 (
      {stage0_19[478]},
      {stage1_19[292]}
   );
   gpc1_1 gpc2087 (
      {stage0_19[479]},
      {stage1_19[293]}
   );
   gpc1_1 gpc2088 (
      {stage0_19[480]},
      {stage1_19[294]}
   );
   gpc1_1 gpc2089 (
      {stage0_19[481]},
      {stage1_19[295]}
   );
   gpc1_1 gpc2090 (
      {stage0_19[482]},
      {stage1_19[296]}
   );
   gpc1_1 gpc2091 (
      {stage0_19[483]},
      {stage1_19[297]}
   );
   gpc1_1 gpc2092 (
      {stage0_19[484]},
      {stage1_19[298]}
   );
   gpc1_1 gpc2093 (
      {stage0_19[485]},
      {stage1_19[299]}
   );
   gpc1_1 gpc2094 (
      {stage0_20[478]},
      {stage1_20[181]}
   );
   gpc1_1 gpc2095 (
      {stage0_20[479]},
      {stage1_20[182]}
   );
   gpc1_1 gpc2096 (
      {stage0_20[480]},
      {stage1_20[183]}
   );
   gpc1_1 gpc2097 (
      {stage0_20[481]},
      {stage1_20[184]}
   );
   gpc1_1 gpc2098 (
      {stage0_20[482]},
      {stage1_20[185]}
   );
   gpc1_1 gpc2099 (
      {stage0_20[483]},
      {stage1_20[186]}
   );
   gpc1_1 gpc2100 (
      {stage0_20[484]},
      {stage1_20[187]}
   );
   gpc1_1 gpc2101 (
      {stage0_20[485]},
      {stage1_20[188]}
   );
   gpc1_1 gpc2102 (
      {stage0_22[422]},
      {stage1_22[187]}
   );
   gpc1_1 gpc2103 (
      {stage0_22[423]},
      {stage1_22[188]}
   );
   gpc1_1 gpc2104 (
      {stage0_22[424]},
      {stage1_22[189]}
   );
   gpc1_1 gpc2105 (
      {stage0_22[425]},
      {stage1_22[190]}
   );
   gpc1_1 gpc2106 (
      {stage0_22[426]},
      {stage1_22[191]}
   );
   gpc1_1 gpc2107 (
      {stage0_22[427]},
      {stage1_22[192]}
   );
   gpc1_1 gpc2108 (
      {stage0_22[428]},
      {stage1_22[193]}
   );
   gpc1_1 gpc2109 (
      {stage0_22[429]},
      {stage1_22[194]}
   );
   gpc1_1 gpc2110 (
      {stage0_22[430]},
      {stage1_22[195]}
   );
   gpc1_1 gpc2111 (
      {stage0_22[431]},
      {stage1_22[196]}
   );
   gpc1_1 gpc2112 (
      {stage0_22[432]},
      {stage1_22[197]}
   );
   gpc1_1 gpc2113 (
      {stage0_22[433]},
      {stage1_22[198]}
   );
   gpc1_1 gpc2114 (
      {stage0_22[434]},
      {stage1_22[199]}
   );
   gpc1_1 gpc2115 (
      {stage0_22[435]},
      {stage1_22[200]}
   );
   gpc1_1 gpc2116 (
      {stage0_22[436]},
      {stage1_22[201]}
   );
   gpc1_1 gpc2117 (
      {stage0_22[437]},
      {stage1_22[202]}
   );
   gpc1_1 gpc2118 (
      {stage0_22[438]},
      {stage1_22[203]}
   );
   gpc1_1 gpc2119 (
      {stage0_22[439]},
      {stage1_22[204]}
   );
   gpc1_1 gpc2120 (
      {stage0_22[440]},
      {stage1_22[205]}
   );
   gpc1_1 gpc2121 (
      {stage0_22[441]},
      {stage1_22[206]}
   );
   gpc1_1 gpc2122 (
      {stage0_22[442]},
      {stage1_22[207]}
   );
   gpc1_1 gpc2123 (
      {stage0_22[443]},
      {stage1_22[208]}
   );
   gpc1_1 gpc2124 (
      {stage0_22[444]},
      {stage1_22[209]}
   );
   gpc1_1 gpc2125 (
      {stage0_22[445]},
      {stage1_22[210]}
   );
   gpc1_1 gpc2126 (
      {stage0_22[446]},
      {stage1_22[211]}
   );
   gpc1_1 gpc2127 (
      {stage0_22[447]},
      {stage1_22[212]}
   );
   gpc1_1 gpc2128 (
      {stage0_22[448]},
      {stage1_22[213]}
   );
   gpc1_1 gpc2129 (
      {stage0_22[449]},
      {stage1_22[214]}
   );
   gpc1_1 gpc2130 (
      {stage0_22[450]},
      {stage1_22[215]}
   );
   gpc1_1 gpc2131 (
      {stage0_22[451]},
      {stage1_22[216]}
   );
   gpc1_1 gpc2132 (
      {stage0_22[452]},
      {stage1_22[217]}
   );
   gpc1_1 gpc2133 (
      {stage0_22[453]},
      {stage1_22[218]}
   );
   gpc1_1 gpc2134 (
      {stage0_22[454]},
      {stage1_22[219]}
   );
   gpc1_1 gpc2135 (
      {stage0_22[455]},
      {stage1_22[220]}
   );
   gpc1_1 gpc2136 (
      {stage0_22[456]},
      {stage1_22[221]}
   );
   gpc1_1 gpc2137 (
      {stage0_22[457]},
      {stage1_22[222]}
   );
   gpc1_1 gpc2138 (
      {stage0_22[458]},
      {stage1_22[223]}
   );
   gpc1_1 gpc2139 (
      {stage0_22[459]},
      {stage1_22[224]}
   );
   gpc1_1 gpc2140 (
      {stage0_22[460]},
      {stage1_22[225]}
   );
   gpc1_1 gpc2141 (
      {stage0_22[461]},
      {stage1_22[226]}
   );
   gpc1_1 gpc2142 (
      {stage0_22[462]},
      {stage1_22[227]}
   );
   gpc1_1 gpc2143 (
      {stage0_22[463]},
      {stage1_22[228]}
   );
   gpc1_1 gpc2144 (
      {stage0_22[464]},
      {stage1_22[229]}
   );
   gpc1_1 gpc2145 (
      {stage0_22[465]},
      {stage1_22[230]}
   );
   gpc1_1 gpc2146 (
      {stage0_22[466]},
      {stage1_22[231]}
   );
   gpc1_1 gpc2147 (
      {stage0_22[467]},
      {stage1_22[232]}
   );
   gpc1_1 gpc2148 (
      {stage0_22[468]},
      {stage1_22[233]}
   );
   gpc1_1 gpc2149 (
      {stage0_22[469]},
      {stage1_22[234]}
   );
   gpc1_1 gpc2150 (
      {stage0_22[470]},
      {stage1_22[235]}
   );
   gpc1_1 gpc2151 (
      {stage0_22[471]},
      {stage1_22[236]}
   );
   gpc1_1 gpc2152 (
      {stage0_22[472]},
      {stage1_22[237]}
   );
   gpc1_1 gpc2153 (
      {stage0_22[473]},
      {stage1_22[238]}
   );
   gpc1_1 gpc2154 (
      {stage0_22[474]},
      {stage1_22[239]}
   );
   gpc1_1 gpc2155 (
      {stage0_22[475]},
      {stage1_22[240]}
   );
   gpc1_1 gpc2156 (
      {stage0_22[476]},
      {stage1_22[241]}
   );
   gpc1_1 gpc2157 (
      {stage0_22[477]},
      {stage1_22[242]}
   );
   gpc1_1 gpc2158 (
      {stage0_22[478]},
      {stage1_22[243]}
   );
   gpc1_1 gpc2159 (
      {stage0_22[479]},
      {stage1_22[244]}
   );
   gpc1_1 gpc2160 (
      {stage0_22[480]},
      {stage1_22[245]}
   );
   gpc1_1 gpc2161 (
      {stage0_22[481]},
      {stage1_22[246]}
   );
   gpc1_1 gpc2162 (
      {stage0_22[482]},
      {stage1_22[247]}
   );
   gpc1_1 gpc2163 (
      {stage0_22[483]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2164 (
      {stage0_22[484]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2165 (
      {stage0_22[485]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2166 (
      {stage0_23[474]},
      {stage1_23[166]}
   );
   gpc1_1 gpc2167 (
      {stage0_23[475]},
      {stage1_23[167]}
   );
   gpc1_1 gpc2168 (
      {stage0_23[476]},
      {stage1_23[168]}
   );
   gpc1_1 gpc2169 (
      {stage0_23[477]},
      {stage1_23[169]}
   );
   gpc1_1 gpc2170 (
      {stage0_23[478]},
      {stage1_23[170]}
   );
   gpc1_1 gpc2171 (
      {stage0_23[479]},
      {stage1_23[171]}
   );
   gpc1_1 gpc2172 (
      {stage0_23[480]},
      {stage1_23[172]}
   );
   gpc1_1 gpc2173 (
      {stage0_23[481]},
      {stage1_23[173]}
   );
   gpc1_1 gpc2174 (
      {stage0_23[482]},
      {stage1_23[174]}
   );
   gpc1_1 gpc2175 (
      {stage0_23[483]},
      {stage1_23[175]}
   );
   gpc1_1 gpc2176 (
      {stage0_23[484]},
      {stage1_23[176]}
   );
   gpc1_1 gpc2177 (
      {stage0_23[485]},
      {stage1_23[177]}
   );
   gpc1_1 gpc2178 (
      {stage0_26[445]},
      {stage1_26[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_26[446]},
      {stage1_26[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_26[447]},
      {stage1_26[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_26[448]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_26[449]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_26[450]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_26[451]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_26[452]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_26[453]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_26[454]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_26[455]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_26[456]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_26[457]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_26[458]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_26[459]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_26[460]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_26[461]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_26[462]},
      {stage1_26[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_26[463]},
      {stage1_26[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_26[464]},
      {stage1_26[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_26[465]},
      {stage1_26[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_26[466]},
      {stage1_26[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_26[467]},
      {stage1_26[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_26[468]},
      {stage1_26[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_26[469]},
      {stage1_26[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_26[470]},
      {stage1_26[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_26[471]},
      {stage1_26[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_26[472]},
      {stage1_26[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_26[473]},
      {stage1_26[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_26[474]},
      {stage1_26[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_26[475]},
      {stage1_26[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_26[476]},
      {stage1_26[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_26[477]},
      {stage1_26[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_26[478]},
      {stage1_26[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_26[479]},
      {stage1_26[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_26[480]},
      {stage1_26[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_26[481]},
      {stage1_26[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_26[482]},
      {stage1_26[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_26[483]},
      {stage1_26[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_26[484]},
      {stage1_26[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_26[485]},
      {stage1_26[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_27[483]},
      {stage1_27[156]}
   );
   gpc1_1 gpc2220 (
      {stage0_27[484]},
      {stage1_27[157]}
   );
   gpc1_1 gpc2221 (
      {stage0_27[485]},
      {stage1_27[158]}
   );
   gpc1_1 gpc2222 (
      {stage0_28[450]},
      {stage1_28[216]}
   );
   gpc1_1 gpc2223 (
      {stage0_28[451]},
      {stage1_28[217]}
   );
   gpc1_1 gpc2224 (
      {stage0_28[452]},
      {stage1_28[218]}
   );
   gpc1_1 gpc2225 (
      {stage0_28[453]},
      {stage1_28[219]}
   );
   gpc1_1 gpc2226 (
      {stage0_28[454]},
      {stage1_28[220]}
   );
   gpc1_1 gpc2227 (
      {stage0_28[455]},
      {stage1_28[221]}
   );
   gpc1_1 gpc2228 (
      {stage0_28[456]},
      {stage1_28[222]}
   );
   gpc1_1 gpc2229 (
      {stage0_28[457]},
      {stage1_28[223]}
   );
   gpc1_1 gpc2230 (
      {stage0_28[458]},
      {stage1_28[224]}
   );
   gpc1_1 gpc2231 (
      {stage0_28[459]},
      {stage1_28[225]}
   );
   gpc1_1 gpc2232 (
      {stage0_28[460]},
      {stage1_28[226]}
   );
   gpc1_1 gpc2233 (
      {stage0_28[461]},
      {stage1_28[227]}
   );
   gpc1_1 gpc2234 (
      {stage0_28[462]},
      {stage1_28[228]}
   );
   gpc1_1 gpc2235 (
      {stage0_28[463]},
      {stage1_28[229]}
   );
   gpc1_1 gpc2236 (
      {stage0_28[464]},
      {stage1_28[230]}
   );
   gpc1_1 gpc2237 (
      {stage0_28[465]},
      {stage1_28[231]}
   );
   gpc1_1 gpc2238 (
      {stage0_28[466]},
      {stage1_28[232]}
   );
   gpc1_1 gpc2239 (
      {stage0_28[467]},
      {stage1_28[233]}
   );
   gpc1_1 gpc2240 (
      {stage0_28[468]},
      {stage1_28[234]}
   );
   gpc1_1 gpc2241 (
      {stage0_28[469]},
      {stage1_28[235]}
   );
   gpc1_1 gpc2242 (
      {stage0_28[470]},
      {stage1_28[236]}
   );
   gpc1_1 gpc2243 (
      {stage0_28[471]},
      {stage1_28[237]}
   );
   gpc1_1 gpc2244 (
      {stage0_28[472]},
      {stage1_28[238]}
   );
   gpc1_1 gpc2245 (
      {stage0_28[473]},
      {stage1_28[239]}
   );
   gpc1_1 gpc2246 (
      {stage0_28[474]},
      {stage1_28[240]}
   );
   gpc1_1 gpc2247 (
      {stage0_28[475]},
      {stage1_28[241]}
   );
   gpc1_1 gpc2248 (
      {stage0_28[476]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2249 (
      {stage0_28[477]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2250 (
      {stage0_28[478]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2251 (
      {stage0_28[479]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2252 (
      {stage0_28[480]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2253 (
      {stage0_28[481]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2254 (
      {stage0_28[482]},
      {stage1_28[248]}
   );
   gpc1_1 gpc2255 (
      {stage0_28[483]},
      {stage1_28[249]}
   );
   gpc1_1 gpc2256 (
      {stage0_28[484]},
      {stage1_28[250]}
   );
   gpc1_1 gpc2257 (
      {stage0_28[485]},
      {stage1_28[251]}
   );
   gpc1_1 gpc2258 (
      {stage0_30[480]},
      {stage1_30[166]}
   );
   gpc1_1 gpc2259 (
      {stage0_30[481]},
      {stage1_30[167]}
   );
   gpc1_1 gpc2260 (
      {stage0_30[482]},
      {stage1_30[168]}
   );
   gpc1_1 gpc2261 (
      {stage0_30[483]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2262 (
      {stage0_30[484]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2263 (
      {stage0_30[485]},
      {stage1_30[171]}
   );
   gpc1163_5 gpc2264 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc2265 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc2266 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2267 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2268 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc2269 (
      {stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc2270 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2271 (
      {stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc2272 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc2273 (
      {stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc2274 (
      {stage1_0[57], stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc2275 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67], stage1_0[68]},
      {stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2276 (
      {stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72], stage1_0[73], stage1_0[74]},
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc2277 (
      {stage1_0[75], stage1_0[76], stage1_0[77], stage1_0[78], stage1_0[79], stage1_0[80]},
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc2278 (
      {stage1_0[81], stage1_0[82], stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86]},
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83], stage1_2[84]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc2279 (
      {stage1_0[87], stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc2280 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97], stage1_0[98]},
      {stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc2281 (
      {stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102], stage1_0[103], stage1_0[104]},
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc2282 (
      {stage1_0[105], stage1_0[106], stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110]},
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107], stage1_2[108]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc2283 (
      {stage1_0[111], stage1_0[112], stage1_0[113], stage1_0[114], stage1_0[115], stage1_0[116]},
      {stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113], stage1_2[114]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc2284 (
      {stage1_0[117], stage1_0[118], stage1_0[119], stage1_0[120], stage1_0[121]},
      {stage1_1[6]},
      {stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc615_5 gpc2285 (
      {stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125], stage1_0[126]},
      {stage1_1[7]},
      {stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc2286 (
      {stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2287 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage2_5[1],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2288 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18]},
      {stage2_5[2],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2289 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage2_5[3],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2290 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30]},
      {stage2_5[4],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2291 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage2_5[5],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2292 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage2_5[6],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2293 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage2_5[7],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2294 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54]},
      {stage2_5[8],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2295 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[9],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc606_5 gpc2296 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137], stage1_2[138]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[10],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc606_5 gpc2297 (
      {stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143], stage1_2[144]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[11],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc606_5 gpc2298 (
      {stage1_2[145], stage1_2[146], stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[12],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc606_5 gpc2299 (
      {stage1_2[151], stage1_2[152], stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[13],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc606_5 gpc2300 (
      {stage1_2[157], stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[14],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc606_5 gpc2301 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167], stage1_2[168]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[15],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc606_5 gpc2302 (
      {stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172], stage1_2[173], stage1_2[174]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[16],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc606_5 gpc2303 (
      {stage1_2[175], stage1_2[176], stage1_2[177], stage1_2[178], stage1_2[179], stage1_2[180]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[17],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc2304 (
      {stage1_2[181], stage1_2[182], stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[18],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc2305 (
      {stage1_2[187], stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[19],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc2306 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197], stage1_2[198]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[20],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc2307 (
      {stage1_2[199], stage1_2[200], stage1_2[201], stage1_2[202], stage1_2[203], stage1_2[204]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[21],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2308 (
      {stage1_2[205], stage1_2[206], stage1_2[207], stage1_2[208], stage1_2[209]},
      {stage1_3[55]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[22],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2309 (
      {stage1_2[210], stage1_2[211], stage1_2[212], stage1_2[213], stage1_2[214]},
      {stage1_3[56]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[23],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2310 (
      {stage1_2[215], stage1_2[216], stage1_2[217], stage1_2[218], stage1_2[219]},
      {stage1_3[57]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[24],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2311 (
      {stage1_2[220], stage1_2[221], stage1_2[222], stage1_2[223], stage1_2[224]},
      {stage1_3[58]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[25],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc2312 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[17],stage2_5[26],stage2_4[48],stage2_3[48]}
   );
   gpc606_5 gpc2313 (
      {stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[18],stage2_5[27],stage2_4[49],stage2_3[49]}
   );
   gpc606_5 gpc2314 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[19],stage2_5[28],stage2_4[50],stage2_3[50]}
   );
   gpc606_5 gpc2315 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[20],stage2_5[29],stage2_4[51],stage2_3[51]}
   );
   gpc606_5 gpc2316 (
      {stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[21],stage2_5[30],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93]},
      {stage1_4[102]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[22],stage2_5[31],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97], stage1_3[98]},
      {stage1_4[103]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[23],stage2_5[32],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage1_4[104]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[24],stage2_5[33],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108]},
      {stage1_4[105]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[25],stage2_5[34],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage1_4[106]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[26],stage2_5[35],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118]},
      {stage1_4[107]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[27],stage2_5[36],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123]},
      {stage1_4[108]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[28],stage2_5[37],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2324 (
      {stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127], stage1_3[128]},
      {stage1_4[109]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[29],stage2_5[38],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2325 (
      {stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage1_4[110]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[30],stage2_5[39],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2326 (
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[111]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[31],stage2_5[40],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2327 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[112]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[32],stage2_5[41],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2328 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[113]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[33],stage2_5[42],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2329 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[114]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[34],stage2_5[43],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2330 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[115]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[35],stage2_5[44],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2331 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[116]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[36],stage2_5[45],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2332 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[117]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[37],stage2_5[46],stage2_4[68],stage2_3[68]}
   );
   gpc1163_5 gpc2333 (
      {stage1_4[118], stage1_4[119], stage1_4[120]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[21],stage2_6[38],stage2_5[47],stage2_4[69]}
   );
   gpc615_5 gpc2334 (
      {stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage1_5[132]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[22],stage2_6[39],stage2_5[48],stage2_4[70]}
   );
   gpc615_5 gpc2335 (
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130]},
      {stage1_5[133]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[23],stage2_6[40],stage2_5[49],stage2_4[71]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_5[134]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[24],stage2_6[41],stage2_5[50],stage2_4[72]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[135]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[25],stage2_6[42],stage2_5[51],stage2_4[73]}
   );
   gpc615_5 gpc2338 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145]},
      {stage1_5[136]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[26],stage2_6[43],stage2_5[52],stage2_4[74]}
   );
   gpc615_5 gpc2339 (
      {stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_5[137]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[27],stage2_6[44],stage2_5[53],stage2_4[75]}
   );
   gpc615_5 gpc2340 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage1_5[138]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[28],stage2_6[45],stage2_5[54],stage2_4[76]}
   );
   gpc615_5 gpc2341 (
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160]},
      {stage1_5[139]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[29],stage2_6[46],stage2_5[55],stage2_4[77]}
   );
   gpc615_5 gpc2342 (
      {stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_5[140]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[30],stage2_6[47],stage2_5[56],stage2_4[78]}
   );
   gpc615_5 gpc2343 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_5[141]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[31],stage2_6[48],stage2_5[57],stage2_4[79]}
   );
   gpc615_5 gpc2344 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175]},
      {stage1_5[142]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[32],stage2_6[49],stage2_5[58],stage2_4[80]}
   );
   gpc615_5 gpc2345 (
      {stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_5[143]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[33],stage2_6[50],stage2_5[59],stage2_4[81]}
   );
   gpc615_5 gpc2346 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage1_5[144]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[34],stage2_6[51],stage2_5[60],stage2_4[82]}
   );
   gpc615_5 gpc2347 (
      {stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190]},
      {stage1_5[145]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[35],stage2_6[52],stage2_5[61],stage2_4[83]}
   );
   gpc615_5 gpc2348 (
      {stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_5[146]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[36],stage2_6[53],stage2_5[62],stage2_4[84]}
   );
   gpc615_5 gpc2349 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_5[147]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[37],stage2_6[54],stage2_5[63],stage2_4[85]}
   );
   gpc615_5 gpc2350 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205]},
      {stage1_5[148]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[38],stage2_6[55],stage2_5[64],stage2_4[86]}
   );
   gpc615_5 gpc2351 (
      {stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_5[149]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[39],stage2_6[56],stage2_5[65],stage2_4[87]}
   );
   gpc615_5 gpc2352 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215]},
      {stage1_5[150]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[40],stage2_6[57],stage2_5[66],stage2_4[88]}
   );
   gpc615_5 gpc2353 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220]},
      {stage1_5[151]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[41],stage2_6[58],stage2_5[67],stage2_4[89]}
   );
   gpc615_5 gpc2354 (
      {stage1_4[221], stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225]},
      {stage1_5[152]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[42],stage2_6[59],stage2_5[68],stage2_4[90]}
   );
   gpc606_5 gpc2355 (
      {stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157], stage1_5[158]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[22],stage2_7[43],stage2_6[60],stage2_5[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163], stage1_5[164]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[23],stage2_7[44],stage2_6[61],stage2_5[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169], stage1_5[170]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[24],stage2_7[45],stage2_6[62],stage2_5[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175], stage1_5[176]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[25],stage2_7[46],stage2_6[63],stage2_5[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181], stage1_5[182]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[26],stage2_7[47],stage2_6[64],stage2_5[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187], stage1_5[188]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[27],stage2_7[48],stage2_6[65],stage2_5[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193], stage1_5[194]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[28],stage2_7[49],stage2_6[66],stage2_5[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199], stage1_5[200]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[29],stage2_7[50],stage2_6[67],stage2_5[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205], stage1_5[206]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[30],stage2_7[51],stage2_6[68],stage2_5[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_5[207], stage1_5[208], stage1_5[209], stage1_5[210], stage1_5[211], stage1_5[212]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[31],stage2_7[52],stage2_6[69],stage2_5[78]}
   );
   gpc615_5 gpc2365 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_7[61]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[10],stage2_8[32],stage2_7[53],stage2_6[70]}
   );
   gpc615_5 gpc2366 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136]},
      {stage1_7[62]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[11],stage2_8[33],stage2_7[54],stage2_6[71]}
   );
   gpc615_5 gpc2367 (
      {stage1_6[137], stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141]},
      {stage1_7[63]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[12],stage2_8[34],stage2_7[55],stage2_6[72]}
   );
   gpc615_5 gpc2368 (
      {stage1_6[142], stage1_6[143], stage1_6[144], stage1_6[145], stage1_6[146]},
      {stage1_7[64]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[13],stage2_8[35],stage2_7[56],stage2_6[73]}
   );
   gpc615_5 gpc2369 (
      {stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150], stage1_6[151]},
      {stage1_7[65]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[14],stage2_8[36],stage2_7[57],stage2_6[74]}
   );
   gpc615_5 gpc2370 (
      {stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_7[66]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[15],stage2_8[37],stage2_7[58],stage2_6[75]}
   );
   gpc615_5 gpc2371 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_7[67]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[16],stage2_8[38],stage2_7[59],stage2_6[76]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166]},
      {stage1_7[68]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[17],stage2_8[39],stage2_7[60],stage2_6[77]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[167], stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171]},
      {stage1_7[69]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[18],stage2_8[40],stage2_7[61],stage2_6[78]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[172], stage1_6[173], stage1_6[174], stage1_6[175], stage1_6[176]},
      {stage1_7[70]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[19],stage2_8[41],stage2_7[62],stage2_6[79]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180], stage1_6[181]},
      {stage1_7[71]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[20],stage2_8[42],stage2_7[63],stage2_6[80]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_7[72]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[21],stage2_8[43],stage2_7[64],stage2_6[81]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_7[73]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[22],stage2_8[44],stage2_7[65],stage2_6[82]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[74]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[23],stage2_8[45],stage2_7[66],stage2_6[83]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[197], stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201]},
      {stage1_7[75]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[24],stage2_8[46],stage2_7[67],stage2_6[84]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[202], stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206]},
      {stage1_7[76]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[25],stage2_8[47],stage2_7[68],stage2_6[85]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[207], stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211]},
      {stage1_7[77]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[26],stage2_8[48],stage2_7[69],stage2_6[86]}
   );
   gpc615_5 gpc2382 (
      {stage1_6[212], stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216]},
      {stage1_7[78]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[27],stage2_8[49],stage2_7[70],stage2_6[87]}
   );
   gpc615_5 gpc2383 (
      {stage1_6[217], stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221]},
      {stage1_7[79]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[28],stage2_8[50],stage2_7[71],stage2_6[88]}
   );
   gpc615_5 gpc2384 (
      {stage1_6[222], stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226]},
      {stage1_7[80]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[29],stage2_8[51],stage2_7[72],stage2_6[89]}
   );
   gpc615_5 gpc2385 (
      {stage1_6[227], stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231]},
      {stage1_7[81]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[30],stage2_8[52],stage2_7[73],stage2_6[90]}
   );
   gpc615_5 gpc2386 (
      {stage1_6[232], stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236]},
      {stage1_7[82]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[31],stage2_8[53],stage2_7[74],stage2_6[91]}
   );
   gpc615_5 gpc2387 (
      {stage1_6[237], stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241]},
      {stage1_7[83]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[32],stage2_8[54],stage2_7[75],stage2_6[92]}
   );
   gpc615_5 gpc2388 (
      {stage1_6[242], stage1_6[243], stage1_6[244], stage1_6[245], stage1_6[246]},
      {stage1_7[84]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[33],stage2_8[55],stage2_7[76],stage2_6[93]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage1_8[144]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[24],stage2_9[34],stage2_8[56],stage2_7[77]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94]},
      {stage1_8[145]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[25],stage2_9[35],stage2_8[57],stage2_7[78]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[95], stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99]},
      {stage1_8[146]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[26],stage2_9[36],stage2_8[58],stage2_7[79]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104]},
      {stage1_8[147]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[27],stage2_9[37],stage2_8[59],stage2_7[80]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage1_8[148]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[28],stage2_9[38],stage2_8[60],stage2_7[81]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_8[149]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[29],stage2_9[39],stage2_8[61],stage2_7[82]}
   );
   gpc615_5 gpc2395 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage1_8[150]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[30],stage2_9[40],stage2_8[62],stage2_7[83]}
   );
   gpc615_5 gpc2396 (
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124]},
      {stage1_8[151]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[31],stage2_9[41],stage2_8[63],stage2_7[84]}
   );
   gpc615_5 gpc2397 (
      {stage1_7[125], stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129]},
      {stage1_8[152]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[32],stage2_9[42],stage2_8[64],stage2_7[85]}
   );
   gpc615_5 gpc2398 (
      {stage1_7[130], stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134]},
      {stage1_8[153]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[33],stage2_9[43],stage2_8[65],stage2_7[86]}
   );
   gpc615_5 gpc2399 (
      {stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139]},
      {stage1_8[154]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[34],stage2_9[44],stage2_8[66],stage2_7[87]}
   );
   gpc615_5 gpc2400 (
      {stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_8[155]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[35],stage2_9[45],stage2_8[67],stage2_7[88]}
   );
   gpc615_5 gpc2401 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149]},
      {stage1_8[156]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[36],stage2_9[46],stage2_8[68],stage2_7[89]}
   );
   gpc615_5 gpc2402 (
      {stage1_7[150], stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154]},
      {stage1_8[157]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[37],stage2_9[47],stage2_8[69],stage2_7[90]}
   );
   gpc615_5 gpc2403 (
      {stage1_7[155], stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159]},
      {stage1_8[158]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[38],stage2_9[48],stage2_8[70],stage2_7[91]}
   );
   gpc615_5 gpc2404 (
      {stage1_7[160], stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164]},
      {stage1_8[159]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[39],stage2_9[49],stage2_8[71],stage2_7[92]}
   );
   gpc615_5 gpc2405 (
      {stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169]},
      {stage1_8[160]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[40],stage2_9[50],stage2_8[72],stage2_7[93]}
   );
   gpc615_5 gpc2406 (
      {stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_8[161]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[41],stage2_9[51],stage2_8[73],stage2_7[94]}
   );
   gpc615_5 gpc2407 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179]},
      {stage1_8[162]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[42],stage2_9[52],stage2_8[74],stage2_7[95]}
   );
   gpc615_5 gpc2408 (
      {stage1_7[180], stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184]},
      {stage1_8[163]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[43],stage2_9[53],stage2_8[75],stage2_7[96]}
   );
   gpc615_5 gpc2409 (
      {stage1_7[185], stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189]},
      {stage1_8[164]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[44],stage2_9[54],stage2_8[76],stage2_7[97]}
   );
   gpc615_5 gpc2410 (
      {stage1_7[190], stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194]},
      {stage1_8[165]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[45],stage2_9[55],stage2_8[77],stage2_7[98]}
   );
   gpc615_5 gpc2411 (
      {stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199]},
      {stage1_8[166]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[46],stage2_9[56],stage2_8[78],stage2_7[99]}
   );
   gpc615_5 gpc2412 (
      {stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_8[167]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[47],stage2_9[57],stage2_8[79],stage2_7[100]}
   );
   gpc615_5 gpc2413 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209]},
      {stage1_8[168]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[48],stage2_9[58],stage2_8[80],stage2_7[101]}
   );
   gpc615_5 gpc2414 (
      {stage1_7[210], stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214]},
      {stage1_8[169]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[49],stage2_9[59],stage2_8[81],stage2_7[102]}
   );
   gpc623_5 gpc2415 (
      {stage1_7[215], stage1_7[216], stage1_7[217]},
      {stage1_8[170], stage1_8[171]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[50],stage2_9[60],stage2_8[82],stage2_7[103]}
   );
   gpc1415_5 gpc2416 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176]},
      {stage1_9[162]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[27],stage2_10[51],stage2_9[61],stage2_8[83]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[177], stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9]},
      {stage2_12[1],stage2_11[28],stage2_10[52],stage2_9[62],stage2_8[84]}
   );
   gpc606_5 gpc2418 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[29],stage2_10[53],stage2_9[63]}
   );
   gpc606_5 gpc2419 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[30],stage2_10[54],stage2_9[64]}
   );
   gpc606_5 gpc2420 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[31],stage2_10[55],stage2_9[65]}
   );
   gpc615_5 gpc2421 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_10[10]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[3],stage2_12[5],stage2_11[32],stage2_10[56],stage2_9[66]}
   );
   gpc615_5 gpc2422 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190]},
      {stage1_10[11]},
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage2_13[4],stage2_12[6],stage2_11[33],stage2_10[57],stage2_9[67]}
   );
   gpc615_5 gpc2423 (
      {stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_10[12]},
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage2_13[5],stage2_12[7],stage2_11[34],stage2_10[58],stage2_9[68]}
   );
   gpc615_5 gpc2424 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200]},
      {stage1_10[13]},
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage2_13[6],stage2_12[8],stage2_11[35],stage2_10[59],stage2_9[69]}
   );
   gpc615_5 gpc2425 (
      {stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205]},
      {stage1_10[14]},
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage2_13[7],stage2_12[9],stage2_11[36],stage2_10[60],stage2_9[70]}
   );
   gpc615_5 gpc2426 (
      {stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_10[15]},
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage2_13[8],stage2_12[10],stage2_11[37],stage2_10[61],stage2_9[71]}
   );
   gpc117_4 gpc2427 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[55]},
      {stage1_12[0]},
      {stage2_13[9],stage2_12[11],stage2_11[38],stage2_10[62]}
   );
   gpc117_4 gpc2428 (
      {stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_11[56]},
      {stage1_12[1]},
      {stage2_13[10],stage2_12[12],stage2_11[39],stage2_10[63]}
   );
   gpc117_4 gpc2429 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[57]},
      {stage1_12[2]},
      {stage2_13[11],stage2_12[13],stage2_11[40],stage2_10[64]}
   );
   gpc117_4 gpc2430 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage1_11[58]},
      {stage1_12[3]},
      {stage2_13[12],stage2_12[14],stage2_11[41],stage2_10[65]}
   );
   gpc117_4 gpc2431 (
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[59]},
      {stage1_12[4]},
      {stage2_13[13],stage2_12[15],stage2_11[42],stage2_10[66]}
   );
   gpc117_4 gpc2432 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57]},
      {stage1_11[60]},
      {stage1_12[5]},
      {stage2_13[14],stage2_12[16],stage2_11[43],stage2_10[67]}
   );
   gpc117_4 gpc2433 (
      {stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64]},
      {stage1_11[61]},
      {stage1_12[6]},
      {stage2_13[15],stage2_12[17],stage2_11[44],stage2_10[68]}
   );
   gpc117_4 gpc2434 (
      {stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_11[62]},
      {stage1_12[7]},
      {stage2_13[16],stage2_12[18],stage2_11[45],stage2_10[69]}
   );
   gpc117_4 gpc2435 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[63]},
      {stage1_12[8]},
      {stage2_13[17],stage2_12[19],stage2_11[46],stage2_10[70]}
   );
   gpc117_4 gpc2436 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage1_11[64]},
      {stage1_12[9]},
      {stage2_13[18],stage2_12[20],stage2_11[47],stage2_10[71]}
   );
   gpc117_4 gpc2437 (
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92]},
      {stage1_11[65]},
      {stage1_12[10]},
      {stage2_13[19],stage2_12[21],stage2_11[48],stage2_10[72]}
   );
   gpc117_4 gpc2438 (
      {stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99]},
      {stage1_11[66]},
      {stage1_12[11]},
      {stage2_13[20],stage2_12[22],stage2_11[49],stage2_10[73]}
   );
   gpc117_4 gpc2439 (
      {stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[67]},
      {stage1_12[12]},
      {stage2_13[21],stage2_12[23],stage2_11[50],stage2_10[74]}
   );
   gpc117_4 gpc2440 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_11[68]},
      {stage1_12[13]},
      {stage2_13[22],stage2_12[24],stage2_11[51],stage2_10[75]}
   );
   gpc117_4 gpc2441 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120]},
      {stage1_11[69]},
      {stage1_12[14]},
      {stage2_13[23],stage2_12[25],stage2_11[52],stage2_10[76]}
   );
   gpc117_4 gpc2442 (
      {stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125], stage1_10[126], stage1_10[127]},
      {stage1_11[70]},
      {stage1_12[15]},
      {stage2_13[24],stage2_12[26],stage2_11[53],stage2_10[77]}
   );
   gpc117_4 gpc2443 (
      {stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[71]},
      {stage1_12[16]},
      {stage2_13[25],stage2_12[27],stage2_11[54],stage2_10[78]}
   );
   gpc117_4 gpc2444 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141]},
      {stage1_11[72]},
      {stage1_12[17]},
      {stage2_13[26],stage2_12[28],stage2_11[55],stage2_10[79]}
   );
   gpc117_4 gpc2445 (
      {stage1_10[142], stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_11[73]},
      {stage1_12[18]},
      {stage2_13[27],stage2_12[29],stage2_11[56],stage2_10[80]}
   );
   gpc117_4 gpc2446 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_11[74]},
      {stage1_12[19]},
      {stage2_13[28],stage2_12[30],stage2_11[57],stage2_10[81]}
   );
   gpc606_5 gpc2447 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[0],stage2_13[29],stage2_12[31],stage2_11[58],stage2_10[82]}
   );
   gpc606_5 gpc2448 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[1],stage2_13[30],stage2_12[32],stage2_11[59],stage2_10[83]}
   );
   gpc606_5 gpc2449 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37]},
      {stage2_14[2],stage2_13[31],stage2_12[33],stage2_11[60],stage2_10[84]}
   );
   gpc606_5 gpc2450 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43]},
      {stage2_14[3],stage2_13[32],stage2_12[34],stage2_11[61],stage2_10[85]}
   );
   gpc606_5 gpc2451 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage2_14[4],stage2_13[33],stage2_12[35],stage2_11[62],stage2_10[86]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78], stage1_11[79]},
      {stage1_12[50]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[34],stage2_12[36],stage2_11[63]}
   );
   gpc615_5 gpc2453 (
      {stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_12[51]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[35],stage2_12[37],stage2_11[64]}
   );
   gpc615_5 gpc2454 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage1_12[52]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[36],stage2_12[38],stage2_11[65]}
   );
   gpc615_5 gpc2455 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[53]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[8],stage2_13[37],stage2_12[39],stage2_11[66]}
   );
   gpc615_5 gpc2456 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[54]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[9],stage2_13[38],stage2_12[40],stage2_11[67]}
   );
   gpc615_5 gpc2457 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[55]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[10],stage2_13[39],stage2_12[41],stage2_11[68]}
   );
   gpc615_5 gpc2458 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[56]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[11],stage2_13[40],stage2_12[42],stage2_11[69]}
   );
   gpc615_5 gpc2459 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[57]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[12],stage2_13[41],stage2_12[43],stage2_11[70]}
   );
   gpc615_5 gpc2460 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[58]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[13],stage2_13[42],stage2_12[44],stage2_11[71]}
   );
   gpc615_5 gpc2461 (
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124]},
      {stage1_12[59]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[14],stage2_13[43],stage2_12[45],stage2_11[72]}
   );
   gpc615_5 gpc2462 (
      {stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[60]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[15],stage2_13[44],stage2_12[46],stage2_11[73]}
   );
   gpc615_5 gpc2463 (
      {stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133], stage1_11[134]},
      {stage1_12[61]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[16],stage2_13[45],stage2_12[47],stage2_11[74]}
   );
   gpc615_5 gpc2464 (
      {stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139]},
      {stage1_12[62]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[17],stage2_13[46],stage2_12[48],stage2_11[75]}
   );
   gpc615_5 gpc2465 (
      {stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[63]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[18],stage2_13[47],stage2_12[49],stage2_11[76]}
   );
   gpc615_5 gpc2466 (
      {stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149]},
      {stage1_12[64]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[19],stage2_13[48],stage2_12[50],stage2_11[77]}
   );
   gpc615_5 gpc2467 (
      {stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154]},
      {stage1_12[65]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[20],stage2_13[49],stage2_12[51],stage2_11[78]}
   );
   gpc615_5 gpc2468 (
      {stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[66]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[21],stage2_13[50],stage2_12[52],stage2_11[79]}
   );
   gpc615_5 gpc2469 (
      {stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163], stage1_11[164]},
      {stage1_12[67]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[22],stage2_13[51],stage2_12[53],stage2_11[80]}
   );
   gpc615_5 gpc2470 (
      {stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168], stage1_11[169]},
      {stage1_12[68]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[23],stage2_13[52],stage2_12[54],stage2_11[81]}
   );
   gpc615_5 gpc2471 (
      {stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173], stage1_11[174]},
      {stage1_12[69]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[24],stage2_13[53],stage2_12[55],stage2_11[82]}
   );
   gpc615_5 gpc2472 (
      {stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178], stage1_11[179]},
      {stage1_12[70]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[25],stage2_13[54],stage2_12[56],stage2_11[83]}
   );
   gpc615_5 gpc2473 (
      {stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183], stage1_11[184]},
      {stage1_12[71]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[26],stage2_13[55],stage2_12[57],stage2_11[84]}
   );
   gpc615_5 gpc2474 (
      {stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188], stage1_11[189]},
      {stage1_12[72]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[27],stage2_13[56],stage2_12[58],stage2_11[85]}
   );
   gpc615_5 gpc2475 (
      {stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193], stage1_11[194]},
      {stage1_12[73]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[28],stage2_13[57],stage2_12[59],stage2_11[86]}
   );
   gpc615_5 gpc2476 (
      {stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198], stage1_11[199]},
      {stage1_12[74]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[29],stage2_13[58],stage2_12[60],stage2_11[87]}
   );
   gpc615_5 gpc2477 (
      {stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203], stage1_11[204]},
      {stage1_12[75]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[30],stage2_13[59],stage2_12[61],stage2_11[88]}
   );
   gpc615_5 gpc2478 (
      {stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208], stage1_11[209]},
      {stage1_12[76]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[31],stage2_13[60],stage2_12[62],stage2_11[89]}
   );
   gpc615_5 gpc2479 (
      {stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213], stage1_11[214]},
      {stage1_12[77]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[32],stage2_13[61],stage2_12[63],stage2_11[90]}
   );
   gpc615_5 gpc2480 (
      {stage1_11[215], stage1_11[216], stage1_11[217], stage1_11[218], stage1_11[219]},
      {stage1_12[78]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[33],stage2_13[62],stage2_12[64],stage2_11[91]}
   );
   gpc606_5 gpc2481 (
      {stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[29],stage2_14[34],stage2_13[63],stage2_12[65]}
   );
   gpc606_5 gpc2482 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89], stage1_12[90]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[30],stage2_14[35],stage2_13[64],stage2_12[66]}
   );
   gpc606_5 gpc2483 (
      {stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95], stage1_12[96]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[31],stage2_14[36],stage2_13[65],stage2_12[67]}
   );
   gpc606_5 gpc2484 (
      {stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[32],stage2_14[37],stage2_13[66],stage2_12[68]}
   );
   gpc606_5 gpc2485 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[33],stage2_14[38],stage2_13[67],stage2_12[69]}
   );
   gpc606_5 gpc2486 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[34],stage2_14[39],stage2_13[68],stage2_12[70]}
   );
   gpc606_5 gpc2487 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[35],stage2_14[40],stage2_13[69],stage2_12[71]}
   );
   gpc606_5 gpc2488 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[36],stage2_14[41],stage2_13[70],stage2_12[72]}
   );
   gpc606_5 gpc2489 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[37],stage2_14[42],stage2_13[71],stage2_12[73]}
   );
   gpc606_5 gpc2490 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[38],stage2_14[43],stage2_13[72],stage2_12[74]}
   );
   gpc606_5 gpc2491 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[39],stage2_14[44],stage2_13[73],stage2_12[75]}
   );
   gpc606_5 gpc2492 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[40],stage2_14[45],stage2_13[74],stage2_12[76]}
   );
   gpc606_5 gpc2493 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[41],stage2_14[46],stage2_13[75],stage2_12[77]}
   );
   gpc606_5 gpc2494 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[42],stage2_14[47],stage2_13[76],stage2_12[78]}
   );
   gpc606_5 gpc2495 (
      {stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[43],stage2_14[48],stage2_13[77],stage2_12[79]}
   );
   gpc606_5 gpc2496 (
      {stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[44],stage2_14[49],stage2_13[78],stage2_12[80]}
   );
   gpc606_5 gpc2497 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[45],stage2_14[50],stage2_13[79],stage2_12[81]}
   );
   gpc606_5 gpc2498 (
      {stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[46],stage2_14[51],stage2_13[80],stage2_12[82]}
   );
   gpc606_5 gpc2499 (
      {stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[47],stage2_14[52],stage2_13[81],stage2_12[83]}
   );
   gpc606_5 gpc2500 (
      {stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[48],stage2_14[53],stage2_13[82],stage2_12[84]}
   );
   gpc606_5 gpc2501 (
      {stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[49],stage2_14[54],stage2_13[83],stage2_12[85]}
   );
   gpc606_5 gpc2502 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209], stage1_12[210]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[50],stage2_14[55],stage2_13[84],stage2_12[86]}
   );
   gpc606_5 gpc2503 (
      {stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214], stage1_12[215], stage1_12[216]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[51],stage2_14[56],stage2_13[85],stage2_12[87]}
   );
   gpc606_5 gpc2504 (
      {stage1_12[217], stage1_12[218], stage1_12[219], stage1_12[220], stage1_12[221], stage1_12[222]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[52],stage2_14[57],stage2_13[86],stage2_12[88]}
   );
   gpc606_5 gpc2505 (
      {stage1_12[223], stage1_12[224], stage1_12[225], stage1_12[226], stage1_12[227], stage1_12[228]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[53],stage2_14[58],stage2_13[87],stage2_12[89]}
   );
   gpc606_5 gpc2506 (
      {stage1_12[229], stage1_12[230], stage1_12[231], stage1_12[232], stage1_12[233], stage1_12[234]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[54],stage2_14[59],stage2_13[88],stage2_12[90]}
   );
   gpc606_5 gpc2507 (
      {stage1_12[235], stage1_12[236], stage1_12[237], stage1_12[238], stage1_12[239], stage1_12[240]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[55],stage2_14[60],stage2_13[89],stage2_12[91]}
   );
   gpc606_5 gpc2508 (
      {stage1_12[241], stage1_12[242], stage1_12[243], stage1_12[244], stage1_12[245], stage1_12[246]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[56],stage2_14[61],stage2_13[90],stage2_12[92]}
   );
   gpc606_5 gpc2509 (
      {stage1_12[247], stage1_12[248], stage1_12[249], stage1_12[250], stage1_12[251], stage1_12[252]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[57],stage2_14[62],stage2_13[91],stage2_12[93]}
   );
   gpc606_5 gpc2510 (
      {stage1_12[253], stage1_12[254], stage1_12[255], stage1_12[256], stage1_12[257], stage1_12[258]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[58],stage2_14[63],stage2_13[92],stage2_12[94]}
   );
   gpc606_5 gpc2511 (
      {stage1_12[259], stage1_12[260], stage1_12[261], stage1_12[262], stage1_12[263], stage1_12[264]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[59],stage2_14[64],stage2_13[93],stage2_12[95]}
   );
   gpc606_5 gpc2512 (
      {stage1_12[265], stage1_12[266], stage1_12[267], stage1_12[268], stage1_12[269], stage1_12[270]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[60],stage2_14[65],stage2_13[94],stage2_12[96]}
   );
   gpc606_5 gpc2513 (
      {stage1_12[271], stage1_12[272], stage1_12[273], stage1_12[274], stage1_12[275], stage1_12[276]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[61],stage2_14[66],stage2_13[95],stage2_12[97]}
   );
   gpc606_5 gpc2514 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[33],stage2_15[62],stage2_14[67],stage2_13[96]}
   );
   gpc615_5 gpc2515 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[198]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[34],stage2_15[63],stage2_14[68],stage2_13[97]}
   );
   gpc615_5 gpc2516 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[199]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[35],stage2_15[64],stage2_14[69],stage2_13[98]}
   );
   gpc615_5 gpc2517 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[200]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[36],stage2_15[65],stage2_14[70],stage2_13[99]}
   );
   gpc615_5 gpc2518 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[201]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[37],stage2_15[66],stage2_14[71],stage2_13[100]}
   );
   gpc615_5 gpc2519 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[202]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[38],stage2_15[67],stage2_14[72],stage2_13[101]}
   );
   gpc615_5 gpc2520 (
      {stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207]},
      {stage1_15[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[6],stage2_16[39],stage2_15[68],stage2_14[73]}
   );
   gpc615_5 gpc2521 (
      {stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211], stage1_14[212]},
      {stage1_15[37]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[7],stage2_16[40],stage2_15[69],stage2_14[74]}
   );
   gpc615_5 gpc2522 (
      {stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216], stage1_14[217]},
      {stage1_15[38]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[8],stage2_16[41],stage2_15[70],stage2_14[75]}
   );
   gpc615_5 gpc2523 (
      {stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221], stage1_14[222]},
      {stage1_15[39]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[9],stage2_16[42],stage2_15[71],stage2_14[76]}
   );
   gpc615_5 gpc2524 (
      {stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226], stage1_14[227]},
      {stage1_15[40]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[10],stage2_16[43],stage2_15[72],stage2_14[77]}
   );
   gpc615_5 gpc2525 (
      {stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231], stage1_14[232]},
      {stage1_15[41]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[11],stage2_16[44],stage2_15[73],stage2_14[78]}
   );
   gpc615_5 gpc2526 (
      {stage1_14[233], stage1_14[234], stage1_14[235], stage1_14[236], stage1_14[237]},
      {stage1_15[42]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[12],stage2_16[45],stage2_15[74],stage2_14[79]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[42]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[46],stage2_15[75]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52]},
      {stage1_16[43]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[47],stage2_15[76]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[53], stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57]},
      {stage1_16[44]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[48],stage2_15[77]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62]},
      {stage1_16[45]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[49],stage2_15[78]}
   );
   gpc615_5 gpc2531 (
      {stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_16[46]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[50],stage2_15[79]}
   );
   gpc615_5 gpc2532 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72]},
      {stage1_16[47]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[51],stage2_15[80]}
   );
   gpc615_5 gpc2533 (
      {stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[48]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[52],stage2_15[81]}
   );
   gpc615_5 gpc2534 (
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82]},
      {stage1_16[49]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[53],stage2_15[82]}
   );
   gpc615_5 gpc2535 (
      {stage1_15[83], stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87]},
      {stage1_16[50]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[54],stage2_15[83]}
   );
   gpc615_5 gpc2536 (
      {stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91], stage1_15[92]},
      {stage1_16[51]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[55],stage2_15[84]}
   );
   gpc615_5 gpc2537 (
      {stage1_15[93], stage1_15[94], stage1_15[95], stage1_15[96], stage1_15[97]},
      {stage1_16[52]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[56],stage2_15[85]}
   );
   gpc615_5 gpc2538 (
      {stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101], stage1_15[102]},
      {stage1_16[53]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[57],stage2_15[86]}
   );
   gpc615_5 gpc2539 (
      {stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[54]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[19],stage2_17[25],stage2_16[58],stage2_15[87]}
   );
   gpc615_5 gpc2540 (
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112]},
      {stage1_16[55]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[20],stage2_17[26],stage2_16[59],stage2_15[88]}
   );
   gpc615_5 gpc2541 (
      {stage1_15[113], stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117]},
      {stage1_16[56]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[21],stage2_17[27],stage2_16[60],stage2_15[89]}
   );
   gpc615_5 gpc2542 (
      {stage1_15[118], stage1_15[119], stage1_15[120], stage1_15[121], stage1_15[122]},
      {stage1_16[57]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[22],stage2_17[28],stage2_16[61],stage2_15[90]}
   );
   gpc615_5 gpc2543 (
      {stage1_15[123], stage1_15[124], stage1_15[125], stage1_15[126], stage1_15[127]},
      {stage1_16[58]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[23],stage2_17[29],stage2_16[62],stage2_15[91]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[59], stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[24],stage2_17[30],stage2_16[63]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[25],stage2_17[31],stage2_16[64]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[26],stage2_17[32],stage2_16[65]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[27],stage2_17[33],stage2_16[66]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[28],stage2_17[34],stage2_16[67]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[89], stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[29],stage2_17[35],stage2_16[68]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[95], stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[30],stage2_17[36],stage2_16[69]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[101], stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[31],stage2_17[37],stage2_16[70]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[107], stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[32],stage2_17[38],stage2_16[71]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[113], stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[33],stage2_17[39],stage2_16[72]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[119], stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[34],stage2_17[40],stage2_16[73]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[125], stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[35],stage2_17[41],stage2_16[74]}
   );
   gpc606_5 gpc2556 (
      {stage1_16[131], stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[36],stage2_17[42],stage2_16[75]}
   );
   gpc606_5 gpc2557 (
      {stage1_16[137], stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[37],stage2_17[43],stage2_16[76]}
   );
   gpc606_5 gpc2558 (
      {stage1_16[143], stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[38],stage2_17[44],stage2_16[77]}
   );
   gpc606_5 gpc2559 (
      {stage1_16[149], stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[39],stage2_17[45],stage2_16[78]}
   );
   gpc606_5 gpc2560 (
      {stage1_16[155], stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[40],stage2_17[46],stage2_16[79]}
   );
   gpc606_5 gpc2561 (
      {stage1_16[161], stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[41],stage2_17[47],stage2_16[80]}
   );
   gpc606_5 gpc2562 (
      {stage1_16[167], stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[42],stage2_17[48],stage2_16[81]}
   );
   gpc606_5 gpc2563 (
      {stage1_16[173], stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[43],stage2_17[49],stage2_16[82]}
   );
   gpc606_5 gpc2564 (
      {stage1_16[179], stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[44],stage2_17[50],stage2_16[83]}
   );
   gpc606_5 gpc2565 (
      {stage1_16[185], stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[45],stage2_17[51],stage2_16[84]}
   );
   gpc606_5 gpc2566 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[46],stage2_17[52],stage2_16[85]}
   );
   gpc606_5 gpc2567 (
      {stage1_16[197], stage1_16[198], stage1_16[199], stage1_16[200], stage1_16[201], stage1_16[202]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[47],stage2_17[53],stage2_16[86]}
   );
   gpc606_5 gpc2568 (
      {stage1_16[203], stage1_16[204], stage1_16[205], stage1_16[206], stage1_16[207], stage1_16[208]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[48],stage2_17[54],stage2_16[87]}
   );
   gpc606_5 gpc2569 (
      {stage1_16[209], stage1_16[210], stage1_16[211], stage1_16[212], stage1_16[213], stage1_16[214]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[49],stage2_17[55],stage2_16[88]}
   );
   gpc606_5 gpc2570 (
      {stage1_16[215], stage1_16[216], stage1_16[217], stage1_16[218], stage1_16[219], stage1_16[220]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[50],stage2_17[56],stage2_16[89]}
   );
   gpc606_5 gpc2571 (
      {stage1_16[221], stage1_16[222], stage1_16[223], stage1_16[224], stage1_16[225], stage1_16[226]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[51],stage2_17[57],stage2_16[90]}
   );
   gpc606_5 gpc2572 (
      {stage1_16[227], stage1_16[228], stage1_16[229], stage1_16[230], stage1_16[231], stage1_16[232]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[52],stage2_17[58],stage2_16[91]}
   );
   gpc606_5 gpc2573 (
      {stage1_16[233], stage1_16[234], stage1_16[235], stage1_16[236], stage1_16[237], stage1_16[238]},
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage2_20[29],stage2_19[46],stage2_18[53],stage2_17[59],stage2_16[92]}
   );
   gpc606_5 gpc2574 (
      {stage1_16[239], stage1_16[240], stage1_16[241], stage1_16[242], stage1_16[243], stage1_16[244]},
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage2_20[30],stage2_19[47],stage2_18[54],stage2_17[60],stage2_16[93]}
   );
   gpc606_5 gpc2575 (
      {stage1_16[245], stage1_16[246], stage1_16[247], stage1_16[248], stage1_16[249], stage1_16[250]},
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190], stage1_18[191]},
      {stage2_20[31],stage2_19[48],stage2_18[55],stage2_17[61],stage2_16[94]}
   );
   gpc606_5 gpc2576 (
      {stage1_16[251], stage1_16[252], stage1_16[253], stage1_16[254], stage1_16[255], stage1_16[256]},
      {stage1_18[192], stage1_18[193], stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197]},
      {stage2_20[32],stage2_19[49],stage2_18[56],stage2_17[62],stage2_16[95]}
   );
   gpc606_5 gpc2577 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[33],stage2_19[50],stage2_18[57],stage2_17[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[34],stage2_19[51],stage2_18[58],stage2_17[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[35],stage2_19[52],stage2_18[59],stage2_17[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[36],stage2_19[53],stage2_18[60],stage2_17[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[37],stage2_19[54],stage2_18[61],stage2_17[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[38],stage2_19[55],stage2_18[62],stage2_17[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[39],stage2_19[56],stage2_18[63],stage2_17[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[40],stage2_19[57],stage2_18[64],stage2_17[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[41],stage2_19[58],stage2_18[65],stage2_17[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[42],stage2_19[59],stage2_18[66],stage2_17[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[43],stage2_19[60],stage2_18[67],stage2_17[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[44],stage2_19[61],stage2_18[68],stage2_17[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[45],stage2_19[62],stage2_18[69],stage2_17[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[46],stage2_19[63],stage2_18[70],stage2_17[76]}
   );
   gpc606_5 gpc2591 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[47],stage2_19[64],stage2_18[71],stage2_17[77]}
   );
   gpc606_5 gpc2592 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[48],stage2_19[65],stage2_18[72],stage2_17[78]}
   );
   gpc606_5 gpc2593 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[49],stage2_19[66],stage2_18[73],stage2_17[79]}
   );
   gpc606_5 gpc2594 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[50],stage2_19[67],stage2_18[74],stage2_17[80]}
   );
   gpc606_5 gpc2595 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[51],stage2_19[68],stage2_18[75],stage2_17[81]}
   );
   gpc606_5 gpc2596 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[52],stage2_19[69],stage2_18[76],stage2_17[82]}
   );
   gpc606_5 gpc2597 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[53],stage2_19[70],stage2_18[77],stage2_17[83]}
   );
   gpc606_5 gpc2598 (
      {stage1_17[228], stage1_17[229], stage1_17[230], stage1_17[231], stage1_17[232], stage1_17[233]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[54],stage2_19[71],stage2_18[78],stage2_17[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[22],stage2_20[55],stage2_19[72]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[23],stage2_20[56],stage2_19[73]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[24],stage2_20[57],stage2_19[74]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[147], stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[25],stage2_20[58],stage2_19[75]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155], stage1_19[156]},
      {stage1_20[4]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[26],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage1_20[5]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[27],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166]},
      {stage1_20[6]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[6],stage2_21[28],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171]},
      {stage1_20[7]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[7],stage2_21[29],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175], stage1_19[176]},
      {stage1_20[8]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[8],stage2_21[30],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180], stage1_19[181]},
      {stage1_20[9]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[9],stage2_21[31],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185], stage1_19[186]},
      {stage1_20[10]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[10],stage2_21[32],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2610 (
      {stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage1_20[11]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[11],stage2_21[33],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2611 (
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196]},
      {stage1_20[12]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[12],stage2_21[34],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2612 (
      {stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201]},
      {stage1_20[13]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[13],stage2_21[35],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2613 (
      {stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205], stage1_19[206]},
      {stage1_20[14]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[14],stage2_21[36],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2614 (
      {stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210], stage1_19[211]},
      {stage1_20[15]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[15],stage2_21[37],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2615 (
      {stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215], stage1_19[216]},
      {stage1_20[16]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[16],stage2_21[38],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2616 (
      {stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage1_20[17]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[17],stage2_21[39],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2617 (
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226]},
      {stage1_20[18]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[18],stage2_21[40],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2618 (
      {stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230], stage1_19[231]},
      {stage1_20[19]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[19],stage2_21[41],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2619 (
      {stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235], stage1_19[236]},
      {stage1_20[20]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[20],stage2_21[42],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2620 (
      {stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240], stage1_19[241]},
      {stage1_20[21]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[21],stage2_21[43],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2621 (
      {stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245], stage1_19[246]},
      {stage1_20[22]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[22],stage2_21[44],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2622 (
      {stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250], stage1_19[251]},
      {stage1_20[23]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[23],stage2_21[45],stage2_20[78],stage2_19[95]}
   );
   gpc615_5 gpc2623 (
      {stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255], stage1_19[256]},
      {stage1_20[24]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[24],stage2_21[46],stage2_20[79],stage2_19[96]}
   );
   gpc615_5 gpc2624 (
      {stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260], stage1_19[261]},
      {stage1_20[25]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[25],stage2_21[47],stage2_20[80],stage2_19[97]}
   );
   gpc615_5 gpc2625 (
      {stage1_19[262], stage1_19[263], stage1_19[264], stage1_19[265], stage1_19[266]},
      {stage1_20[26]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[26],stage2_21[48],stage2_20[81],stage2_19[98]}
   );
   gpc615_5 gpc2626 (
      {stage1_19[267], stage1_19[268], stage1_19[269], stage1_19[270], stage1_19[271]},
      {stage1_20[27]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[27],stage2_21[49],stage2_20[82],stage2_19[99]}
   );
   gpc615_5 gpc2627 (
      {stage1_19[272], stage1_19[273], stage1_19[274], stage1_19[275], stage1_19[276]},
      {stage1_20[28]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[28],stage2_21[50],stage2_20[83],stage2_19[100]}
   );
   gpc615_5 gpc2628 (
      {stage1_19[277], stage1_19[278], stage1_19[279], stage1_19[280], stage1_19[281]},
      {stage1_20[29]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[29],stage2_21[51],stage2_20[84],stage2_19[101]}
   );
   gpc615_5 gpc2629 (
      {stage1_19[282], stage1_19[283], stage1_19[284], stage1_19[285], stage1_19[286]},
      {stage1_20[30]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[30],stage2_21[52],stage2_20[85],stage2_19[102]}
   );
   gpc615_5 gpc2630 (
      {stage1_19[287], stage1_19[288], stage1_19[289], stage1_19[290], stage1_19[291]},
      {stage1_20[31]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[31],stage2_21[53],stage2_20[86],stage2_19[103]}
   );
   gpc623_5 gpc2631 (
      {stage1_19[292], stage1_19[293], stage1_19[294]},
      {stage1_20[32], stage1_20[33]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[32],stage2_21[54],stage2_20[87],stage2_19[104]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[34], stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[33],stage2_22[33],stage2_21[55],stage2_20[88]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[40], stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[34],stage2_22[34],stage2_21[56],stage2_20[89]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[46], stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[35],stage2_22[35],stage2_21[57],stage2_20[90]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[52], stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[36],stage2_22[36],stage2_21[58],stage2_20[91]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[58], stage1_20[59], stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[37],stage2_22[37],stage2_21[59],stage2_20[92]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[64], stage1_20[65], stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[38],stage2_22[38],stage2_21[60],stage2_20[93]}
   );
   gpc606_5 gpc2638 (
      {stage1_20[70], stage1_20[71], stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[39],stage2_22[39],stage2_21[61],stage2_20[94]}
   );
   gpc606_5 gpc2639 (
      {stage1_20[76], stage1_20[77], stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[40],stage2_22[40],stage2_21[62],stage2_20[95]}
   );
   gpc606_5 gpc2640 (
      {stage1_20[82], stage1_20[83], stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[41],stage2_22[41],stage2_21[63],stage2_20[96]}
   );
   gpc606_5 gpc2641 (
      {stage1_20[88], stage1_20[89], stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[42],stage2_22[42],stage2_21[64],stage2_20[97]}
   );
   gpc606_5 gpc2642 (
      {stage1_20[94], stage1_20[95], stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[43],stage2_22[43],stage2_21[65],stage2_20[98]}
   );
   gpc606_5 gpc2643 (
      {stage1_20[100], stage1_20[101], stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[44],stage2_22[44],stage2_21[66],stage2_20[99]}
   );
   gpc606_5 gpc2644 (
      {stage1_20[106], stage1_20[107], stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[45],stage2_22[45],stage2_21[67],stage2_20[100]}
   );
   gpc606_5 gpc2645 (
      {stage1_20[112], stage1_20[113], stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[46],stage2_22[46],stage2_21[68],stage2_20[101]}
   );
   gpc606_5 gpc2646 (
      {stage1_20[118], stage1_20[119], stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[47],stage2_22[47],stage2_21[69],stage2_20[102]}
   );
   gpc606_5 gpc2647 (
      {stage1_20[124], stage1_20[125], stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[48],stage2_22[48],stage2_21[70],stage2_20[103]}
   );
   gpc606_5 gpc2648 (
      {stage1_20[130], stage1_20[131], stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[49],stage2_22[49],stage2_21[71],stage2_20[104]}
   );
   gpc606_5 gpc2649 (
      {stage1_20[136], stage1_20[137], stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[50],stage2_22[50],stage2_21[72],stage2_20[105]}
   );
   gpc606_5 gpc2650 (
      {stage1_20[142], stage1_20[143], stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[51],stage2_22[51],stage2_21[73],stage2_20[106]}
   );
   gpc606_5 gpc2651 (
      {stage1_20[148], stage1_20[149], stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[52],stage2_22[52],stage2_21[74],stage2_20[107]}
   );
   gpc606_5 gpc2652 (
      {stage1_20[154], stage1_20[155], stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[53],stage2_22[53],stage2_21[75],stage2_20[108]}
   );
   gpc606_5 gpc2653 (
      {stage1_20[160], stage1_20[161], stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[54],stage2_22[54],stage2_21[76],stage2_20[109]}
   );
   gpc606_5 gpc2654 (
      {stage1_20[166], stage1_20[167], stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[55],stage2_22[55],stage2_21[77],stage2_20[110]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142]},
      {stage1_23[0]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[0],stage2_24[23],stage2_23[56],stage2_22[56]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[143], stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147]},
      {stage1_23[1]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[1],stage2_24[24],stage2_23[57],stage2_22[57]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[148], stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152]},
      {stage1_23[2]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[2],stage2_24[25],stage2_23[58],stage2_22[58]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[153], stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157]},
      {stage1_23[3]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[3],stage2_24[26],stage2_23[59],stage2_22[59]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162]},
      {stage1_23[4]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[4],stage2_24[27],stage2_23[60],stage2_22[60]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage1_23[5]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[5],stage2_24[28],stage2_23[61],stage2_22[61]}
   );
   gpc615_5 gpc2661 (
      {stage1_22[168], stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172]},
      {stage1_23[6]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[6],stage2_24[29],stage2_23[62],stage2_22[62]}
   );
   gpc615_5 gpc2662 (
      {stage1_22[173], stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177]},
      {stage1_23[7]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[7],stage2_24[30],stage2_23[63],stage2_22[63]}
   );
   gpc615_5 gpc2663 (
      {stage1_22[178], stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182]},
      {stage1_23[8]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[8],stage2_24[31],stage2_23[64],stage2_22[64]}
   );
   gpc615_5 gpc2664 (
      {stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187]},
      {stage1_23[9]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[9],stage2_24[32],stage2_23[65],stage2_22[65]}
   );
   gpc615_5 gpc2665 (
      {stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_23[10]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[10],stage2_24[33],stage2_23[66],stage2_22[66]}
   );
   gpc615_5 gpc2666 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[11]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[11],stage2_24[34],stage2_23[67],stage2_22[67]}
   );
   gpc615_5 gpc2667 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[12]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[12],stage2_24[35],stage2_23[68],stage2_22[68]}
   );
   gpc615_5 gpc2668 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[13]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[13],stage2_24[36],stage2_23[69],stage2_22[69]}
   );
   gpc615_5 gpc2669 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[14]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[14],stage2_24[37],stage2_23[70],stage2_22[70]}
   );
   gpc615_5 gpc2670 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[15]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[15],stage2_24[38],stage2_23[71],stage2_22[71]}
   );
   gpc615_5 gpc2671 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[16]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[16],stage2_24[39],stage2_23[72],stage2_22[72]}
   );
   gpc615_5 gpc2672 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[17]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[17],stage2_24[40],stage2_23[73],stage2_22[73]}
   );
   gpc615_5 gpc2673 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[18]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[18],stage2_24[41],stage2_23[74],stage2_22[74]}
   );
   gpc615_5 gpc2674 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[19]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[19],stage2_24[42],stage2_23[75],stage2_22[75]}
   );
   gpc615_5 gpc2675 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[20]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[20],stage2_24[43],stage2_23[76],stage2_22[76]}
   );
   gpc615_5 gpc2676 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[21]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[21],stage2_24[44],stage2_23[77],stage2_22[77]}
   );
   gpc615_5 gpc2677 (
      {stage1_22[248], stage1_22[249], stage1_22[250], 1'b0, 1'b0},
      {stage1_23[22]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[22],stage2_24[45],stage2_23[78],stage2_22[78]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[23], stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27]},
      {stage1_24[138]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[23],stage2_25[23],stage2_24[46],stage2_23[79]}
   );
   gpc615_5 gpc2679 (
      {stage1_23[28], stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32]},
      {stage1_24[139]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[24],stage2_25[24],stage2_24[47],stage2_23[80]}
   );
   gpc615_5 gpc2680 (
      {stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36], stage1_23[37]},
      {stage1_24[140]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[25],stage2_25[25],stage2_24[48],stage2_23[81]}
   );
   gpc615_5 gpc2681 (
      {stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_24[141]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[26],stage2_25[26],stage2_24[49],stage2_23[82]}
   );
   gpc615_5 gpc2682 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[142]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[27],stage2_25[27],stage2_24[50],stage2_23[83]}
   );
   gpc615_5 gpc2683 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52]},
      {stage1_24[143]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[28],stage2_25[28],stage2_24[51],stage2_23[84]}
   );
   gpc615_5 gpc2684 (
      {stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57]},
      {stage1_24[144]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[29],stage2_25[29],stage2_24[52],stage2_23[85]}
   );
   gpc615_5 gpc2685 (
      {stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_24[145]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[30],stage2_25[30],stage2_24[53],stage2_23[86]}
   );
   gpc615_5 gpc2686 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67]},
      {stage1_24[146]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[31],stage2_25[31],stage2_24[54],stage2_23[87]}
   );
   gpc615_5 gpc2687 (
      {stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_24[147]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[32],stage2_25[32],stage2_24[55],stage2_23[88]}
   );
   gpc615_5 gpc2688 (
      {stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_24[148]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[33],stage2_25[33],stage2_24[56],stage2_23[89]}
   );
   gpc615_5 gpc2689 (
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82]},
      {stage1_24[149]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[34],stage2_25[34],stage2_24[57],stage2_23[90]}
   );
   gpc615_5 gpc2690 (
      {stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87]},
      {stage1_24[150]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[35],stage2_25[35],stage2_24[58],stage2_23[91]}
   );
   gpc615_5 gpc2691 (
      {stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_24[151]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[36],stage2_25[36],stage2_24[59],stage2_23[92]}
   );
   gpc615_5 gpc2692 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97]},
      {stage1_24[152]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[37],stage2_25[37],stage2_24[60],stage2_23[93]}
   );
   gpc615_5 gpc2693 (
      {stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_24[153]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[38],stage2_25[38],stage2_24[61],stage2_23[94]}
   );
   gpc615_5 gpc2694 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage1_24[154]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[39],stage2_25[39],stage2_24[62],stage2_23[95]}
   );
   gpc615_5 gpc2695 (
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112]},
      {stage1_24[155]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[40],stage2_25[40],stage2_24[63],stage2_23[96]}
   );
   gpc615_5 gpc2696 (
      {stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117]},
      {stage1_24[156]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[41],stage2_25[41],stage2_24[64],stage2_23[97]}
   );
   gpc615_5 gpc2697 (
      {stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_24[157]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[42],stage2_25[42],stage2_24[65],stage2_23[98]}
   );
   gpc615_5 gpc2698 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127]},
      {stage1_24[158]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[43],stage2_25[43],stage2_24[66],stage2_23[99]}
   );
   gpc615_5 gpc2699 (
      {stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132]},
      {stage1_24[159]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[44],stage2_25[44],stage2_24[67],stage2_23[100]}
   );
   gpc615_5 gpc2700 (
      {stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage1_24[160]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[45],stage2_25[45],stage2_24[68],stage2_23[101]}
   );
   gpc615_5 gpc2701 (
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142]},
      {stage1_24[161]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[46],stage2_25[46],stage2_24[69],stage2_23[102]}
   );
   gpc615_5 gpc2702 (
      {stage1_23[143], stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147]},
      {stage1_24[162]},
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage2_27[24],stage2_26[47],stage2_25[47],stage2_24[70],stage2_23[103]}
   );
   gpc615_5 gpc2703 (
      {stage1_23[148], stage1_23[149], stage1_23[150], stage1_23[151], stage1_23[152]},
      {stage1_24[163]},
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage2_27[25],stage2_26[48],stage2_25[48],stage2_24[71],stage2_23[104]}
   );
   gpc615_5 gpc2704 (
      {stage1_23[153], stage1_23[154], stage1_23[155], stage1_23[156], stage1_23[157]},
      {stage1_24[164]},
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage2_27[26],stage2_26[49],stage2_25[49],stage2_24[72],stage2_23[105]}
   );
   gpc615_5 gpc2705 (
      {stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161], stage1_23[162]},
      {stage1_24[165]},
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage2_27[27],stage2_26[50],stage2_25[50],stage2_24[73],stage2_23[106]}
   );
   gpc615_5 gpc2706 (
      {stage1_23[163], stage1_23[164], stage1_23[165], stage1_23[166], stage1_23[167]},
      {stage1_24[166]},
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage2_27[28],stage2_26[51],stage2_25[51],stage2_24[74],stage2_23[107]}
   );
   gpc615_5 gpc2707 (
      {stage1_23[168], stage1_23[169], stage1_23[170], stage1_23[171], stage1_23[172]},
      {stage1_24[167]},
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage2_27[29],stage2_26[52],stage2_25[52],stage2_24[75],stage2_23[108]}
   );
   gpc615_5 gpc2708 (
      {stage1_23[173], stage1_23[174], stage1_23[175], stage1_23[176], stage1_23[177]},
      {stage1_24[168]},
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage2_27[30],stage2_26[53],stage2_25[53],stage2_24[76],stage2_23[109]}
   );
   gpc615_5 gpc2709 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[186]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[31],stage2_26[54],stage2_25[54],stage2_24[77]}
   );
   gpc615_5 gpc2710 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[187]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[32],stage2_26[55],stage2_25[55],stage2_24[78]}
   );
   gpc615_5 gpc2711 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[188]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[33],stage2_26[56],stage2_25[56],stage2_24[79]}
   );
   gpc615_5 gpc2712 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[189]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[34],stage2_26[57],stage2_25[57],stage2_24[80]}
   );
   gpc615_5 gpc2713 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[190]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[35],stage2_26[58],stage2_25[58],stage2_24[81]}
   );
   gpc606_5 gpc2714 (
      {stage1_25[191], stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[5],stage2_27[36],stage2_26[59],stage2_25[59]}
   );
   gpc606_5 gpc2715 (
      {stage1_25[197], stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[6],stage2_27[37],stage2_26[60],stage2_25[60]}
   );
   gpc606_5 gpc2716 (
      {stage1_25[203], stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[7],stage2_27[38],stage2_26[61],stage2_25[61]}
   );
   gpc615_5 gpc2717 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34]},
      {stage1_27[18]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[3],stage2_28[8],stage2_27[39],stage2_26[62]}
   );
   gpc615_5 gpc2718 (
      {stage1_26[35], stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39]},
      {stage1_27[19]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[4],stage2_28[9],stage2_27[40],stage2_26[63]}
   );
   gpc615_5 gpc2719 (
      {stage1_26[40], stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44]},
      {stage1_27[20]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[5],stage2_28[10],stage2_27[41],stage2_26[64]}
   );
   gpc615_5 gpc2720 (
      {stage1_26[45], stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49]},
      {stage1_27[21]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[6],stage2_28[11],stage2_27[42],stage2_26[65]}
   );
   gpc615_5 gpc2721 (
      {stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54]},
      {stage1_27[22]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[7],stage2_28[12],stage2_27[43],stage2_26[66]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage1_27[23]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[8],stage2_28[13],stage2_27[44],stage2_26[67]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64]},
      {stage1_27[24]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[9],stage2_28[14],stage2_27[45],stage2_26[68]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69]},
      {stage1_27[25]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[10],stage2_28[15],stage2_27[46],stage2_26[69]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74]},
      {stage1_27[26]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[11],stage2_28[16],stage2_27[47],stage2_26[70]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[75], stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79]},
      {stage1_27[27]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[12],stage2_28[17],stage2_27[48],stage2_26[71]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84]},
      {stage1_27[28]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[13],stage2_28[18],stage2_27[49],stage2_26[72]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage1_27[29]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[14],stage2_28[19],stage2_27[50],stage2_26[73]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94]},
      {stage1_27[30]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[15],stage2_28[20],stage2_27[51],stage2_26[74]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[95], stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99]},
      {stage1_27[31]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[16],stage2_28[21],stage2_27[52],stage2_26[75]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[100], stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104]},
      {stage1_27[32]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[17],stage2_28[22],stage2_27[53],stage2_26[76]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[105], stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109]},
      {stage1_27[33]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[18],stage2_28[23],stage2_27[54],stage2_26[77]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114]},
      {stage1_27[34]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[19],stage2_28[24],stage2_27[55],stage2_26[78]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage1_27[35]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[20],stage2_28[25],stage2_27[56],stage2_26[79]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124]},
      {stage1_27[36]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[21],stage2_28[26],stage2_27[57],stage2_26[80]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[125], stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129]},
      {stage1_27[37]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[22],stage2_28[27],stage2_27[58],stage2_26[81]}
   );
   gpc615_5 gpc2737 (
      {stage1_26[130], stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134]},
      {stage1_27[38]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[23],stage2_28[28],stage2_27[59],stage2_26[82]}
   );
   gpc615_5 gpc2738 (
      {stage1_26[135], stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139]},
      {stage1_27[39]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[24],stage2_28[29],stage2_27[60],stage2_26[83]}
   );
   gpc615_5 gpc2739 (
      {stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144]},
      {stage1_27[40]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[25],stage2_28[30],stage2_27[61],stage2_26[84]}
   );
   gpc615_5 gpc2740 (
      {stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage1_27[41]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[26],stage2_28[31],stage2_27[62],stage2_26[85]}
   );
   gpc615_5 gpc2741 (
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154]},
      {stage1_27[42]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[27],stage2_28[32],stage2_27[63],stage2_26[86]}
   );
   gpc615_5 gpc2742 (
      {stage1_26[155], stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159]},
      {stage1_27[43]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[28],stage2_28[33],stage2_27[64],stage2_26[87]}
   );
   gpc615_5 gpc2743 (
      {stage1_26[160], stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164]},
      {stage1_27[44]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[29],stage2_28[34],stage2_27[65],stage2_26[88]}
   );
   gpc615_5 gpc2744 (
      {stage1_26[165], stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169]},
      {stage1_27[45]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[30],stage2_28[35],stage2_27[66],stage2_26[89]}
   );
   gpc615_5 gpc2745 (
      {stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174]},
      {stage1_27[46]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[31],stage2_28[36],stage2_27[67],stage2_26[90]}
   );
   gpc615_5 gpc2746 (
      {stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage1_27[47]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[32],stage2_28[37],stage2_27[68],stage2_26[91]}
   );
   gpc615_5 gpc2747 (
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184]},
      {stage1_27[48]},
      {stage1_28[180], stage1_28[181], stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185]},
      {stage2_30[30],stage2_29[33],stage2_28[38],stage2_27[69],stage2_26[92]}
   );
   gpc615_5 gpc2748 (
      {stage1_26[185], stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189]},
      {stage1_27[49]},
      {stage1_28[186], stage1_28[187], stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191]},
      {stage2_30[31],stage2_29[34],stage2_28[39],stage2_27[70],stage2_26[93]}
   );
   gpc615_5 gpc2749 (
      {stage1_26[190], stage1_26[191], stage1_26[192], stage1_26[193], stage1_26[194]},
      {stage1_27[50]},
      {stage1_28[192], stage1_28[193], stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197]},
      {stage2_30[32],stage2_29[35],stage2_28[40],stage2_27[71],stage2_26[94]}
   );
   gpc615_5 gpc2750 (
      {stage1_26[195], stage1_26[196], stage1_26[197], stage1_26[198], stage1_26[199]},
      {stage1_27[51]},
      {stage1_28[198], stage1_28[199], stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203]},
      {stage2_30[33],stage2_29[36],stage2_28[41],stage2_27[72],stage2_26[95]}
   );
   gpc615_5 gpc2751 (
      {stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203], stage1_26[204]},
      {stage1_27[52]},
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage2_30[34],stage2_29[37],stage2_28[42],stage2_27[73],stage2_26[96]}
   );
   gpc615_5 gpc2752 (
      {stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208], stage1_26[209]},
      {stage1_27[53]},
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage2_30[35],stage2_29[38],stage2_28[43],stage2_27[74],stage2_26[97]}
   );
   gpc615_5 gpc2753 (
      {stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213], stage1_26[214]},
      {stage1_27[54]},
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage2_30[36],stage2_29[39],stage2_28[44],stage2_27[75],stage2_26[98]}
   );
   gpc615_5 gpc2754 (
      {stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage1_28[222]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[37],stage2_29[40],stage2_28[45],stage2_27[76]}
   );
   gpc615_5 gpc2755 (
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64]},
      {stage1_28[223]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[38],stage2_29[41],stage2_28[46],stage2_27[77]}
   );
   gpc615_5 gpc2756 (
      {stage1_27[65], stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69]},
      {stage1_28[224]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[39],stage2_29[42],stage2_28[47],stage2_27[78]}
   );
   gpc615_5 gpc2757 (
      {stage1_27[70], stage1_27[71], stage1_27[72], stage1_27[73], stage1_27[74]},
      {stage1_28[225]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[40],stage2_29[43],stage2_28[48],stage2_27[79]}
   );
   gpc615_5 gpc2758 (
      {stage1_27[75], stage1_27[76], stage1_27[77], stage1_27[78], stage1_27[79]},
      {stage1_28[226]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[41],stage2_29[44],stage2_28[49],stage2_27[80]}
   );
   gpc615_5 gpc2759 (
      {stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83], stage1_27[84]},
      {stage1_28[227]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[42],stage2_29[45],stage2_28[50],stage2_27[81]}
   );
   gpc615_5 gpc2760 (
      {stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage1_28[228]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[43],stage2_29[46],stage2_28[51],stage2_27[82]}
   );
   gpc615_5 gpc2761 (
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94]},
      {stage1_28[229]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[44],stage2_29[47],stage2_28[52],stage2_27[83]}
   );
   gpc615_5 gpc2762 (
      {stage1_27[95], stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99]},
      {stage1_28[230]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[45],stage2_29[48],stage2_28[53],stage2_27[84]}
   );
   gpc615_5 gpc2763 (
      {stage1_27[100], stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104]},
      {stage1_28[231]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[46],stage2_29[49],stage2_28[54],stage2_27[85]}
   );
   gpc615_5 gpc2764 (
      {stage1_27[105], stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109]},
      {stage1_28[232]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[47],stage2_29[50],stage2_28[55],stage2_27[86]}
   );
   gpc615_5 gpc2765 (
      {stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114]},
      {stage1_28[233]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[48],stage2_29[51],stage2_28[56],stage2_27[87]}
   );
   gpc615_5 gpc2766 (
      {stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage1_28[234]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[49],stage2_29[52],stage2_28[57],stage2_27[88]}
   );
   gpc615_5 gpc2767 (
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124]},
      {stage1_28[235]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[50],stage2_29[53],stage2_28[58],stage2_27[89]}
   );
   gpc615_5 gpc2768 (
      {stage1_27[125], stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129]},
      {stage1_28[236]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[51],stage2_29[54],stage2_28[59],stage2_27[90]}
   );
   gpc615_5 gpc2769 (
      {stage1_27[130], stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134]},
      {stage1_28[237]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[52],stage2_29[55],stage2_28[60],stage2_27[91]}
   );
   gpc615_5 gpc2770 (
      {stage1_27[135], stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139]},
      {stage1_28[238]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[53],stage2_29[56],stage2_28[61],stage2_27[92]}
   );
   gpc615_5 gpc2771 (
      {stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144]},
      {stage1_28[239]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[54],stage2_29[57],stage2_28[62],stage2_27[93]}
   );
   gpc615_5 gpc2772 (
      {stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage1_28[240]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[55],stage2_29[58],stage2_28[63],stage2_27[94]}
   );
   gpc615_5 gpc2773 (
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154]},
      {stage1_28[241]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[56],stage2_29[59],stage2_28[64],stage2_27[95]}
   );
   gpc615_5 gpc2774 (
      {stage1_27[155], stage1_27[156], stage1_27[157], stage1_27[158], 1'b0},
      {stage1_28[242]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[57],stage2_29[60],stage2_28[65],stage2_27[96]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[0],stage2_31[21],stage2_30[58],stage2_29[61]}
   );
   gpc606_5 gpc2776 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[1],stage2_31[22],stage2_30[59],stage2_29[62]}
   );
   gpc606_5 gpc2777 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[2],stage2_31[23],stage2_30[60],stage2_29[63]}
   );
   gpc606_5 gpc2778 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[3],stage2_31[24],stage2_30[61],stage2_29[64]}
   );
   gpc606_5 gpc2779 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[4],stage2_31[25],stage2_30[62],stage2_29[65]}
   );
   gpc606_5 gpc2780 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[5],stage2_31[26],stage2_30[63],stage2_29[66]}
   );
   gpc606_5 gpc2781 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[6],stage2_31[27],stage2_30[64],stage2_29[67]}
   );
   gpc606_5 gpc2782 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[7],stage2_31[28],stage2_30[65],stage2_29[68]}
   );
   gpc606_5 gpc2783 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[8],stage2_31[29],stage2_30[66],stage2_29[69]}
   );
   gpc606_5 gpc2784 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[9],stage2_31[30],stage2_30[67],stage2_29[70]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[10],stage2_32[10],stage2_31[31],stage2_30[68]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[11],stage2_32[11],stage2_31[32],stage2_30[69]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[12],stage2_32[12],stage2_31[33],stage2_30[70]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[13],stage2_32[13],stage2_31[34],stage2_30[71]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[14],stage2_32[14],stage2_31[35],stage2_30[72]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[15],stage2_32[15],stage2_31[36],stage2_30[73]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[16],stage2_32[16],stage2_31[37],stage2_30[74]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[17],stage2_32[17],stage2_31[38],stage2_30[75]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[18],stage2_32[18],stage2_31[39],stage2_30[76]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[19],stage2_32[19],stage2_31[40],stage2_30[77]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[20],stage2_32[20],stage2_31[41],stage2_30[78]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[21],stage2_32[21],stage2_31[42],stage2_30[79]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[22],stage2_32[22],stage2_31[43],stage2_30[80]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[23],stage2_32[23],stage2_31[44],stage2_30[81]}
   );
   gpc606_5 gpc2799 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[24],stage2_32[24],stage2_31[45],stage2_30[82]}
   );
   gpc606_5 gpc2800 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[25],stage2_32[25],stage2_31[46],stage2_30[83]}
   );
   gpc606_5 gpc2801 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[26],stage2_32[26],stage2_31[47],stage2_30[84]}
   );
   gpc606_5 gpc2802 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[27],stage2_32[27],stage2_31[48],stage2_30[85]}
   );
   gpc606_5 gpc2803 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[28],stage2_32[28],stage2_31[49],stage2_30[86]}
   );
   gpc606_5 gpc2804 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[29],stage2_32[29],stage2_31[50],stage2_30[87]}
   );
   gpc606_5 gpc2805 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[30],stage2_32[30],stage2_31[51],stage2_30[88]}
   );
   gpc606_5 gpc2806 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[31],stage2_32[31],stage2_31[52],stage2_30[89]}
   );
   gpc606_5 gpc2807 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[22],stage2_33[32],stage2_32[32],stage2_31[53]}
   );
   gpc606_5 gpc2808 (
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[23],stage2_33[33],stage2_32[33],stage2_31[54]}
   );
   gpc606_5 gpc2809 (
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[24],stage2_33[34],stage2_32[34],stage2_31[55]}
   );
   gpc606_5 gpc2810 (
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[25],stage2_33[35],stage2_32[35],stage2_31[56]}
   );
   gpc606_5 gpc2811 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[26],stage2_33[36],stage2_32[36],stage2_31[57]}
   );
   gpc606_5 gpc2812 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[27],stage2_33[37],stage2_32[37],stage2_31[58]}
   );
   gpc606_5 gpc2813 (
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[28],stage2_33[38],stage2_32[38],stage2_31[59]}
   );
   gpc606_5 gpc2814 (
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[29],stage2_33[39],stage2_32[39],stage2_31[60]}
   );
   gpc606_5 gpc2815 (
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[30],stage2_33[40],stage2_32[40],stage2_31[61]}
   );
   gpc606_5 gpc2816 (
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[31],stage2_33[41],stage2_32[41],stage2_31[62]}
   );
   gpc606_5 gpc2817 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[32],stage2_33[42],stage2_32[42],stage2_31[63]}
   );
   gpc606_5 gpc2818 (
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[33],stage2_33[43],stage2_32[43],stage2_31[64]}
   );
   gpc606_5 gpc2819 (
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[34],stage2_33[44],stage2_32[44],stage2_31[65]}
   );
   gpc606_5 gpc2820 (
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage1_33[78], stage1_33[79], stage1_33[80], 1'b0, 1'b0, 1'b0},
      {stage2_35[13],stage2_34[35],stage2_33[45],stage2_32[45],stage2_31[66]}
   );
   gpc1_1 gpc2821 (
      {stage1_1[62]},
      {stage2_1[31]}
   );
   gpc1_1 gpc2822 (
      {stage1_1[63]},
      {stage2_1[32]}
   );
   gpc1_1 gpc2823 (
      {stage1_1[64]},
      {stage2_1[33]}
   );
   gpc1_1 gpc2824 (
      {stage1_1[65]},
      {stage2_1[34]}
   );
   gpc1_1 gpc2825 (
      {stage1_1[66]},
      {stage2_1[35]}
   );
   gpc1_1 gpc2826 (
      {stage1_1[67]},
      {stage2_1[36]}
   );
   gpc1_1 gpc2827 (
      {stage1_1[68]},
      {stage2_1[37]}
   );
   gpc1_1 gpc2828 (
      {stage1_1[69]},
      {stage2_1[38]}
   );
   gpc1_1 gpc2829 (
      {stage1_1[70]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2830 (
      {stage1_1[71]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2831 (
      {stage1_1[72]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2832 (
      {stage1_1[73]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2833 (
      {stage1_1[74]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2834 (
      {stage1_1[75]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2835 (
      {stage1_1[76]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2836 (
      {stage1_1[77]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2837 (
      {stage1_1[78]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2838 (
      {stage1_1[79]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2839 (
      {stage1_1[80]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2840 (
      {stage1_1[81]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2841 (
      {stage1_1[82]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2842 (
      {stage1_1[83]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2843 (
      {stage1_1[84]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2844 (
      {stage1_1[85]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2845 (
      {stage1_1[86]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2846 (
      {stage1_1[87]},
      {stage2_1[56]}
   );
   gpc1_1 gpc2847 (
      {stage1_1[88]},
      {stage2_1[57]}
   );
   gpc1_1 gpc2848 (
      {stage1_1[89]},
      {stage2_1[58]}
   );
   gpc1_1 gpc2849 (
      {stage1_1[90]},
      {stage2_1[59]}
   );
   gpc1_1 gpc2850 (
      {stage1_1[91]},
      {stage2_1[60]}
   );
   gpc1_1 gpc2851 (
      {stage1_1[92]},
      {stage2_1[61]}
   );
   gpc1_1 gpc2852 (
      {stage1_1[93]},
      {stage2_1[62]}
   );
   gpc1_1 gpc2853 (
      {stage1_1[94]},
      {stage2_1[63]}
   );
   gpc1_1 gpc2854 (
      {stage1_1[95]},
      {stage2_1[64]}
   );
   gpc1_1 gpc2855 (
      {stage1_1[96]},
      {stage2_1[65]}
   );
   gpc1_1 gpc2856 (
      {stage1_1[97]},
      {stage2_1[66]}
   );
   gpc1_1 gpc2857 (
      {stage1_1[98]},
      {stage2_1[67]}
   );
   gpc1_1 gpc2858 (
      {stage1_1[99]},
      {stage2_1[68]}
   );
   gpc1_1 gpc2859 (
      {stage1_1[100]},
      {stage2_1[69]}
   );
   gpc1_1 gpc2860 (
      {stage1_1[101]},
      {stage2_1[70]}
   );
   gpc1_1 gpc2861 (
      {stage1_1[102]},
      {stage2_1[71]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[103]},
      {stage2_1[72]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[104]},
      {stage2_1[73]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[105]},
      {stage2_1[74]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[106]},
      {stage2_1[75]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[107]},
      {stage2_1[76]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[108]},
      {stage2_1[77]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[109]},
      {stage2_1[78]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[110]},
      {stage2_1[79]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[111]},
      {stage2_1[80]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[112]},
      {stage2_1[81]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[113]},
      {stage2_1[82]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[114]},
      {stage2_1[83]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[115]},
      {stage2_1[84]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[116]},
      {stage2_1[85]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[117]},
      {stage2_1[86]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[118]},
      {stage2_1[87]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[119]},
      {stage2_1[88]}
   );
   gpc1_1 gpc2879 (
      {stage1_1[120]},
      {stage2_1[89]}
   );
   gpc1_1 gpc2880 (
      {stage1_1[121]},
      {stage2_1[90]}
   );
   gpc1_1 gpc2881 (
      {stage1_1[122]},
      {stage2_1[91]}
   );
   gpc1_1 gpc2882 (
      {stage1_1[123]},
      {stage2_1[92]}
   );
   gpc1_1 gpc2883 (
      {stage1_1[124]},
      {stage2_1[93]}
   );
   gpc1_1 gpc2884 (
      {stage1_1[125]},
      {stage2_1[94]}
   );
   gpc1_1 gpc2885 (
      {stage1_1[126]},
      {stage2_1[95]}
   );
   gpc1_1 gpc2886 (
      {stage1_1[127]},
      {stage2_1[96]}
   );
   gpc1_1 gpc2887 (
      {stage1_1[128]},
      {stage2_1[97]}
   );
   gpc1_1 gpc2888 (
      {stage1_1[129]},
      {stage2_1[98]}
   );
   gpc1_1 gpc2889 (
      {stage1_1[130]},
      {stage2_1[99]}
   );
   gpc1_1 gpc2890 (
      {stage1_1[131]},
      {stage2_1[100]}
   );
   gpc1_1 gpc2891 (
      {stage1_1[132]},
      {stage2_1[101]}
   );
   gpc1_1 gpc2892 (
      {stage1_1[133]},
      {stage2_1[102]}
   );
   gpc1_1 gpc2893 (
      {stage1_1[134]},
      {stage2_1[103]}
   );
   gpc1_1 gpc2894 (
      {stage1_1[135]},
      {stage2_1[104]}
   );
   gpc1_1 gpc2895 (
      {stage1_1[136]},
      {stage2_1[105]}
   );
   gpc1_1 gpc2896 (
      {stage1_1[137]},
      {stage2_1[106]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[225]},
      {stage2_2[48]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[226]},
      {stage2_2[49]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[227]},
      {stage2_2[50]}
   );
   gpc1_1 gpc2900 (
      {stage1_3[169]},
      {stage2_3[69]}
   );
   gpc1_1 gpc2901 (
      {stage1_3[170]},
      {stage2_3[70]}
   );
   gpc1_1 gpc2902 (
      {stage1_3[171]},
      {stage2_3[71]}
   );
   gpc1_1 gpc2903 (
      {stage1_3[172]},
      {stage2_3[72]}
   );
   gpc1_1 gpc2904 (
      {stage1_3[173]},
      {stage2_3[73]}
   );
   gpc1_1 gpc2905 (
      {stage1_3[174]},
      {stage2_3[74]}
   );
   gpc1_1 gpc2906 (
      {stage1_3[175]},
      {stage2_3[75]}
   );
   gpc1_1 gpc2907 (
      {stage1_3[176]},
      {stage2_3[76]}
   );
   gpc1_1 gpc2908 (
      {stage1_3[177]},
      {stage2_3[77]}
   );
   gpc1_1 gpc2909 (
      {stage1_3[178]},
      {stage2_3[78]}
   );
   gpc1_1 gpc2910 (
      {stage1_3[179]},
      {stage2_3[79]}
   );
   gpc1_1 gpc2911 (
      {stage1_3[180]},
      {stage2_3[80]}
   );
   gpc1_1 gpc2912 (
      {stage1_3[181]},
      {stage2_3[81]}
   );
   gpc1_1 gpc2913 (
      {stage1_3[182]},
      {stage2_3[82]}
   );
   gpc1_1 gpc2914 (
      {stage1_3[183]},
      {stage2_3[83]}
   );
   gpc1_1 gpc2915 (
      {stage1_3[184]},
      {stage2_3[84]}
   );
   gpc1_1 gpc2916 (
      {stage1_3[185]},
      {stage2_3[85]}
   );
   gpc1_1 gpc2917 (
      {stage1_3[186]},
      {stage2_3[86]}
   );
   gpc1_1 gpc2918 (
      {stage1_3[187]},
      {stage2_3[87]}
   );
   gpc1_1 gpc2919 (
      {stage1_5[213]},
      {stage2_5[79]}
   );
   gpc1_1 gpc2920 (
      {stage1_5[214]},
      {stage2_5[80]}
   );
   gpc1_1 gpc2921 (
      {stage1_5[215]},
      {stage2_5[81]}
   );
   gpc1_1 gpc2922 (
      {stage1_5[216]},
      {stage2_5[82]}
   );
   gpc1_1 gpc2923 (
      {stage1_5[217]},
      {stage2_5[83]}
   );
   gpc1_1 gpc2924 (
      {stage1_7[218]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2925 (
      {stage1_7[219]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2926 (
      {stage1_7[220]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2927 (
      {stage1_7[221]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2928 (
      {stage1_7[222]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2929 (
      {stage1_7[223]},
      {stage2_7[109]}
   );
   gpc1_1 gpc2930 (
      {stage1_8[183]},
      {stage2_8[85]}
   );
   gpc1_1 gpc2931 (
      {stage1_8[184]},
      {stage2_8[86]}
   );
   gpc1_1 gpc2932 (
      {stage1_8[185]},
      {stage2_8[87]}
   );
   gpc1_1 gpc2933 (
      {stage1_8[186]},
      {stage2_8[88]}
   );
   gpc1_1 gpc2934 (
      {stage1_8[187]},
      {stage2_8[89]}
   );
   gpc1_1 gpc2935 (
      {stage1_8[188]},
      {stage2_8[90]}
   );
   gpc1_1 gpc2936 (
      {stage1_8[189]},
      {stage2_8[91]}
   );
   gpc1_1 gpc2937 (
      {stage1_8[190]},
      {stage2_8[92]}
   );
   gpc1_1 gpc2938 (
      {stage1_8[191]},
      {stage2_8[93]}
   );
   gpc1_1 gpc2939 (
      {stage1_8[192]},
      {stage2_8[94]}
   );
   gpc1_1 gpc2940 (
      {stage1_8[193]},
      {stage2_8[95]}
   );
   gpc1_1 gpc2941 (
      {stage1_8[194]},
      {stage2_8[96]}
   );
   gpc1_1 gpc2942 (
      {stage1_8[195]},
      {stage2_8[97]}
   );
   gpc1_1 gpc2943 (
      {stage1_8[196]},
      {stage2_8[98]}
   );
   gpc1_1 gpc2944 (
      {stage1_8[197]},
      {stage2_8[99]}
   );
   gpc1_1 gpc2945 (
      {stage1_8[198]},
      {stage2_8[100]}
   );
   gpc1_1 gpc2946 (
      {stage1_8[199]},
      {stage2_8[101]}
   );
   gpc1_1 gpc2947 (
      {stage1_8[200]},
      {stage2_8[102]}
   );
   gpc1_1 gpc2948 (
      {stage1_8[201]},
      {stage2_8[103]}
   );
   gpc1_1 gpc2949 (
      {stage1_8[202]},
      {stage2_8[104]}
   );
   gpc1_1 gpc2950 (
      {stage1_8[203]},
      {stage2_8[105]}
   );
   gpc1_1 gpc2951 (
      {stage1_8[204]},
      {stage2_8[106]}
   );
   gpc1_1 gpc2952 (
      {stage1_8[205]},
      {stage2_8[107]}
   );
   gpc1_1 gpc2953 (
      {stage1_9[211]},
      {stage2_9[72]}
   );
   gpc1_1 gpc2954 (
      {stage1_9[212]},
      {stage2_9[73]}
   );
   gpc1_1 gpc2955 (
      {stage1_9[213]},
      {stage2_9[74]}
   );
   gpc1_1 gpc2956 (
      {stage1_10[186]},
      {stage2_10[87]}
   );
   gpc1_1 gpc2957 (
      {stage1_10[187]},
      {stage2_10[88]}
   );
   gpc1_1 gpc2958 (
      {stage1_12[277]},
      {stage2_12[98]}
   );
   gpc1_1 gpc2959 (
      {stage1_12[278]},
      {stage2_12[99]}
   );
   gpc1_1 gpc2960 (
      {stage1_12[279]},
      {stage2_12[100]}
   );
   gpc1_1 gpc2961 (
      {stage1_12[280]},
      {stage2_12[101]}
   );
   gpc1_1 gpc2962 (
      {stage1_12[281]},
      {stage2_12[102]}
   );
   gpc1_1 gpc2963 (
      {stage1_14[238]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2964 (
      {stage1_14[239]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2965 (
      {stage1_14[240]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2966 (
      {stage1_14[241]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2967 (
      {stage1_14[242]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2968 (
      {stage1_14[243]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2969 (
      {stage1_14[244]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2970 (
      {stage1_14[245]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2971 (
      {stage1_14[246]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2972 (
      {stage1_14[247]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2973 (
      {stage1_14[248]},
      {stage2_14[90]}
   );
   gpc1_1 gpc2974 (
      {stage1_14[249]},
      {stage2_14[91]}
   );
   gpc1_1 gpc2975 (
      {stage1_14[250]},
      {stage2_14[92]}
   );
   gpc1_1 gpc2976 (
      {stage1_14[251]},
      {stage2_14[93]}
   );
   gpc1_1 gpc2977 (
      {stage1_14[252]},
      {stage2_14[94]}
   );
   gpc1_1 gpc2978 (
      {stage1_14[253]},
      {stage2_14[95]}
   );
   gpc1_1 gpc2979 (
      {stage1_14[254]},
      {stage2_14[96]}
   );
   gpc1_1 gpc2980 (
      {stage1_14[255]},
      {stage2_14[97]}
   );
   gpc1_1 gpc2981 (
      {stage1_14[256]},
      {stage2_14[98]}
   );
   gpc1_1 gpc2982 (
      {stage1_14[257]},
      {stage2_14[99]}
   );
   gpc1_1 gpc2983 (
      {stage1_14[258]},
      {stage2_14[100]}
   );
   gpc1_1 gpc2984 (
      {stage1_14[259]},
      {stage2_14[101]}
   );
   gpc1_1 gpc2985 (
      {stage1_14[260]},
      {stage2_14[102]}
   );
   gpc1_1 gpc2986 (
      {stage1_14[261]},
      {stage2_14[103]}
   );
   gpc1_1 gpc2987 (
      {stage1_14[262]},
      {stage2_14[104]}
   );
   gpc1_1 gpc2988 (
      {stage1_14[263]},
      {stage2_14[105]}
   );
   gpc1_1 gpc2989 (
      {stage1_14[264]},
      {stage2_14[106]}
   );
   gpc1_1 gpc2990 (
      {stage1_14[265]},
      {stage2_14[107]}
   );
   gpc1_1 gpc2991 (
      {stage1_14[266]},
      {stage2_14[108]}
   );
   gpc1_1 gpc2992 (
      {stage1_14[267]},
      {stage2_14[109]}
   );
   gpc1_1 gpc2993 (
      {stage1_14[268]},
      {stage2_14[110]}
   );
   gpc1_1 gpc2994 (
      {stage1_14[269]},
      {stage2_14[111]}
   );
   gpc1_1 gpc2995 (
      {stage1_14[270]},
      {stage2_14[112]}
   );
   gpc1_1 gpc2996 (
      {stage1_14[271]},
      {stage2_14[113]}
   );
   gpc1_1 gpc2997 (
      {stage1_14[272]},
      {stage2_14[114]}
   );
   gpc1_1 gpc2998 (
      {stage1_14[273]},
      {stage2_14[115]}
   );
   gpc1_1 gpc2999 (
      {stage1_14[274]},
      {stage2_14[116]}
   );
   gpc1_1 gpc3000 (
      {stage1_14[275]},
      {stage2_14[117]}
   );
   gpc1_1 gpc3001 (
      {stage1_14[276]},
      {stage2_14[118]}
   );
   gpc1_1 gpc3002 (
      {stage1_14[277]},
      {stage2_14[119]}
   );
   gpc1_1 gpc3003 (
      {stage1_14[278]},
      {stage2_14[120]}
   );
   gpc1_1 gpc3004 (
      {stage1_14[279]},
      {stage2_14[121]}
   );
   gpc1_1 gpc3005 (
      {stage1_14[280]},
      {stage2_14[122]}
   );
   gpc1_1 gpc3006 (
      {stage1_14[281]},
      {stage2_14[123]}
   );
   gpc1_1 gpc3007 (
      {stage1_14[282]},
      {stage2_14[124]}
   );
   gpc1_1 gpc3008 (
      {stage1_14[283]},
      {stage2_14[125]}
   );
   gpc1_1 gpc3009 (
      {stage1_14[284]},
      {stage2_14[126]}
   );
   gpc1_1 gpc3010 (
      {stage1_14[285]},
      {stage2_14[127]}
   );
   gpc1_1 gpc3011 (
      {stage1_14[286]},
      {stage2_14[128]}
   );
   gpc1_1 gpc3012 (
      {stage1_14[287]},
      {stage2_14[129]}
   );
   gpc1_1 gpc3013 (
      {stage1_14[288]},
      {stage2_14[130]}
   );
   gpc1_1 gpc3014 (
      {stage1_14[289]},
      {stage2_14[131]}
   );
   gpc1_1 gpc3015 (
      {stage1_14[290]},
      {stage2_14[132]}
   );
   gpc1_1 gpc3016 (
      {stage1_14[291]},
      {stage2_14[133]}
   );
   gpc1_1 gpc3017 (
      {stage1_14[292]},
      {stage2_14[134]}
   );
   gpc1_1 gpc3018 (
      {stage1_14[293]},
      {stage2_14[135]}
   );
   gpc1_1 gpc3019 (
      {stage1_14[294]},
      {stage2_14[136]}
   );
   gpc1_1 gpc3020 (
      {stage1_14[295]},
      {stage2_14[137]}
   );
   gpc1_1 gpc3021 (
      {stage1_14[296]},
      {stage2_14[138]}
   );
   gpc1_1 gpc3022 (
      {stage1_15[128]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3023 (
      {stage1_15[129]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3024 (
      {stage1_15[130]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3025 (
      {stage1_15[131]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3026 (
      {stage1_15[132]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3027 (
      {stage1_15[133]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3028 (
      {stage1_15[134]},
      {stage2_15[98]}
   );
   gpc1_1 gpc3029 (
      {stage1_15[135]},
      {stage2_15[99]}
   );
   gpc1_1 gpc3030 (
      {stage1_15[136]},
      {stage2_15[100]}
   );
   gpc1_1 gpc3031 (
      {stage1_15[137]},
      {stage2_15[101]}
   );
   gpc1_1 gpc3032 (
      {stage1_15[138]},
      {stage2_15[102]}
   );
   gpc1_1 gpc3033 (
      {stage1_15[139]},
      {stage2_15[103]}
   );
   gpc1_1 gpc3034 (
      {stage1_15[140]},
      {stage2_15[104]}
   );
   gpc1_1 gpc3035 (
      {stage1_15[141]},
      {stage2_15[105]}
   );
   gpc1_1 gpc3036 (
      {stage1_15[142]},
      {stage2_15[106]}
   );
   gpc1_1 gpc3037 (
      {stage1_15[143]},
      {stage2_15[107]}
   );
   gpc1_1 gpc3038 (
      {stage1_15[144]},
      {stage2_15[108]}
   );
   gpc1_1 gpc3039 (
      {stage1_15[145]},
      {stage2_15[109]}
   );
   gpc1_1 gpc3040 (
      {stage1_15[146]},
      {stage2_15[110]}
   );
   gpc1_1 gpc3041 (
      {stage1_15[147]},
      {stage2_15[111]}
   );
   gpc1_1 gpc3042 (
      {stage1_15[148]},
      {stage2_15[112]}
   );
   gpc1_1 gpc3043 (
      {stage1_15[149]},
      {stage2_15[113]}
   );
   gpc1_1 gpc3044 (
      {stage1_15[150]},
      {stage2_15[114]}
   );
   gpc1_1 gpc3045 (
      {stage1_15[151]},
      {stage2_15[115]}
   );
   gpc1_1 gpc3046 (
      {stage1_15[152]},
      {stage2_15[116]}
   );
   gpc1_1 gpc3047 (
      {stage1_15[153]},
      {stage2_15[117]}
   );
   gpc1_1 gpc3048 (
      {stage1_15[154]},
      {stage2_15[118]}
   );
   gpc1_1 gpc3049 (
      {stage1_15[155]},
      {stage2_15[119]}
   );
   gpc1_1 gpc3050 (
      {stage1_15[156]},
      {stage2_15[120]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[157]},
      {stage2_15[121]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[158]},
      {stage2_15[122]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[159]},
      {stage2_15[123]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[160]},
      {stage2_15[124]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[161]},
      {stage2_15[125]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[162]},
      {stage2_15[126]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[163]},
      {stage2_15[127]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[164]},
      {stage2_15[128]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[165]},
      {stage2_15[129]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[166]},
      {stage2_15[130]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[167]},
      {stage2_15[131]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[168]},
      {stage2_15[132]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[169]},
      {stage2_15[133]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[170]},
      {stage2_15[134]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[171]},
      {stage2_15[135]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[257]},
      {stage2_16[96]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[258]},
      {stage2_16[97]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[259]},
      {stage2_16[98]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[260]},
      {stage2_16[99]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[261]},
      {stage2_16[100]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[262]},
      {stage2_16[101]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[263]},
      {stage2_16[102]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[264]},
      {stage2_16[103]}
   );
   gpc1_1 gpc3074 (
      {stage1_17[234]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3075 (
      {stage1_17[235]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3076 (
      {stage1_17[236]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3077 (
      {stage1_17[237]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3078 (
      {stage1_17[238]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3079 (
      {stage1_17[239]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3080 (
      {stage1_17[240]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3081 (
      {stage1_17[241]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3082 (
      {stage1_17[242]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3083 (
      {stage1_17[243]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[244]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[245]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[246]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[247]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[248]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[249]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[250]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[251]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[252]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[253]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[254]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[255]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[256]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[257]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[258]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[259]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[260]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[261]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[262]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[263]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[264]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[265]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[266]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[267]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[268]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[269]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[270]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3111 (
      {stage1_18[198]},
      {stage2_18[79]}
   );
   gpc1_1 gpc3112 (
      {stage1_18[199]},
      {stage2_18[80]}
   );
   gpc1_1 gpc3113 (
      {stage1_18[200]},
      {stage2_18[81]}
   );
   gpc1_1 gpc3114 (
      {stage1_19[295]},
      {stage2_19[105]}
   );
   gpc1_1 gpc3115 (
      {stage1_19[296]},
      {stage2_19[106]}
   );
   gpc1_1 gpc3116 (
      {stage1_19[297]},
      {stage2_19[107]}
   );
   gpc1_1 gpc3117 (
      {stage1_19[298]},
      {stage2_19[108]}
   );
   gpc1_1 gpc3118 (
      {stage1_19[299]},
      {stage2_19[109]}
   );
   gpc1_1 gpc3119 (
      {stage1_20[172]},
      {stage2_20[111]}
   );
   gpc1_1 gpc3120 (
      {stage1_20[173]},
      {stage2_20[112]}
   );
   gpc1_1 gpc3121 (
      {stage1_20[174]},
      {stage2_20[113]}
   );
   gpc1_1 gpc3122 (
      {stage1_20[175]},
      {stage2_20[114]}
   );
   gpc1_1 gpc3123 (
      {stage1_20[176]},
      {stage2_20[115]}
   );
   gpc1_1 gpc3124 (
      {stage1_20[177]},
      {stage2_20[116]}
   );
   gpc1_1 gpc3125 (
      {stage1_20[178]},
      {stage2_20[117]}
   );
   gpc1_1 gpc3126 (
      {stage1_20[179]},
      {stage2_20[118]}
   );
   gpc1_1 gpc3127 (
      {stage1_20[180]},
      {stage2_20[119]}
   );
   gpc1_1 gpc3128 (
      {stage1_20[181]},
      {stage2_20[120]}
   );
   gpc1_1 gpc3129 (
      {stage1_20[182]},
      {stage2_20[121]}
   );
   gpc1_1 gpc3130 (
      {stage1_20[183]},
      {stage2_20[122]}
   );
   gpc1_1 gpc3131 (
      {stage1_20[184]},
      {stage2_20[123]}
   );
   gpc1_1 gpc3132 (
      {stage1_20[185]},
      {stage2_20[124]}
   );
   gpc1_1 gpc3133 (
      {stage1_20[186]},
      {stage2_20[125]}
   );
   gpc1_1 gpc3134 (
      {stage1_20[187]},
      {stage2_20[126]}
   );
   gpc1_1 gpc3135 (
      {stage1_20[188]},
      {stage2_20[127]}
   );
   gpc1_1 gpc3136 (
      {stage1_21[198]},
      {stage2_21[78]}
   );
   gpc1_1 gpc3137 (
      {stage1_24[194]},
      {stage2_24[82]}
   );
   gpc1_1 gpc3138 (
      {stage1_24[195]},
      {stage2_24[83]}
   );
   gpc1_1 gpc3139 (
      {stage1_24[196]},
      {stage2_24[84]}
   );
   gpc1_1 gpc3140 (
      {stage1_24[197]},
      {stage2_24[85]}
   );
   gpc1_1 gpc3141 (
      {stage1_24[198]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3142 (
      {stage1_24[199]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3143 (
      {stage1_24[200]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3144 (
      {stage1_24[201]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3145 (
      {stage1_24[202]},
      {stage2_24[90]}
   );
   gpc1_1 gpc3146 (
      {stage1_24[203]},
      {stage2_24[91]}
   );
   gpc1_1 gpc3147 (
      {stage1_24[204]},
      {stage2_24[92]}
   );
   gpc1_1 gpc3148 (
      {stage1_24[205]},
      {stage2_24[93]}
   );
   gpc1_1 gpc3149 (
      {stage1_24[206]},
      {stage2_24[94]}
   );
   gpc1_1 gpc3150 (
      {stage1_24[207]},
      {stage2_24[95]}
   );
   gpc1_1 gpc3151 (
      {stage1_24[208]},
      {stage2_24[96]}
   );
   gpc1_1 gpc3152 (
      {stage1_24[209]},
      {stage2_24[97]}
   );
   gpc1_1 gpc3153 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc3154 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc3155 (
      {stage1_25[209]},
      {stage2_25[62]}
   );
   gpc1_1 gpc3156 (
      {stage1_25[210]},
      {stage2_25[63]}
   );
   gpc1_1 gpc3157 (
      {stage1_25[211]},
      {stage2_25[64]}
   );
   gpc1_1 gpc3158 (
      {stage1_25[212]},
      {stage2_25[65]}
   );
   gpc1_1 gpc3159 (
      {stage1_25[213]},
      {stage2_25[66]}
   );
   gpc1_1 gpc3160 (
      {stage1_25[214]},
      {stage2_25[67]}
   );
   gpc1_1 gpc3161 (
      {stage1_25[215]},
      {stage2_25[68]}
   );
   gpc1_1 gpc3162 (
      {stage1_25[216]},
      {stage2_25[69]}
   );
   gpc1_1 gpc3163 (
      {stage1_25[217]},
      {stage2_25[70]}
   );
   gpc1_1 gpc3164 (
      {stage1_25[218]},
      {stage2_25[71]}
   );
   gpc1_1 gpc3165 (
      {stage1_25[219]},
      {stage2_25[72]}
   );
   gpc1_1 gpc3166 (
      {stage1_25[220]},
      {stage2_25[73]}
   );
   gpc1_1 gpc3167 (
      {stage1_25[221]},
      {stage2_25[74]}
   );
   gpc1_1 gpc3168 (
      {stage1_25[222]},
      {stage2_25[75]}
   );
   gpc1_1 gpc3169 (
      {stage1_25[223]},
      {stage2_25[76]}
   );
   gpc1_1 gpc3170 (
      {stage1_25[224]},
      {stage2_25[77]}
   );
   gpc1_1 gpc3171 (
      {stage1_25[225]},
      {stage2_25[78]}
   );
   gpc1_1 gpc3172 (
      {stage1_25[226]},
      {stage2_25[79]}
   );
   gpc1_1 gpc3173 (
      {stage1_25[227]},
      {stage2_25[80]}
   );
   gpc1_1 gpc3174 (
      {stage1_25[228]},
      {stage2_25[81]}
   );
   gpc1_1 gpc3175 (
      {stage1_25[229]},
      {stage2_25[82]}
   );
   gpc1_1 gpc3176 (
      {stage1_25[230]},
      {stage2_25[83]}
   );
   gpc1_1 gpc3177 (
      {stage1_25[231]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3178 (
      {stage1_25[232]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3179 (
      {stage1_25[233]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3180 (
      {stage1_25[234]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3181 (
      {stage1_28[243]},
      {stage2_28[66]}
   );
   gpc1_1 gpc3182 (
      {stage1_28[244]},
      {stage2_28[67]}
   );
   gpc1_1 gpc3183 (
      {stage1_28[245]},
      {stage2_28[68]}
   );
   gpc1_1 gpc3184 (
      {stage1_28[246]},
      {stage2_28[69]}
   );
   gpc1_1 gpc3185 (
      {stage1_28[247]},
      {stage2_28[70]}
   );
   gpc1_1 gpc3186 (
      {stage1_28[248]},
      {stage2_28[71]}
   );
   gpc1_1 gpc3187 (
      {stage1_28[249]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3188 (
      {stage1_28[250]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3189 (
      {stage1_28[251]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3190 (
      {stage1_29[186]},
      {stage2_29[71]}
   );
   gpc1_1 gpc3191 (
      {stage1_29[187]},
      {stage2_29[72]}
   );
   gpc1_1 gpc3192 (
      {stage1_29[188]},
      {stage2_29[73]}
   );
   gpc1_1 gpc3193 (
      {stage1_29[189]},
      {stage2_29[74]}
   );
   gpc1_1 gpc3194 (
      {stage1_29[190]},
      {stage2_29[75]}
   );
   gpc1_1 gpc3195 (
      {stage1_29[191]},
      {stage2_29[76]}
   );
   gpc1_1 gpc3196 (
      {stage1_29[192]},
      {stage2_29[77]}
   );
   gpc1_1 gpc3197 (
      {stage1_29[193]},
      {stage2_29[78]}
   );
   gpc1_1 gpc3198 (
      {stage1_29[194]},
      {stage2_29[79]}
   );
   gpc1_1 gpc3199 (
      {stage1_29[195]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3200 (
      {stage1_29[196]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3201 (
      {stage1_29[197]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3202 (
      {stage1_29[198]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3203 (
      {stage1_29[199]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3204 (
      {stage1_29[200]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3205 (
      {stage1_29[201]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3206 (
      {stage1_29[202]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3207 (
      {stage1_29[203]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3208 (
      {stage1_29[204]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3209 (
      {stage1_29[205]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3210 (
      {stage1_29[206]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3211 (
      {stage1_29[207]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3212 (
      {stage1_29[208]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3213 (
      {stage1_29[209]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3214 (
      {stage1_29[210]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3215 (
      {stage1_29[211]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3216 (
      {stage1_29[212]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3217 (
      {stage1_29[213]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3218 (
      {stage1_29[214]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3219 (
      {stage1_29[215]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3220 (
      {stage1_29[216]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3221 (
      {stage1_29[217]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3222 (
      {stage1_29[218]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3223 (
      {stage1_29[219]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3224 (
      {stage1_29[220]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3225 (
      {stage1_29[221]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3226 (
      {stage1_29[222]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3227 (
      {stage1_29[223]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3228 (
      {stage1_29[224]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3229 (
      {stage1_29[225]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3230 (
      {stage1_29[226]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3231 (
      {stage1_29[227]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3232 (
      {stage1_29[228]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3233 (
      {stage1_29[229]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3234 (
      {stage1_29[230]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3235 (
      {stage1_29[231]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3236 (
      {stage1_29[232]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3237 (
      {stage1_29[233]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3238 (
      {stage1_29[234]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3239 (
      {stage1_29[235]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3240 (
      {stage1_30[132]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3241 (
      {stage1_30[133]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3242 (
      {stage1_30[134]},
      {stage2_30[92]}
   );
   gpc1_1 gpc3243 (
      {stage1_30[135]},
      {stage2_30[93]}
   );
   gpc1_1 gpc3244 (
      {stage1_30[136]},
      {stage2_30[94]}
   );
   gpc1_1 gpc3245 (
      {stage1_30[137]},
      {stage2_30[95]}
   );
   gpc1_1 gpc3246 (
      {stage1_30[138]},
      {stage2_30[96]}
   );
   gpc1_1 gpc3247 (
      {stage1_30[139]},
      {stage2_30[97]}
   );
   gpc1_1 gpc3248 (
      {stage1_30[140]},
      {stage2_30[98]}
   );
   gpc1_1 gpc3249 (
      {stage1_30[141]},
      {stage2_30[99]}
   );
   gpc1_1 gpc3250 (
      {stage1_30[142]},
      {stage2_30[100]}
   );
   gpc1_1 gpc3251 (
      {stage1_30[143]},
      {stage2_30[101]}
   );
   gpc1_1 gpc3252 (
      {stage1_30[144]},
      {stage2_30[102]}
   );
   gpc1_1 gpc3253 (
      {stage1_30[145]},
      {stage2_30[103]}
   );
   gpc1_1 gpc3254 (
      {stage1_30[146]},
      {stage2_30[104]}
   );
   gpc1_1 gpc3255 (
      {stage1_30[147]},
      {stage2_30[105]}
   );
   gpc1_1 gpc3256 (
      {stage1_30[148]},
      {stage2_30[106]}
   );
   gpc1_1 gpc3257 (
      {stage1_30[149]},
      {stage2_30[107]}
   );
   gpc1_1 gpc3258 (
      {stage1_30[150]},
      {stage2_30[108]}
   );
   gpc1_1 gpc3259 (
      {stage1_30[151]},
      {stage2_30[109]}
   );
   gpc1_1 gpc3260 (
      {stage1_30[152]},
      {stage2_30[110]}
   );
   gpc1_1 gpc3261 (
      {stage1_30[153]},
      {stage2_30[111]}
   );
   gpc1_1 gpc3262 (
      {stage1_30[154]},
      {stage2_30[112]}
   );
   gpc1_1 gpc3263 (
      {stage1_30[155]},
      {stage2_30[113]}
   );
   gpc1_1 gpc3264 (
      {stage1_30[156]},
      {stage2_30[114]}
   );
   gpc1_1 gpc3265 (
      {stage1_30[157]},
      {stage2_30[115]}
   );
   gpc1_1 gpc3266 (
      {stage1_30[158]},
      {stage2_30[116]}
   );
   gpc1_1 gpc3267 (
      {stage1_30[159]},
      {stage2_30[117]}
   );
   gpc1_1 gpc3268 (
      {stage1_30[160]},
      {stage2_30[118]}
   );
   gpc1_1 gpc3269 (
      {stage1_30[161]},
      {stage2_30[119]}
   );
   gpc1_1 gpc3270 (
      {stage1_30[162]},
      {stage2_30[120]}
   );
   gpc1_1 gpc3271 (
      {stage1_30[163]},
      {stage2_30[121]}
   );
   gpc1_1 gpc3272 (
      {stage1_30[164]},
      {stage2_30[122]}
   );
   gpc1_1 gpc3273 (
      {stage1_30[165]},
      {stage2_30[123]}
   );
   gpc1_1 gpc3274 (
      {stage1_30[166]},
      {stage2_30[124]}
   );
   gpc1_1 gpc3275 (
      {stage1_30[167]},
      {stage2_30[125]}
   );
   gpc1_1 gpc3276 (
      {stage1_30[168]},
      {stage2_30[126]}
   );
   gpc1_1 gpc3277 (
      {stage1_30[169]},
      {stage2_30[127]}
   );
   gpc1_1 gpc3278 (
      {stage1_30[170]},
      {stage2_30[128]}
   );
   gpc1_1 gpc3279 (
      {stage1_30[171]},
      {stage2_30[129]}
   );
   gpc1_1 gpc3280 (
      {stage1_31[144]},
      {stage2_31[67]}
   );
   gpc1_1 gpc3281 (
      {stage1_31[145]},
      {stage2_31[68]}
   );
   gpc1_1 gpc3282 (
      {stage1_31[146]},
      {stage2_31[69]}
   );
   gpc1_1 gpc3283 (
      {stage1_31[147]},
      {stage2_31[70]}
   );
   gpc1_1 gpc3284 (
      {stage1_31[148]},
      {stage2_31[71]}
   );
   gpc1_1 gpc3285 (
      {stage1_31[149]},
      {stage2_31[72]}
   );
   gpc1_1 gpc3286 (
      {stage1_31[150]},
      {stage2_31[73]}
   );
   gpc1_1 gpc3287 (
      {stage1_31[151]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3288 (
      {stage1_31[152]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3289 (
      {stage1_31[153]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3290 (
      {stage1_31[154]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3291 (
      {stage1_31[155]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3292 (
      {stage1_31[156]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3293 (
      {stage1_31[157]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3294 (
      {stage1_31[158]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3295 (
      {stage1_31[159]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3296 (
      {stage1_31[160]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3297 (
      {stage1_32[132]},
      {stage2_32[46]}
   );
   gpc1_1 gpc3298 (
      {stage1_32[133]},
      {stage2_32[47]}
   );
   gpc1_1 gpc3299 (
      {stage1_32[134]},
      {stage2_32[48]}
   );
   gpc1_1 gpc3300 (
      {stage1_32[135]},
      {stage2_32[49]}
   );
   gpc1_1 gpc3301 (
      {stage1_32[136]},
      {stage2_32[50]}
   );
   gpc1_1 gpc3302 (
      {stage1_32[137]},
      {stage2_32[51]}
   );
   gpc1_1 gpc3303 (
      {stage1_32[138]},
      {stage2_32[52]}
   );
   gpc1_1 gpc3304 (
      {stage1_32[139]},
      {stage2_32[53]}
   );
   gpc1_1 gpc3305 (
      {stage1_32[140]},
      {stage2_32[54]}
   );
   gpc1_1 gpc3306 (
      {stage1_32[141]},
      {stage2_32[55]}
   );
   gpc1_1 gpc3307 (
      {stage1_32[142]},
      {stage2_32[56]}
   );
   gpc1_1 gpc3308 (
      {stage1_32[143]},
      {stage2_32[57]}
   );
   gpc1_1 gpc3309 (
      {stage1_32[144]},
      {stage2_32[58]}
   );
   gpc1_1 gpc3310 (
      {stage1_32[145]},
      {stage2_32[59]}
   );
   gpc1_1 gpc3311 (
      {stage1_32[146]},
      {stage2_32[60]}
   );
   gpc1_1 gpc3312 (
      {stage1_32[147]},
      {stage2_32[61]}
   );
   gpc1_1 gpc3313 (
      {stage1_32[148]},
      {stage2_32[62]}
   );
   gpc1_1 gpc3314 (
      {stage1_32[149]},
      {stage2_32[63]}
   );
   gpc1_1 gpc3315 (
      {stage1_32[150]},
      {stage2_32[64]}
   );
   gpc1163_5 gpc3316 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc3317 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc3318 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc3319 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc1163_5 gpc3320 (
      {stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_2[4]},
      {stage2_3[4]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc1163_5 gpc3321 (
      {stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_2[5]},
      {stage2_3[5]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1163_5 gpc3322 (
      {stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[6]},
      {stage2_3[6]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3323 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[0],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc3324 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[1],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc3325 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[2],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc3326 (
      {stage2_1[60], stage2_1[61], stage2_1[62], stage2_1[63], stage2_1[64], stage2_1[65]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[3],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc3327 (
      {stage2_1[66], stage2_1[67], stage2_1[68], stage2_1[69], stage2_1[70], stage2_1[71]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[4],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3328 (
      {stage2_1[72], stage2_1[73], stage2_1[74], stage2_1[75], stage2_1[76], stage2_1[77]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[5],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3329 (
      {stage2_1[78], stage2_1[79], stage2_1[80], stage2_1[81], stage2_1[82], stage2_1[83]},
      {stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage3_5[6],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3330 (
      {stage2_1[84], stage2_1[85], stage2_1[86], stage2_1[87], stage2_1[88], stage2_1[89]},
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage3_5[7],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3331 (
      {stage2_1[90], stage2_1[91], stage2_1[92], stage2_1[93], stage2_1[94], stage2_1[95]},
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60]},
      {stage3_5[8],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3332 (
      {stage2_1[96], stage2_1[97], stage2_1[98], stage2_1[99], stage2_1[100], stage2_1[101]},
      {stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage3_5[9],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3333 (
      {stage2_1[102], stage2_1[103], stage2_1[104], stage2_1[105], stage2_1[106], 1'b0},
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage3_5[10],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc606_5 gpc3334 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[11],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc606_5 gpc3335 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[12],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc606_5 gpc3336 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[13],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc606_5 gpc3337 (
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[14],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc606_5 gpc3338 (
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[15],stage3_4[22],stage3_3[22],stage3_2[22]}
   );
   gpc606_5 gpc3339 (
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[16],stage3_4[23],stage3_3[23],stage3_2[23]}
   );
   gpc615_5 gpc3340 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[17],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3341 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[18],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3342 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[19],stage3_4[26],stage3_3[26]}
   );
   gpc606_5 gpc3343 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[20],stage3_4[27]}
   );
   gpc606_5 gpc3344 (
      {stage2_4[45], stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[21],stage3_4[28]}
   );
   gpc606_5 gpc3345 (
      {stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[22],stage3_4[29]}
   );
   gpc615_5 gpc3346 (
      {stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[12],stage3_5[23],stage3_4[30]}
   );
   gpc615_5 gpc3347 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[13],stage3_5[24],stage3_4[31]}
   );
   gpc615_5 gpc3348 (
      {stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[14],stage3_5[25],stage3_4[32]}
   );
   gpc615_5 gpc3349 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[15],stage3_5[26],stage3_4[33]}
   );
   gpc615_5 gpc3350 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[16],stage3_5[27],stage3_4[34]}
   );
   gpc606_5 gpc3351 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[17],stage3_5[28]}
   );
   gpc606_5 gpc3352 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[18],stage3_5[29]}
   );
   gpc606_5 gpc3353 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[19],stage3_5[30]}
   );
   gpc606_5 gpc3354 (
      {stage2_5[41], stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[11],stage3_7[14],stage3_6[20],stage3_5[31]}
   );
   gpc606_5 gpc3355 (
      {stage2_5[47], stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[12],stage3_7[15],stage3_6[21],stage3_5[32]}
   );
   gpc606_5 gpc3356 (
      {stage2_5[53], stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[13],stage3_7[16],stage3_6[22],stage3_5[33]}
   );
   gpc606_5 gpc3357 (
      {stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[14],stage3_7[17],stage3_6[23],stage3_5[34]}
   );
   gpc606_5 gpc3358 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[15],stage3_7[18],stage3_6[24],stage3_5[35]}
   );
   gpc615_5 gpc3359 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[48]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[8],stage3_8[16],stage3_7[19],stage3_6[25]}
   );
   gpc615_5 gpc3360 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[49]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[9],stage3_8[17],stage3_7[20],stage3_6[26]}
   );
   gpc615_5 gpc3361 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[50]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[10],stage3_8[18],stage3_7[21],stage3_6[27]}
   );
   gpc615_5 gpc3362 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[51]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[11],stage3_8[19],stage3_7[22],stage3_6[28]}
   );
   gpc615_5 gpc3363 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[52]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[12],stage3_8[20],stage3_7[23],stage3_6[29]}
   );
   gpc615_5 gpc3364 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[53]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[13],stage3_8[21],stage3_7[24],stage3_6[30]}
   );
   gpc615_5 gpc3365 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[54]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[14],stage3_8[22],stage3_7[25],stage3_6[31]}
   );
   gpc615_5 gpc3366 (
      {stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage2_8[42]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[7],stage3_9[15],stage3_8[23],stage3_7[26]}
   );
   gpc615_5 gpc3367 (
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64]},
      {stage2_8[43]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[8],stage3_9[16],stage3_8[24],stage3_7[27]}
   );
   gpc615_5 gpc3368 (
      {stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69]},
      {stage2_8[44]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[9],stage3_9[17],stage3_8[25],stage3_7[28]}
   );
   gpc1343_5 gpc3369 (
      {stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[3],stage3_10[10],stage3_9[18],stage3_8[26]}
   );
   gpc1343_5 gpc3370 (
      {stage2_8[48], stage2_8[49], stage2_8[50]},
      {stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25]},
      {stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_11[1]},
      {stage3_12[1],stage3_11[4],stage3_10[11],stage3_9[19],stage3_8[27]}
   );
   gpc1343_5 gpc3371 (
      {stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_10[6], stage2_10[7], stage2_10[8]},
      {stage2_11[2]},
      {stage3_12[2],stage3_11[5],stage3_10[12],stage3_9[20],stage3_8[28]}
   );
   gpc606_5 gpc3372 (
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13], stage2_10[14]},
      {stage3_12[3],stage3_11[6],stage3_10[13],stage3_9[21],stage3_8[29]}
   );
   gpc606_5 gpc3373 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage3_12[4],stage3_11[7],stage3_10[14],stage3_9[22],stage3_8[30]}
   );
   gpc606_5 gpc3374 (
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25], stage2_10[26]},
      {stage3_12[5],stage3_11[8],stage3_10[15],stage3_9[23],stage3_8[31]}
   );
   gpc606_5 gpc3375 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31], stage2_10[32]},
      {stage3_12[6],stage3_11[9],stage3_10[16],stage3_9[24],stage3_8[32]}
   );
   gpc606_5 gpc3376 (
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage3_12[7],stage3_11[10],stage3_10[17],stage3_9[25],stage3_8[33]}
   );
   gpc606_5 gpc3377 (
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage3_12[8],stage3_11[11],stage3_10[18],stage3_9[26],stage3_8[34]}
   );
   gpc606_5 gpc3378 (
      {stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94], stage2_8[95]},
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage3_12[9],stage3_11[12],stage3_10[19],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc3379 (
      {stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100], stage2_8[101]},
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage3_12[10],stage3_11[13],stage3_10[20],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc3380 (
      {stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106], stage2_8[107]},
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage3_12[11],stage3_11[14],stage3_10[21],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc3381 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage3_13[0],stage3_12[12],stage3_11[15],stage3_10[22],stage3_9[30]}
   );
   gpc615_5 gpc3382 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67]},
      {stage2_11[9]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[13],stage3_11[16],stage3_10[23]}
   );
   gpc615_5 gpc3383 (
      {stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72]},
      {stage2_11[10]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[14],stage3_11[17],stage3_10[24]}
   );
   gpc615_5 gpc3384 (
      {stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage2_11[11]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[15],stage3_11[18],stage3_10[25]}
   );
   gpc615_5 gpc3385 (
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82]},
      {stage2_11[12]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[16],stage3_11[19],stage3_10[26]}
   );
   gpc615_5 gpc3386 (
      {stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87]},
      {stage2_11[13]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[17],stage3_11[20],stage3_10[27]}
   );
   gpc606_5 gpc3387 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[5],stage3_13[6],stage3_12[18],stage3_11[21]}
   );
   gpc606_5 gpc3388 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[6],stage3_13[7],stage3_12[19],stage3_11[22]}
   );
   gpc606_5 gpc3389 (
      {stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[7],stage3_13[8],stage3_12[20],stage3_11[23]}
   );
   gpc606_5 gpc3390 (
      {stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[8],stage3_13[9],stage3_12[21],stage3_11[24]}
   );
   gpc606_5 gpc3391 (
      {stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[9],stage3_13[10],stage3_12[22],stage3_11[25]}
   );
   gpc606_5 gpc3392 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[10],stage3_13[11],stage3_12[23],stage3_11[26]}
   );
   gpc606_5 gpc3393 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[11],stage3_13[12],stage3_12[24],stage3_11[27]}
   );
   gpc606_5 gpc3394 (
      {stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[12],stage3_13[13],stage3_12[25],stage3_11[28]}
   );
   gpc606_5 gpc3395 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[13],stage3_13[14],stage3_12[26],stage3_11[29]}
   );
   gpc606_5 gpc3396 (
      {stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[14],stage3_13[15],stage3_12[27],stage3_11[30]}
   );
   gpc606_5 gpc3397 (
      {stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[15],stage3_13[16],stage3_12[28],stage3_11[31]}
   );
   gpc606_5 gpc3398 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[11],stage3_14[16],stage3_13[17],stage3_12[29]}
   );
   gpc606_5 gpc3399 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[12],stage3_14[17],stage3_13[18],stage3_12[30]}
   );
   gpc606_5 gpc3400 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[13],stage3_14[18],stage3_13[19],stage3_12[31]}
   );
   gpc606_5 gpc3401 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[14],stage3_14[19],stage3_13[20],stage3_12[32]}
   );
   gpc606_5 gpc3402 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[15],stage3_14[20],stage3_13[21],stage3_12[33]}
   );
   gpc606_5 gpc3403 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[16],stage3_14[21],stage3_13[22],stage3_12[34]}
   );
   gpc606_5 gpc3404 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[17],stage3_14[22],stage3_13[23],stage3_12[35]}
   );
   gpc606_5 gpc3405 (
      {stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[18],stage3_14[23],stage3_13[24],stage3_12[36]}
   );
   gpc606_5 gpc3406 (
      {stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[19],stage3_14[24],stage3_13[25],stage3_12[37]}
   );
   gpc606_5 gpc3407 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[20],stage3_14[25],stage3_13[26],stage3_12[38]}
   );
   gpc606_5 gpc3408 (
      {stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94], stage2_12[95]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[21],stage3_14[26],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc3409 (
      {stage2_12[96], stage2_12[97], stage2_12[98], stage2_12[99], stage2_12[100], stage2_12[101]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[22],stage3_14[27],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc3410 (
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[23],stage3_14[28],stage3_13[29]}
   );
   gpc606_5 gpc3411 (
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[24],stage3_14[29],stage3_13[30]}
   );
   gpc606_5 gpc3412 (
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[25],stage3_14[30],stage3_13[31]}
   );
   gpc606_5 gpc3413 (
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[26],stage3_14[31],stage3_13[32]}
   );
   gpc615_5 gpc3414 (
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94]},
      {stage2_14[72]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[27],stage3_14[32],stage3_13[33]}
   );
   gpc615_5 gpc3415 (
      {stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_15[30]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[5],stage3_16[17],stage3_15[28],stage3_14[33]}
   );
   gpc615_5 gpc3416 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[31]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[6],stage3_16[18],stage3_15[29],stage3_14[34]}
   );
   gpc615_5 gpc3417 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[32]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[7],stage3_16[19],stage3_15[30],stage3_14[35]}
   );
   gpc615_5 gpc3418 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[33]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[8],stage3_16[20],stage3_15[31],stage3_14[36]}
   );
   gpc615_5 gpc3419 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[34]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[9],stage3_16[21],stage3_15[32],stage3_14[37]}
   );
   gpc615_5 gpc3420 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], stage2_14[102]},
      {stage2_15[35]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[10],stage3_16[22],stage3_15[33],stage3_14[38]}
   );
   gpc615_5 gpc3421 (
      {stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_15[36]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[11],stage3_16[23],stage3_15[34],stage3_14[39]}
   );
   gpc615_5 gpc3422 (
      {stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111], stage2_14[112]},
      {stage2_15[37]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[12],stage3_16[24],stage3_15[35],stage3_14[40]}
   );
   gpc615_5 gpc3423 (
      {stage2_14[113], stage2_14[114], stage2_14[115], stage2_14[116], stage2_14[117]},
      {stage2_15[38]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[13],stage3_16[25],stage3_15[36],stage3_14[41]}
   );
   gpc615_5 gpc3424 (
      {stage2_14[118], stage2_14[119], stage2_14[120], stage2_14[121], stage2_14[122]},
      {stage2_15[39]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[14],stage3_16[26],stage3_15[37],stage3_14[42]}
   );
   gpc615_5 gpc3425 (
      {stage2_14[123], stage2_14[124], stage2_14[125], stage2_14[126], stage2_14[127]},
      {stage2_15[40]},
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage3_18[10],stage3_17[15],stage3_16[27],stage3_15[38],stage3_14[43]}
   );
   gpc615_5 gpc3426 (
      {stage2_14[128], stage2_14[129], stage2_14[130], stage2_14[131], stage2_14[132]},
      {stage2_15[41]},
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage3_18[11],stage3_17[16],stage3_16[28],stage3_15[39],stage3_14[44]}
   );
   gpc2135_5 gpc3427 (
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46]},
      {stage2_16[72], stage2_16[73], stage2_16[74]},
      {stage2_17[0]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[12],stage3_17[17],stage3_16[29],stage3_15[40]}
   );
   gpc606_5 gpc3428 (
      {stage2_15[47], stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[1],stage3_18[13],stage3_17[18],stage3_16[30],stage3_15[41]}
   );
   gpc606_5 gpc3429 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[2],stage3_18[14],stage3_17[19],stage3_16[31],stage3_15[42]}
   );
   gpc606_5 gpc3430 (
      {stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[3],stage3_18[15],stage3_17[20],stage3_16[32],stage3_15[43]}
   );
   gpc606_5 gpc3431 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69], stage2_15[70]},
      {stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24]},
      {stage3_19[4],stage3_18[16],stage3_17[21],stage3_16[33],stage3_15[44]}
   );
   gpc606_5 gpc3432 (
      {stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76]},
      {stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30]},
      {stage3_19[5],stage3_18[17],stage3_17[22],stage3_16[34],stage3_15[45]}
   );
   gpc606_5 gpc3433 (
      {stage2_15[77], stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36]},
      {stage3_19[6],stage3_18[18],stage3_17[23],stage3_16[35],stage3_15[46]}
   );
   gpc606_5 gpc3434 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87], stage2_15[88]},
      {stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42]},
      {stage3_19[7],stage3_18[19],stage3_17[24],stage3_16[36],stage3_15[47]}
   );
   gpc606_5 gpc3435 (
      {stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92], stage2_15[93], stage2_15[94]},
      {stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48]},
      {stage3_19[8],stage3_18[20],stage3_17[25],stage3_16[37],stage3_15[48]}
   );
   gpc606_5 gpc3436 (
      {stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80]},
      {stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6], stage2_18[7]},
      {stage3_20[0],stage3_19[9],stage3_18[21],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc3437 (
      {stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[10],stage3_18[22],stage3_17[27]}
   );
   gpc606_5 gpc3438 (
      {stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[11],stage3_18[23],stage3_17[28]}
   );
   gpc606_5 gpc3439 (
      {stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[12],stage3_18[24],stage3_17[29]}
   );
   gpc606_5 gpc3440 (
      {stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[13],stage3_18[25],stage3_17[30]}
   );
   gpc606_5 gpc3441 (
      {stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[5],stage3_19[14],stage3_18[26],stage3_17[31]}
   );
   gpc606_5 gpc3442 (
      {stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83], stage2_17[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage3_21[5],stage3_20[6],stage3_19[15],stage3_18[27],stage3_17[32]}
   );
   gpc606_5 gpc3443 (
      {stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89], stage2_17[90]},
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage3_21[6],stage3_20[7],stage3_19[16],stage3_18[28],stage3_17[33]}
   );
   gpc606_5 gpc3444 (
      {stage2_17[91], stage2_17[92], stage2_17[93], stage2_17[94], stage2_17[95], stage2_17[96]},
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage3_21[7],stage3_20[8],stage3_19[17],stage3_18[29],stage3_17[34]}
   );
   gpc606_5 gpc3445 (
      {stage2_17[97], stage2_17[98], stage2_17[99], stage2_17[100], stage2_17[101], stage2_17[102]},
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage3_21[8],stage3_20[9],stage3_19[18],stage3_18[30],stage3_17[35]}
   );
   gpc606_5 gpc3446 (
      {stage2_17[103], stage2_17[104], stage2_17[105], stage2_17[106], stage2_17[107], stage2_17[108]},
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage3_21[9],stage3_20[10],stage3_19[19],stage3_18[31],stage3_17[36]}
   );
   gpc1343_5 gpc3447 (
      {stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[10],stage3_20[11],stage3_19[20],stage3_18[32]}
   );
   gpc1343_5 gpc3448 (
      {stage2_18[11], stage2_18[12], stage2_18[13]},
      {stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[11],stage3_20[12],stage3_19[21],stage3_18[33]}
   );
   gpc1343_5 gpc3449 (
      {stage2_18[14], stage2_18[15], stage2_18[16]},
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71]},
      {stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_21[2]},
      {stage3_22[2],stage3_21[12],stage3_20[13],stage3_19[22],stage3_18[34]}
   );
   gpc1343_5 gpc3450 (
      {stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[72], stage2_19[73], stage2_19[74], stage2_19[75]},
      {stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage2_21[3]},
      {stage3_22[3],stage3_21[13],stage3_20[14],stage3_19[23],stage3_18[35]}
   );
   gpc615_5 gpc3451 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[76]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[4],stage3_21[14],stage3_20[15],stage3_19[24],stage3_18[36]}
   );
   gpc615_5 gpc3452 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[77]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[5],stage3_21[15],stage3_20[16],stage3_19[25],stage3_18[37]}
   );
   gpc615_5 gpc3453 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[78]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[6],stage3_21[16],stage3_20[17],stage3_19[26],stage3_18[38]}
   );
   gpc615_5 gpc3454 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[79]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[7],stage3_21[17],stage3_20[18],stage3_19[27],stage3_18[39]}
   );
   gpc615_5 gpc3455 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[80]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[8],stage3_21[18],stage3_20[19],stage3_19[28],stage3_18[40]}
   );
   gpc615_5 gpc3456 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[81]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[9],stage3_21[19],stage3_20[20],stage3_19[29],stage3_18[41]}
   );
   gpc615_5 gpc3457 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[82]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[10],stage3_21[20],stage3_20[21],stage3_19[30],stage3_18[42]}
   );
   gpc615_5 gpc3458 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[83]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[11],stage3_21[21],stage3_20[22],stage3_19[31],stage3_18[43]}
   );
   gpc615_5 gpc3459 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[84]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[12],stage3_21[22],stage3_20[23],stage3_19[32],stage3_18[44]}
   );
   gpc615_5 gpc3460 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[85]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[13],stage3_21[23],stage3_20[24],stage3_19[33],stage3_18[45]}
   );
   gpc615_5 gpc3461 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[86]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[14],stage3_21[24],stage3_20[25],stage3_19[34],stage3_18[46]}
   );
   gpc615_5 gpc3462 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[87]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[15],stage3_21[25],stage3_20[26],stage3_19[35],stage3_18[47]}
   );
   gpc615_5 gpc3463 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[84]},
      {stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage3_23[0],stage3_22[16],stage3_21[26],stage3_20[27],stage3_19[36]}
   );
   gpc615_5 gpc3464 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[85]},
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage3_23[1],stage3_22[17],stage3_21[27],stage3_20[28],stage3_19[37]}
   );
   gpc606_5 gpc3465 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[18],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3466 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[3],stage3_22[19],stage3_21[29],stage3_20[30]}
   );
   gpc606_5 gpc3467 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[4],stage3_22[20],stage3_21[30],stage3_20[31]}
   );
   gpc606_5 gpc3468 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[5],stage3_22[21],stage3_21[31],stage3_20[32]}
   );
   gpc606_5 gpc3469 (
      {stage2_20[110], stage2_20[111], stage2_20[112], stage2_20[113], stage2_20[114], stage2_20[115]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[6],stage3_22[22],stage3_21[32],stage3_20[33]}
   );
   gpc1163_5 gpc3470 (
      {stage2_21[16], stage2_21[17], stage2_21[18]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage2_23[0]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[5],stage3_23[7],stage3_22[23],stage3_21[33]}
   );
   gpc1163_5 gpc3471 (
      {stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[1]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[6],stage3_23[8],stage3_22[24],stage3_21[34]}
   );
   gpc1163_5 gpc3472 (
      {stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage2_23[2]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[7],stage3_23[9],stage3_22[25],stage3_21[35]}
   );
   gpc1163_5 gpc3473 (
      {stage2_21[25], stage2_21[26], stage2_21[27]},
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53]},
      {stage2_23[3]},
      {stage2_24[3]},
      {stage3_25[3],stage3_24[8],stage3_23[10],stage3_22[26],stage3_21[36]}
   );
   gpc1163_5 gpc3474 (
      {stage2_21[28], stage2_21[29], stage2_21[30]},
      {stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[4]},
      {stage2_24[4]},
      {stage3_25[4],stage3_24[9],stage3_23[11],stage3_22[27],stage3_21[37]}
   );
   gpc1163_5 gpc3475 (
      {stage2_21[31], stage2_21[32], stage2_21[33]},
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65]},
      {stage2_23[5]},
      {stage2_24[5]},
      {stage3_25[5],stage3_24[10],stage3_23[12],stage3_22[28],stage3_21[38]}
   );
   gpc606_5 gpc3476 (
      {stage2_21[34], stage2_21[35], stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[6],stage3_24[11],stage3_23[13],stage3_22[29],stage3_21[39]}
   );
   gpc606_5 gpc3477 (
      {stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[7],stage3_24[12],stage3_23[14],stage3_22[30],stage3_21[40]}
   );
   gpc606_5 gpc3478 (
      {stage2_21[46], stage2_21[47], stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[8],stage3_24[13],stage3_23[15],stage3_22[31],stage3_21[41]}
   );
   gpc606_5 gpc3479 (
      {stage2_21[52], stage2_21[53], stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[9],stage3_24[14],stage3_23[16],stage3_22[32],stage3_21[42]}
   );
   gpc606_5 gpc3480 (
      {stage2_21[58], stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[10],stage3_24[15],stage3_23[17],stage3_22[33],stage3_21[43]}
   );
   gpc615_5 gpc3481 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40]},
      {stage2_24[6]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[11],stage3_24[16],stage3_23[18]}
   );
   gpc615_5 gpc3482 (
      {stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45]},
      {stage2_24[7]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[1],stage3_25[12],stage3_24[17],stage3_23[19]}
   );
   gpc615_5 gpc3483 (
      {stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_24[8]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[2],stage3_25[13],stage3_24[18],stage3_23[20]}
   );
   gpc615_5 gpc3484 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55]},
      {stage2_24[9]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[3],stage3_25[14],stage3_24[19],stage3_23[21]}
   );
   gpc615_5 gpc3485 (
      {stage2_23[56], stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60]},
      {stage2_24[10]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[4],stage3_25[15],stage3_24[20],stage3_23[22]}
   );
   gpc615_5 gpc3486 (
      {stage2_23[61], stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65]},
      {stage2_24[11]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[5],stage3_25[16],stage3_24[21],stage3_23[23]}
   );
   gpc615_5 gpc3487 (
      {stage2_23[66], stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70]},
      {stage2_24[12]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[6],stage3_25[17],stage3_24[22],stage3_23[24]}
   );
   gpc615_5 gpc3488 (
      {stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75]},
      {stage2_24[13]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[7],stage3_25[18],stage3_24[23],stage3_23[25]}
   );
   gpc615_5 gpc3489 (
      {stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_24[14]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[8],stage3_25[19],stage3_24[24],stage3_23[26]}
   );
   gpc615_5 gpc3490 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85]},
      {stage2_24[15]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[9],stage3_25[20],stage3_24[25],stage3_23[27]}
   );
   gpc615_5 gpc3491 (
      {stage2_23[86], stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90]},
      {stage2_24[16]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[10],stage3_25[21],stage3_24[26],stage3_23[28]}
   );
   gpc606_5 gpc3492 (
      {stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[11],stage3_26[11],stage3_25[22],stage3_24[27]}
   );
   gpc606_5 gpc3493 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[12],stage3_26[12],stage3_25[23],stage3_24[28]}
   );
   gpc606_5 gpc3494 (
      {stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[13],stage3_26[13],stage3_25[24],stage3_24[29]}
   );
   gpc606_5 gpc3495 (
      {stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[14],stage3_26[14],stage3_25[25],stage3_24[30]}
   );
   gpc606_5 gpc3496 (
      {stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[15],stage3_26[15],stage3_25[26],stage3_24[31]}
   );
   gpc606_5 gpc3497 (
      {stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[16],stage3_26[16],stage3_25[27],stage3_24[32]}
   );
   gpc606_5 gpc3498 (
      {stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[17],stage3_26[17],stage3_25[28],stage3_24[33]}
   );
   gpc606_5 gpc3499 (
      {stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[18],stage3_26[18],stage3_25[29],stage3_24[34]}
   );
   gpc606_5 gpc3500 (
      {stage2_24[65], stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70]},
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53]},
      {stage3_28[8],stage3_27[19],stage3_26[19],stage3_25[30],stage3_24[35]}
   );
   gpc606_5 gpc3501 (
      {stage2_24[71], stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76]},
      {stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59]},
      {stage3_28[9],stage3_27[20],stage3_26[20],stage3_25[31],stage3_24[36]}
   );
   gpc606_5 gpc3502 (
      {stage2_24[77], stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82]},
      {stage2_26[60], stage2_26[61], stage2_26[62], stage2_26[63], stage2_26[64], stage2_26[65]},
      {stage3_28[10],stage3_27[21],stage3_26[21],stage3_25[32],stage3_24[37]}
   );
   gpc606_5 gpc3503 (
      {stage2_24[83], stage2_24[84], stage2_24[85], stage2_24[86], stage2_24[87], stage2_24[88]},
      {stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71]},
      {stage3_28[11],stage3_27[22],stage3_26[22],stage3_25[33],stage3_24[38]}
   );
   gpc606_5 gpc3504 (
      {stage2_24[89], stage2_24[90], stage2_24[91], stage2_24[92], stage2_24[93], stage2_24[94]},
      {stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76], stage2_26[77]},
      {stage3_28[12],stage3_27[23],stage3_26[23],stage3_25[34],stage3_24[39]}
   );
   gpc606_5 gpc3505 (
      {stage2_24[95], stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], 1'b0},
      {stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage3_28[13],stage3_27[24],stage3_26[24],stage3_25[35],stage3_24[40]}
   );
   gpc606_5 gpc3506 (
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[14],stage3_27[25],stage3_26[25],stage3_25[36]}
   );
   gpc606_5 gpc3507 (
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[15],stage3_27[26],stage3_26[26],stage3_25[37]}
   );
   gpc606_5 gpc3508 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[16],stage3_27[27],stage3_26[27],stage3_25[38]}
   );
   gpc606_5 gpc3509 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], 1'b0, 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[17],stage3_27[28],stage3_26[28],stage3_25[39]}
   );
   gpc615_5 gpc3510 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88]},
      {stage2_27[24]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[4],stage3_28[18],stage3_27[29],stage3_26[29]}
   );
   gpc615_5 gpc3511 (
      {stage2_26[89], stage2_26[90], stage2_26[91], stage2_26[92], stage2_26[93]},
      {stage2_27[25]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[5],stage3_28[19],stage3_27[30],stage3_26[30]}
   );
   gpc615_5 gpc3512 (
      {stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97], stage2_26[98]},
      {stage2_27[26]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[6],stage3_28[20],stage3_27[31],stage3_26[31]}
   );
   gpc606_5 gpc3513 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[3],stage3_29[7],stage3_28[21],stage3_27[32]}
   );
   gpc606_5 gpc3514 (
      {stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[4],stage3_29[8],stage3_28[22],stage3_27[33]}
   );
   gpc606_5 gpc3515 (
      {stage2_27[39], stage2_27[40], stage2_27[41], stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[5],stage3_29[9],stage3_28[23],stage3_27[34]}
   );
   gpc615_5 gpc3516 (
      {stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48], stage2_27[49]},
      {stage2_28[18]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[6],stage3_29[10],stage3_28[24],stage3_27[35]}
   );
   gpc615_5 gpc3517 (
      {stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54]},
      {stage2_28[19]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[7],stage3_29[11],stage3_28[25],stage3_27[36]}
   );
   gpc615_5 gpc3518 (
      {stage2_27[55], stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[20]},
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage3_31[5],stage3_30[8],stage3_29[12],stage3_28[26],stage3_27[37]}
   );
   gpc615_5 gpc3519 (
      {stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63], stage2_27[64]},
      {stage2_28[21]},
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage3_31[6],stage3_30[9],stage3_29[13],stage3_28[27],stage3_27[38]}
   );
   gpc615_5 gpc3520 (
      {stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_28[22]},
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage3_31[7],stage3_30[10],stage3_29[14],stage3_28[28],stage3_27[39]}
   );
   gpc606_5 gpc3521 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[8],stage3_30[11],stage3_29[15],stage3_28[29]}
   );
   gpc606_5 gpc3522 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[9],stage3_30[12],stage3_29[16],stage3_28[30]}
   );
   gpc606_5 gpc3523 (
      {stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[10],stage3_30[13],stage3_29[17],stage3_28[31]}
   );
   gpc606_5 gpc3524 (
      {stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[11],stage3_30[14],stage3_29[18],stage3_28[32]}
   );
   gpc606_5 gpc3525 (
      {stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[12],stage3_30[15],stage3_29[19],stage3_28[33]}
   );
   gpc606_5 gpc3526 (
      {stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[13],stage3_30[16],stage3_29[20],stage3_28[34]}
   );
   gpc615_5 gpc3527 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[48]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[14],stage3_30[17],stage3_29[21],stage3_28[35]}
   );
   gpc615_5 gpc3528 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[49]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[15],stage3_30[18],stage3_29[22],stage3_28[36]}
   );
   gpc1163_5 gpc3529 (
      {stage2_29[50], stage2_29[51], stage2_29[52]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[8],stage3_31[16],stage3_30[19],stage3_29[23]}
   );
   gpc1163_5 gpc3530 (
      {stage2_29[53], stage2_29[54], stage2_29[55]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[9],stage3_31[17],stage3_30[20],stage3_29[24]}
   );
   gpc1163_5 gpc3531 (
      {stage2_29[56], stage2_29[57], stage2_29[58]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[10],stage3_31[18],stage3_30[21],stage3_29[25]}
   );
   gpc1163_5 gpc3532 (
      {stage2_29[59], stage2_29[60], stage2_29[61]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[11],stage3_31[19],stage3_30[22],stage3_29[26]}
   );
   gpc1163_5 gpc3533 (
      {stage2_29[62], stage2_29[63], stage2_29[64]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[12],stage3_31[20],stage3_30[23],stage3_29[27]}
   );
   gpc606_5 gpc3534 (
      {stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[13],stage3_31[21],stage3_30[24],stage3_29[28]}
   );
   gpc606_5 gpc3535 (
      {stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[14],stage3_31[22],stage3_30[25],stage3_29[29]}
   );
   gpc606_5 gpc3536 (
      {stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[15],stage3_31[23],stage3_30[26],stage3_29[30]}
   );
   gpc606_5 gpc3537 (
      {stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[16],stage3_31[24],stage3_30[27],stage3_29[31]}
   );
   gpc606_5 gpc3538 (
      {stage2_29[89], stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[17],stage3_31[25],stage3_30[28],stage3_29[32]}
   );
   gpc606_5 gpc3539 (
      {stage2_29[95], stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[18],stage3_31[26],stage3_30[29],stage3_29[33]}
   );
   gpc606_5 gpc3540 (
      {stage2_29[101], stage2_29[102], stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[19],stage3_31[27],stage3_30[30],stage3_29[34]}
   );
   gpc606_5 gpc3541 (
      {stage2_29[107], stage2_29[108], stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[20],stage3_31[28],stage3_30[31],stage3_29[35]}
   );
   gpc606_5 gpc3542 (
      {stage2_29[113], stage2_29[114], stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[21],stage3_31[29],stage3_30[32],stage3_29[36]}
   );
   gpc606_5 gpc3543 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_32[5], stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10]},
      {stage3_34[0],stage3_33[14],stage3_32[22],stage3_31[30],stage3_30[33]}
   );
   gpc606_5 gpc3544 (
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_32[11], stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16]},
      {stage3_34[1],stage3_33[15],stage3_32[23],stage3_31[31],stage3_30[34]}
   );
   gpc606_5 gpc3545 (
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22]},
      {stage3_34[2],stage3_33[16],stage3_32[24],stage3_31[32],stage3_30[35]}
   );
   gpc606_5 gpc3546 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101]},
      {stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28]},
      {stage3_34[3],stage3_33[17],stage3_32[25],stage3_31[33],stage3_30[36]}
   );
   gpc606_5 gpc3547 (
      {stage2_30[102], stage2_30[103], stage2_30[104], stage2_30[105], stage2_30[106], stage2_30[107]},
      {stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34]},
      {stage3_34[4],stage3_33[18],stage3_32[26],stage3_31[34],stage3_30[37]}
   );
   gpc606_5 gpc3548 (
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[5],stage3_33[19],stage3_32[27],stage3_31[35]}
   );
   gpc606_5 gpc3549 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[6],stage3_33[20],stage3_32[28],stage3_31[36]}
   );
   gpc606_5 gpc3550 (
      {stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[7],stage3_33[21],stage3_32[29],stage3_31[37]}
   );
   gpc606_5 gpc3551 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[8],stage3_33[22],stage3_32[30],stage3_31[38]}
   );
   gpc606_5 gpc3552 (
      {stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[9],stage3_33[23],stage3_32[31]}
   );
   gpc606_5 gpc3553 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45], stage2_32[46]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[10],stage3_33[24],stage3_32[32]}
   );
   gpc606_5 gpc3554 (
      {stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50], stage2_32[51], stage2_32[52]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[6],stage3_34[11],stage3_33[25],stage3_32[33]}
   );
   gpc606_5 gpc3555 (
      {stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56], stage2_32[57], stage2_32[58]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[7],stage3_34[12],stage3_33[26],stage3_32[34]}
   );
   gpc606_5 gpc3556 (
      {stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62], stage2_32[63], stage2_32[64]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[8],stage3_34[13],stage3_33[27],stage3_32[35]}
   );
   gpc606_5 gpc3557 (
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[5],stage3_35[9],stage3_34[14],stage3_33[28]}
   );
   gpc606_5 gpc3558 (
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[6],stage3_35[10],stage3_34[15],stage3_33[29]}
   );
   gpc1_1 gpc3559 (
      {stage2_0[21]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3560 (
      {stage2_2[43]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3561 (
      {stage2_2[44]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3562 (
      {stage2_2[45]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3563 (
      {stage2_2[46]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3564 (
      {stage2_2[47]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3565 (
      {stage2_2[48]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3566 (
      {stage2_2[49]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3567 (
      {stage2_2[50]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3568 (
      {stage2_4[82]},
      {stage3_4[35]}
   );
   gpc1_1 gpc3569 (
      {stage2_4[83]},
      {stage3_4[36]}
   );
   gpc1_1 gpc3570 (
      {stage2_4[84]},
      {stage3_4[37]}
   );
   gpc1_1 gpc3571 (
      {stage2_4[85]},
      {stage3_4[38]}
   );
   gpc1_1 gpc3572 (
      {stage2_4[86]},
      {stage3_4[39]}
   );
   gpc1_1 gpc3573 (
      {stage2_4[87]},
      {stage3_4[40]}
   );
   gpc1_1 gpc3574 (
      {stage2_4[88]},
      {stage3_4[41]}
   );
   gpc1_1 gpc3575 (
      {stage2_4[89]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3576 (
      {stage2_4[90]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3577 (
      {stage2_5[71]},
      {stage3_5[36]}
   );
   gpc1_1 gpc3578 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3579 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3580 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3581 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3582 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3583 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3584 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3585 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3586 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3587 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3588 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3589 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3590 (
      {stage2_6[83]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3591 (
      {stage2_6[84]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3592 (
      {stage2_6[85]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3593 (
      {stage2_6[86]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3594 (
      {stage2_6[87]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3595 (
      {stage2_6[88]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3596 (
      {stage2_6[89]},
      {stage3_6[38]}
   );
   gpc1_1 gpc3597 (
      {stage2_6[90]},
      {stage3_6[39]}
   );
   gpc1_1 gpc3598 (
      {stage2_6[91]},
      {stage3_6[40]}
   );
   gpc1_1 gpc3599 (
      {stage2_6[92]},
      {stage3_6[41]}
   );
   gpc1_1 gpc3600 (
      {stage2_6[93]},
      {stage3_6[42]}
   );
   gpc1_1 gpc3601 (
      {stage2_7[70]},
      {stage3_7[29]}
   );
   gpc1_1 gpc3602 (
      {stage2_7[71]},
      {stage3_7[30]}
   );
   gpc1_1 gpc3603 (
      {stage2_7[72]},
      {stage3_7[31]}
   );
   gpc1_1 gpc3604 (
      {stage2_7[73]},
      {stage3_7[32]}
   );
   gpc1_1 gpc3605 (
      {stage2_7[74]},
      {stage3_7[33]}
   );
   gpc1_1 gpc3606 (
      {stage2_7[75]},
      {stage3_7[34]}
   );
   gpc1_1 gpc3607 (
      {stage2_7[76]},
      {stage3_7[35]}
   );
   gpc1_1 gpc3608 (
      {stage2_7[77]},
      {stage3_7[36]}
   );
   gpc1_1 gpc3609 (
      {stage2_7[78]},
      {stage3_7[37]}
   );
   gpc1_1 gpc3610 (
      {stage2_7[79]},
      {stage3_7[38]}
   );
   gpc1_1 gpc3611 (
      {stage2_7[80]},
      {stage3_7[39]}
   );
   gpc1_1 gpc3612 (
      {stage2_7[81]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3613 (
      {stage2_7[82]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3614 (
      {stage2_7[83]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3615 (
      {stage2_7[84]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3616 (
      {stage2_7[85]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3617 (
      {stage2_7[86]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3618 (
      {stage2_7[87]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3619 (
      {stage2_7[88]},
      {stage3_7[47]}
   );
   gpc1_1 gpc3620 (
      {stage2_7[89]},
      {stage3_7[48]}
   );
   gpc1_1 gpc3621 (
      {stage2_7[90]},
      {stage3_7[49]}
   );
   gpc1_1 gpc3622 (
      {stage2_7[91]},
      {stage3_7[50]}
   );
   gpc1_1 gpc3623 (
      {stage2_7[92]},
      {stage3_7[51]}
   );
   gpc1_1 gpc3624 (
      {stage2_7[93]},
      {stage3_7[52]}
   );
   gpc1_1 gpc3625 (
      {stage2_7[94]},
      {stage3_7[53]}
   );
   gpc1_1 gpc3626 (
      {stage2_7[95]},
      {stage3_7[54]}
   );
   gpc1_1 gpc3627 (
      {stage2_7[96]},
      {stage3_7[55]}
   );
   gpc1_1 gpc3628 (
      {stage2_7[97]},
      {stage3_7[56]}
   );
   gpc1_1 gpc3629 (
      {stage2_7[98]},
      {stage3_7[57]}
   );
   gpc1_1 gpc3630 (
      {stage2_7[99]},
      {stage3_7[58]}
   );
   gpc1_1 gpc3631 (
      {stage2_7[100]},
      {stage3_7[59]}
   );
   gpc1_1 gpc3632 (
      {stage2_7[101]},
      {stage3_7[60]}
   );
   gpc1_1 gpc3633 (
      {stage2_7[102]},
      {stage3_7[61]}
   );
   gpc1_1 gpc3634 (
      {stage2_7[103]},
      {stage3_7[62]}
   );
   gpc1_1 gpc3635 (
      {stage2_7[104]},
      {stage3_7[63]}
   );
   gpc1_1 gpc3636 (
      {stage2_7[105]},
      {stage3_7[64]}
   );
   gpc1_1 gpc3637 (
      {stage2_7[106]},
      {stage3_7[65]}
   );
   gpc1_1 gpc3638 (
      {stage2_7[107]},
      {stage3_7[66]}
   );
   gpc1_1 gpc3639 (
      {stage2_7[108]},
      {stage3_7[67]}
   );
   gpc1_1 gpc3640 (
      {stage2_7[109]},
      {stage3_7[68]}
   );
   gpc1_1 gpc3641 (
      {stage2_9[36]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3642 (
      {stage2_9[37]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3643 (
      {stage2_9[38]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3644 (
      {stage2_9[39]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3645 (
      {stage2_9[40]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3646 (
      {stage2_9[41]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3647 (
      {stage2_9[42]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3648 (
      {stage2_9[43]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3649 (
      {stage2_9[44]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3650 (
      {stage2_9[45]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3651 (
      {stage2_9[46]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3652 (
      {stage2_9[47]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3653 (
      {stage2_9[48]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[49]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[50]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[51]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[52]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3658 (
      {stage2_9[53]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3659 (
      {stage2_9[54]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3660 (
      {stage2_9[55]},
      {stage3_9[50]}
   );
   gpc1_1 gpc3661 (
      {stage2_9[56]},
      {stage3_9[51]}
   );
   gpc1_1 gpc3662 (
      {stage2_9[57]},
      {stage3_9[52]}
   );
   gpc1_1 gpc3663 (
      {stage2_9[58]},
      {stage3_9[53]}
   );
   gpc1_1 gpc3664 (
      {stage2_9[59]},
      {stage3_9[54]}
   );
   gpc1_1 gpc3665 (
      {stage2_9[60]},
      {stage3_9[55]}
   );
   gpc1_1 gpc3666 (
      {stage2_9[61]},
      {stage3_9[56]}
   );
   gpc1_1 gpc3667 (
      {stage2_9[62]},
      {stage3_9[57]}
   );
   gpc1_1 gpc3668 (
      {stage2_9[63]},
      {stage3_9[58]}
   );
   gpc1_1 gpc3669 (
      {stage2_9[64]},
      {stage3_9[59]}
   );
   gpc1_1 gpc3670 (
      {stage2_9[65]},
      {stage3_9[60]}
   );
   gpc1_1 gpc3671 (
      {stage2_9[66]},
      {stage3_9[61]}
   );
   gpc1_1 gpc3672 (
      {stage2_9[67]},
      {stage3_9[62]}
   );
   gpc1_1 gpc3673 (
      {stage2_9[68]},
      {stage3_9[63]}
   );
   gpc1_1 gpc3674 (
      {stage2_9[69]},
      {stage3_9[64]}
   );
   gpc1_1 gpc3675 (
      {stage2_9[70]},
      {stage3_9[65]}
   );
   gpc1_1 gpc3676 (
      {stage2_9[71]},
      {stage3_9[66]}
   );
   gpc1_1 gpc3677 (
      {stage2_9[72]},
      {stage3_9[67]}
   );
   gpc1_1 gpc3678 (
      {stage2_9[73]},
      {stage3_9[68]}
   );
   gpc1_1 gpc3679 (
      {stage2_9[74]},
      {stage3_9[69]}
   );
   gpc1_1 gpc3680 (
      {stage2_10[88]},
      {stage3_10[28]}
   );
   gpc1_1 gpc3681 (
      {stage2_11[80]},
      {stage3_11[32]}
   );
   gpc1_1 gpc3682 (
      {stage2_11[81]},
      {stage3_11[33]}
   );
   gpc1_1 gpc3683 (
      {stage2_11[82]},
      {stage3_11[34]}
   );
   gpc1_1 gpc3684 (
      {stage2_11[83]},
      {stage3_11[35]}
   );
   gpc1_1 gpc3685 (
      {stage2_11[84]},
      {stage3_11[36]}
   );
   gpc1_1 gpc3686 (
      {stage2_11[85]},
      {stage3_11[37]}
   );
   gpc1_1 gpc3687 (
      {stage2_11[86]},
      {stage3_11[38]}
   );
   gpc1_1 gpc3688 (
      {stage2_11[87]},
      {stage3_11[39]}
   );
   gpc1_1 gpc3689 (
      {stage2_11[88]},
      {stage3_11[40]}
   );
   gpc1_1 gpc3690 (
      {stage2_11[89]},
      {stage3_11[41]}
   );
   gpc1_1 gpc3691 (
      {stage2_11[90]},
      {stage3_11[42]}
   );
   gpc1_1 gpc3692 (
      {stage2_11[91]},
      {stage3_11[43]}
   );
   gpc1_1 gpc3693 (
      {stage2_12[102]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3694 (
      {stage2_13[95]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3695 (
      {stage2_13[96]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3696 (
      {stage2_13[97]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3697 (
      {stage2_13[98]},
      {stage3_13[37]}
   );
   gpc1_1 gpc3698 (
      {stage2_13[99]},
      {stage3_13[38]}
   );
   gpc1_1 gpc3699 (
      {stage2_13[100]},
      {stage3_13[39]}
   );
   gpc1_1 gpc3700 (
      {stage2_13[101]},
      {stage3_13[40]}
   );
   gpc1_1 gpc3701 (
      {stage2_14[133]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3702 (
      {stage2_14[134]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3703 (
      {stage2_14[135]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3704 (
      {stage2_14[136]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3705 (
      {stage2_14[137]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3706 (
      {stage2_14[138]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[95]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[96]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[97]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[98]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[99]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[100]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[101]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[102]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[103]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[104]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3717 (
      {stage2_15[105]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3718 (
      {stage2_15[106]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3719 (
      {stage2_15[107]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3720 (
      {stage2_15[108]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3721 (
      {stage2_15[109]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3722 (
      {stage2_15[110]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3723 (
      {stage2_15[111]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3724 (
      {stage2_15[112]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3725 (
      {stage2_15[113]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3726 (
      {stage2_15[114]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3727 (
      {stage2_15[115]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3728 (
      {stage2_15[116]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3729 (
      {stage2_15[117]},
      {stage3_15[71]}
   );
   gpc1_1 gpc3730 (
      {stage2_15[118]},
      {stage3_15[72]}
   );
   gpc1_1 gpc3731 (
      {stage2_15[119]},
      {stage3_15[73]}
   );
   gpc1_1 gpc3732 (
      {stage2_15[120]},
      {stage3_15[74]}
   );
   gpc1_1 gpc3733 (
      {stage2_15[121]},
      {stage3_15[75]}
   );
   gpc1_1 gpc3734 (
      {stage2_15[122]},
      {stage3_15[76]}
   );
   gpc1_1 gpc3735 (
      {stage2_15[123]},
      {stage3_15[77]}
   );
   gpc1_1 gpc3736 (
      {stage2_15[124]},
      {stage3_15[78]}
   );
   gpc1_1 gpc3737 (
      {stage2_15[125]},
      {stage3_15[79]}
   );
   gpc1_1 gpc3738 (
      {stage2_15[126]},
      {stage3_15[80]}
   );
   gpc1_1 gpc3739 (
      {stage2_15[127]},
      {stage3_15[81]}
   );
   gpc1_1 gpc3740 (
      {stage2_15[128]},
      {stage3_15[82]}
   );
   gpc1_1 gpc3741 (
      {stage2_15[129]},
      {stage3_15[83]}
   );
   gpc1_1 gpc3742 (
      {stage2_15[130]},
      {stage3_15[84]}
   );
   gpc1_1 gpc3743 (
      {stage2_15[131]},
      {stage3_15[85]}
   );
   gpc1_1 gpc3744 (
      {stage2_15[132]},
      {stage3_15[86]}
   );
   gpc1_1 gpc3745 (
      {stage2_15[133]},
      {stage3_15[87]}
   );
   gpc1_1 gpc3746 (
      {stage2_15[134]},
      {stage3_15[88]}
   );
   gpc1_1 gpc3747 (
      {stage2_15[135]},
      {stage3_15[89]}
   );
   gpc1_1 gpc3748 (
      {stage2_16[81]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3749 (
      {stage2_16[82]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3750 (
      {stage2_16[83]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3751 (
      {stage2_16[84]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3752 (
      {stage2_16[85]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3753 (
      {stage2_16[86]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3754 (
      {stage2_16[87]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3755 (
      {stage2_16[88]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3756 (
      {stage2_16[89]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3757 (
      {stage2_16[90]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3758 (
      {stage2_16[91]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3759 (
      {stage2_16[92]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3760 (
      {stage2_16[93]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3761 (
      {stage2_16[94]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3762 (
      {stage2_16[95]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3763 (
      {stage2_16[96]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3764 (
      {stage2_16[97]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3765 (
      {stage2_16[98]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3766 (
      {stage2_16[99]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3767 (
      {stage2_16[100]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3768 (
      {stage2_16[101]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3769 (
      {stage2_16[102]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3770 (
      {stage2_16[103]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3771 (
      {stage2_17[109]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3772 (
      {stage2_17[110]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3773 (
      {stage2_17[111]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3774 (
      {stage2_17[112]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3775 (
      {stage2_17[113]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3776 (
      {stage2_17[114]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3777 (
      {stage2_17[115]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3778 (
      {stage2_17[116]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3779 (
      {stage2_17[117]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3780 (
      {stage2_17[118]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3781 (
      {stage2_17[119]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3782 (
      {stage2_17[120]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3783 (
      {stage2_17[121]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3784 (
      {stage2_18[80]},
      {stage3_18[48]}
   );
   gpc1_1 gpc3785 (
      {stage2_18[81]},
      {stage3_18[49]}
   );
   gpc1_1 gpc3786 (
      {stage2_19[98]},
      {stage3_19[38]}
   );
   gpc1_1 gpc3787 (
      {stage2_19[99]},
      {stage3_19[39]}
   );
   gpc1_1 gpc3788 (
      {stage2_19[100]},
      {stage3_19[40]}
   );
   gpc1_1 gpc3789 (
      {stage2_19[101]},
      {stage3_19[41]}
   );
   gpc1_1 gpc3790 (
      {stage2_19[102]},
      {stage3_19[42]}
   );
   gpc1_1 gpc3791 (
      {stage2_19[103]},
      {stage3_19[43]}
   );
   gpc1_1 gpc3792 (
      {stage2_19[104]},
      {stage3_19[44]}
   );
   gpc1_1 gpc3793 (
      {stage2_19[105]},
      {stage3_19[45]}
   );
   gpc1_1 gpc3794 (
      {stage2_19[106]},
      {stage3_19[46]}
   );
   gpc1_1 gpc3795 (
      {stage2_19[107]},
      {stage3_19[47]}
   );
   gpc1_1 gpc3796 (
      {stage2_19[108]},
      {stage3_19[48]}
   );
   gpc1_1 gpc3797 (
      {stage2_19[109]},
      {stage3_19[49]}
   );
   gpc1_1 gpc3798 (
      {stage2_20[116]},
      {stage3_20[34]}
   );
   gpc1_1 gpc3799 (
      {stage2_20[117]},
      {stage3_20[35]}
   );
   gpc1_1 gpc3800 (
      {stage2_20[118]},
      {stage3_20[36]}
   );
   gpc1_1 gpc3801 (
      {stage2_20[119]},
      {stage3_20[37]}
   );
   gpc1_1 gpc3802 (
      {stage2_20[120]},
      {stage3_20[38]}
   );
   gpc1_1 gpc3803 (
      {stage2_20[121]},
      {stage3_20[39]}
   );
   gpc1_1 gpc3804 (
      {stage2_20[122]},
      {stage3_20[40]}
   );
   gpc1_1 gpc3805 (
      {stage2_20[123]},
      {stage3_20[41]}
   );
   gpc1_1 gpc3806 (
      {stage2_20[124]},
      {stage3_20[42]}
   );
   gpc1_1 gpc3807 (
      {stage2_20[125]},
      {stage3_20[43]}
   );
   gpc1_1 gpc3808 (
      {stage2_20[126]},
      {stage3_20[44]}
   );
   gpc1_1 gpc3809 (
      {stage2_20[127]},
      {stage3_20[45]}
   );
   gpc1_1 gpc3810 (
      {stage2_21[64]},
      {stage3_21[44]}
   );
   gpc1_1 gpc3811 (
      {stage2_21[65]},
      {stage3_21[45]}
   );
   gpc1_1 gpc3812 (
      {stage2_21[66]},
      {stage3_21[46]}
   );
   gpc1_1 gpc3813 (
      {stage2_21[67]},
      {stage3_21[47]}
   );
   gpc1_1 gpc3814 (
      {stage2_21[68]},
      {stage3_21[48]}
   );
   gpc1_1 gpc3815 (
      {stage2_21[69]},
      {stage3_21[49]}
   );
   gpc1_1 gpc3816 (
      {stage2_21[70]},
      {stage3_21[50]}
   );
   gpc1_1 gpc3817 (
      {stage2_21[71]},
      {stage3_21[51]}
   );
   gpc1_1 gpc3818 (
      {stage2_21[72]},
      {stage3_21[52]}
   );
   gpc1_1 gpc3819 (
      {stage2_21[73]},
      {stage3_21[53]}
   );
   gpc1_1 gpc3820 (
      {stage2_21[74]},
      {stage3_21[54]}
   );
   gpc1_1 gpc3821 (
      {stage2_21[75]},
      {stage3_21[55]}
   );
   gpc1_1 gpc3822 (
      {stage2_21[76]},
      {stage3_21[56]}
   );
   gpc1_1 gpc3823 (
      {stage2_21[77]},
      {stage3_21[57]}
   );
   gpc1_1 gpc3824 (
      {stage2_21[78]},
      {stage3_21[58]}
   );
   gpc1_1 gpc3825 (
      {stage2_22[66]},
      {stage3_22[34]}
   );
   gpc1_1 gpc3826 (
      {stage2_22[67]},
      {stage3_22[35]}
   );
   gpc1_1 gpc3827 (
      {stage2_22[68]},
      {stage3_22[36]}
   );
   gpc1_1 gpc3828 (
      {stage2_22[69]},
      {stage3_22[37]}
   );
   gpc1_1 gpc3829 (
      {stage2_22[70]},
      {stage3_22[38]}
   );
   gpc1_1 gpc3830 (
      {stage2_22[71]},
      {stage3_22[39]}
   );
   gpc1_1 gpc3831 (
      {stage2_22[72]},
      {stage3_22[40]}
   );
   gpc1_1 gpc3832 (
      {stage2_22[73]},
      {stage3_22[41]}
   );
   gpc1_1 gpc3833 (
      {stage2_22[74]},
      {stage3_22[42]}
   );
   gpc1_1 gpc3834 (
      {stage2_22[75]},
      {stage3_22[43]}
   );
   gpc1_1 gpc3835 (
      {stage2_22[76]},
      {stage3_22[44]}
   );
   gpc1_1 gpc3836 (
      {stage2_22[77]},
      {stage3_22[45]}
   );
   gpc1_1 gpc3837 (
      {stage2_22[78]},
      {stage3_22[46]}
   );
   gpc1_1 gpc3838 (
      {stage2_23[91]},
      {stage3_23[29]}
   );
   gpc1_1 gpc3839 (
      {stage2_23[92]},
      {stage3_23[30]}
   );
   gpc1_1 gpc3840 (
      {stage2_23[93]},
      {stage3_23[31]}
   );
   gpc1_1 gpc3841 (
      {stage2_23[94]},
      {stage3_23[32]}
   );
   gpc1_1 gpc3842 (
      {stage2_23[95]},
      {stage3_23[33]}
   );
   gpc1_1 gpc3843 (
      {stage2_23[96]},
      {stage3_23[34]}
   );
   gpc1_1 gpc3844 (
      {stage2_23[97]},
      {stage3_23[35]}
   );
   gpc1_1 gpc3845 (
      {stage2_23[98]},
      {stage3_23[36]}
   );
   gpc1_1 gpc3846 (
      {stage2_23[99]},
      {stage3_23[37]}
   );
   gpc1_1 gpc3847 (
      {stage2_23[100]},
      {stage3_23[38]}
   );
   gpc1_1 gpc3848 (
      {stage2_23[101]},
      {stage3_23[39]}
   );
   gpc1_1 gpc3849 (
      {stage2_23[102]},
      {stage3_23[40]}
   );
   gpc1_1 gpc3850 (
      {stage2_23[103]},
      {stage3_23[41]}
   );
   gpc1_1 gpc3851 (
      {stage2_23[104]},
      {stage3_23[42]}
   );
   gpc1_1 gpc3852 (
      {stage2_23[105]},
      {stage3_23[43]}
   );
   gpc1_1 gpc3853 (
      {stage2_23[106]},
      {stage3_23[44]}
   );
   gpc1_1 gpc3854 (
      {stage2_23[107]},
      {stage3_23[45]}
   );
   gpc1_1 gpc3855 (
      {stage2_23[108]},
      {stage3_23[46]}
   );
   gpc1_1 gpc3856 (
      {stage2_23[109]},
      {stage3_23[47]}
   );
   gpc1_1 gpc3857 (
      {stage2_27[70]},
      {stage3_27[40]}
   );
   gpc1_1 gpc3858 (
      {stage2_27[71]},
      {stage3_27[41]}
   );
   gpc1_1 gpc3859 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc3860 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc3861 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc3862 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc3863 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc3864 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc3865 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc3866 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc3867 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc3868 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc3869 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc3870 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc3871 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc3872 (
      {stage2_27[85]},
      {stage3_27[55]}
   );
   gpc1_1 gpc3873 (
      {stage2_27[86]},
      {stage3_27[56]}
   );
   gpc1_1 gpc3874 (
      {stage2_27[87]},
      {stage3_27[57]}
   );
   gpc1_1 gpc3875 (
      {stage2_27[88]},
      {stage3_27[58]}
   );
   gpc1_1 gpc3876 (
      {stage2_27[89]},
      {stage3_27[59]}
   );
   gpc1_1 gpc3877 (
      {stage2_27[90]},
      {stage3_27[60]}
   );
   gpc1_1 gpc3878 (
      {stage2_27[91]},
      {stage3_27[61]}
   );
   gpc1_1 gpc3879 (
      {stage2_27[92]},
      {stage3_27[62]}
   );
   gpc1_1 gpc3880 (
      {stage2_27[93]},
      {stage3_27[63]}
   );
   gpc1_1 gpc3881 (
      {stage2_27[94]},
      {stage3_27[64]}
   );
   gpc1_1 gpc3882 (
      {stage2_27[95]},
      {stage3_27[65]}
   );
   gpc1_1 gpc3883 (
      {stage2_27[96]},
      {stage3_27[66]}
   );
   gpc1_1 gpc3884 (
      {stage2_28[69]},
      {stage3_28[37]}
   );
   gpc1_1 gpc3885 (
      {stage2_28[70]},
      {stage3_28[38]}
   );
   gpc1_1 gpc3886 (
      {stage2_28[71]},
      {stage3_28[39]}
   );
   gpc1_1 gpc3887 (
      {stage2_28[72]},
      {stage3_28[40]}
   );
   gpc1_1 gpc3888 (
      {stage2_28[73]},
      {stage3_28[41]}
   );
   gpc1_1 gpc3889 (
      {stage2_28[74]},
      {stage3_28[42]}
   );
   gpc1_1 gpc3890 (
      {stage2_29[119]},
      {stage3_29[37]}
   );
   gpc1_1 gpc3891 (
      {stage2_29[120]},
      {stage3_29[38]}
   );
   gpc1_1 gpc3892 (
      {stage2_30[108]},
      {stage3_30[38]}
   );
   gpc1_1 gpc3893 (
      {stage2_30[109]},
      {stage3_30[39]}
   );
   gpc1_1 gpc3894 (
      {stage2_30[110]},
      {stage3_30[40]}
   );
   gpc1_1 gpc3895 (
      {stage2_30[111]},
      {stage3_30[41]}
   );
   gpc1_1 gpc3896 (
      {stage2_30[112]},
      {stage3_30[42]}
   );
   gpc1_1 gpc3897 (
      {stage2_30[113]},
      {stage3_30[43]}
   );
   gpc1_1 gpc3898 (
      {stage2_30[114]},
      {stage3_30[44]}
   );
   gpc1_1 gpc3899 (
      {stage2_30[115]},
      {stage3_30[45]}
   );
   gpc1_1 gpc3900 (
      {stage2_30[116]},
      {stage3_30[46]}
   );
   gpc1_1 gpc3901 (
      {stage2_30[117]},
      {stage3_30[47]}
   );
   gpc1_1 gpc3902 (
      {stage2_30[118]},
      {stage3_30[48]}
   );
   gpc1_1 gpc3903 (
      {stage2_30[119]},
      {stage3_30[49]}
   );
   gpc1_1 gpc3904 (
      {stage2_30[120]},
      {stage3_30[50]}
   );
   gpc1_1 gpc3905 (
      {stage2_30[121]},
      {stage3_30[51]}
   );
   gpc1_1 gpc3906 (
      {stage2_30[122]},
      {stage3_30[52]}
   );
   gpc1_1 gpc3907 (
      {stage2_30[123]},
      {stage3_30[53]}
   );
   gpc1_1 gpc3908 (
      {stage2_30[124]},
      {stage3_30[54]}
   );
   gpc1_1 gpc3909 (
      {stage2_30[125]},
      {stage3_30[55]}
   );
   gpc1_1 gpc3910 (
      {stage2_30[126]},
      {stage3_30[56]}
   );
   gpc1_1 gpc3911 (
      {stage2_30[127]},
      {stage3_30[57]}
   );
   gpc1_1 gpc3912 (
      {stage2_30[128]},
      {stage3_30[58]}
   );
   gpc1_1 gpc3913 (
      {stage2_30[129]},
      {stage3_30[59]}
   );
   gpc1_1 gpc3914 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc3915 (
      {stage2_33[36]},
      {stage3_33[30]}
   );
   gpc1_1 gpc3916 (
      {stage2_33[37]},
      {stage3_33[31]}
   );
   gpc1_1 gpc3917 (
      {stage2_33[38]},
      {stage3_33[32]}
   );
   gpc1_1 gpc3918 (
      {stage2_33[39]},
      {stage3_33[33]}
   );
   gpc1_1 gpc3919 (
      {stage2_33[40]},
      {stage3_33[34]}
   );
   gpc1_1 gpc3920 (
      {stage2_33[41]},
      {stage3_33[35]}
   );
   gpc1_1 gpc3921 (
      {stage2_33[42]},
      {stage3_33[36]}
   );
   gpc1_1 gpc3922 (
      {stage2_33[43]},
      {stage3_33[37]}
   );
   gpc1_1 gpc3923 (
      {stage2_33[44]},
      {stage3_33[38]}
   );
   gpc1_1 gpc3924 (
      {stage2_33[45]},
      {stage3_33[39]}
   );
   gpc1_1 gpc3925 (
      {stage2_34[30]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3926 (
      {stage2_34[31]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3927 (
      {stage2_34[32]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3928 (
      {stage2_34[33]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3929 (
      {stage2_34[34]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3930 (
      {stage2_34[35]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3931 (
      {stage2_35[12]},
      {stage3_35[11]}
   );
   gpc1_1 gpc3932 (
      {stage2_35[13]},
      {stage3_35[12]}
   );
   gpc606_5 gpc3933 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc3934 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc3935 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc3936 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc3937 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc3938 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc3939 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc615_5 gpc3940 (
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc3941 (
      {stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21]},
      {stage3_4[25]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[5],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc3942 (
      {stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25], stage3_3[26]},
      {stage3_4[26]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[6],stage4_5[8],stage4_4[9],stage4_3[9]}
   );
   gpc606_5 gpc3943 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[7],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc3944 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[8],stage4_5[10],stage4_4[11]}
   );
   gpc1163_5 gpc3945 (
      {stage3_5[18], stage3_5[19], stage3_5[20]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[0]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[2],stage4_7[5],stage4_6[9],stage4_5[11]}
   );
   gpc1163_5 gpc3946 (
      {stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[1]},
      {stage3_8[1]},
      {stage4_9[1],stage4_8[3],stage4_7[6],stage4_6[10],stage4_5[12]}
   );
   gpc606_5 gpc3947 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage4_9[2],stage4_8[4],stage4_7[7],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc3948 (
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage4_9[3],stage4_8[5],stage4_7[8],stage4_6[12],stage4_5[14]}
   );
   gpc606_5 gpc3949 (
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage4_9[4],stage4_8[6],stage4_7[9],stage4_6[13],stage4_5[15]}
   );
   gpc615_5 gpc3950 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[20]},
      {stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6], stage3_8[7]},
      {stage4_10[0],stage4_9[5],stage4_8[7],stage4_7[10],stage4_6[14]}
   );
   gpc615_5 gpc3951 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[21]},
      {stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13]},
      {stage4_10[1],stage4_9[6],stage4_8[8],stage4_7[11],stage4_6[15]}
   );
   gpc615_5 gpc3952 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[22]},
      {stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19]},
      {stage4_10[2],stage4_9[7],stage4_8[9],stage4_7[12],stage4_6[16]}
   );
   gpc615_5 gpc3953 (
      {stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27]},
      {stage3_8[20]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[8],stage4_8[10],stage4_7[13]}
   );
   gpc615_5 gpc3954 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[21]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[9],stage4_8[11],stage4_7[14]}
   );
   gpc615_5 gpc3955 (
      {stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36], stage3_7[37]},
      {stage3_8[22]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[10],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc3956 (
      {stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41], stage3_7[42]},
      {stage3_8[23]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[11],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc3957 (
      {stage3_7[43], stage3_7[44], stage3_7[45], stage3_7[46], stage3_7[47]},
      {stage3_8[24]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[12],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc3958 (
      {stage3_7[48], stage3_7[49], stage3_7[50], stage3_7[51], stage3_7[52]},
      {stage3_8[25]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[8],stage4_9[13],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc3959 (
      {stage3_7[53], stage3_7[54], stage3_7[55], stage3_7[56], stage3_7[57]},
      {stage3_8[26]},
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage4_11[6],stage4_10[9],stage4_9[14],stage4_8[16],stage4_7[19]}
   );
   gpc615_5 gpc3960 (
      {stage3_7[58], stage3_7[59], stage3_7[60], stage3_7[61], stage3_7[62]},
      {stage3_8[27]},
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage4_11[7],stage4_10[10],stage4_9[15],stage4_8[17],stage4_7[20]}
   );
   gpc606_5 gpc3961 (
      {stage3_8[28], stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[8],stage4_10[11],stage4_9[16],stage4_8[18]}
   );
   gpc623_5 gpc3962 (
      {stage3_9[48], stage3_9[49], stage3_9[50]},
      {stage3_10[6], stage3_10[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[9],stage4_10[12],stage4_9[17]}
   );
   gpc623_5 gpc3963 (
      {stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_10[8], stage3_10[9]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[2],stage4_11[10],stage4_10[13],stage4_9[18]}
   );
   gpc623_5 gpc3964 (
      {stage3_9[54], stage3_9[55], stage3_9[56]},
      {stage3_10[10], stage3_10[11]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[3],stage4_11[11],stage4_10[14],stage4_9[19]}
   );
   gpc623_5 gpc3965 (
      {stage3_9[57], stage3_9[58], stage3_9[59]},
      {stage3_10[12], stage3_10[13]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[4],stage4_11[12],stage4_10[15],stage4_9[20]}
   );
   gpc623_5 gpc3966 (
      {stage3_9[60], stage3_9[61], stage3_9[62]},
      {stage3_10[14], stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[5],stage4_11[13],stage4_10[16],stage4_9[21]}
   );
   gpc623_5 gpc3967 (
      {stage3_9[63], stage3_9[64], stage3_9[65]},
      {stage3_10[16], stage3_10[17]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[6],stage4_11[14],stage4_10[17],stage4_9[22]}
   );
   gpc1163_5 gpc3968 (
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[6],stage4_12[7],stage4_11[15]}
   );
   gpc606_5 gpc3969 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[7],stage4_12[8]}
   );
   gpc606_5 gpc3970 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage4_16[1],stage4_15[2],stage4_14[2],stage4_13[8],stage4_12[9]}
   );
   gpc606_5 gpc3971 (
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18]},
      {stage4_16[2],stage4_15[3],stage4_14[3],stage4_13[9],stage4_12[10]}
   );
   gpc606_5 gpc3972 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage4_16[3],stage4_15[4],stage4_14[4],stage4_13[10],stage4_12[11]}
   );
   gpc606_5 gpc3973 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage4_16[4],stage4_15[5],stage4_14[5],stage4_13[11],stage4_12[12]}
   );
   gpc606_5 gpc3974 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], stage3_14[36]},
      {stage4_16[5],stage4_15[6],stage4_14[6],stage4_13[12],stage4_12[13]}
   );
   gpc2135_5 gpc3975 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[37], stage3_14[38], stage3_14[39]},
      {stage3_15[0]},
      {stage3_16[0], stage3_16[1]},
      {stage4_17[0],stage4_16[6],stage4_15[7],stage4_14[7],stage4_13[13]}
   );
   gpc2135_5 gpc3976 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[40], stage3_14[41], stage3_14[42]},
      {stage3_15[1]},
      {stage3_16[2], stage3_16[3]},
      {stage4_17[1],stage4_16[7],stage4_15[8],stage4_14[8],stage4_13[14]}
   );
   gpc2135_5 gpc3977 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[43], stage3_14[44], stage3_14[45]},
      {stage3_15[2]},
      {stage3_16[4], stage3_16[5]},
      {stage4_17[2],stage4_16[8],stage4_15[9],stage4_14[9],stage4_13[15]}
   );
   gpc2135_5 gpc3978 (
      {stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_14[46], stage3_14[47], stage3_14[48]},
      {stage3_15[3]},
      {stage3_16[6], stage3_16[7]},
      {stage4_17[3],stage4_16[9],stage4_15[10],stage4_14[10],stage4_13[16]}
   );
   gpc2135_5 gpc3979 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_14[49], stage3_14[50], 1'b0},
      {stage3_15[4]},
      {stage3_16[8], stage3_16[9]},
      {stage4_17[4],stage4_16[10],stage4_15[11],stage4_14[11],stage4_13[17]}
   );
   gpc606_5 gpc3980 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10]},
      {stage4_17[5],stage4_16[11],stage4_15[12],stage4_14[12],stage4_13[18]}
   );
   gpc2135_5 gpc3981 (
      {stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage3_16[10], stage3_16[11], stage3_16[12]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[6],stage4_16[12],stage4_15[13]}
   );
   gpc2135_5 gpc3982 (
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage3_17[1]},
      {stage3_18[2], stage3_18[3]},
      {stage4_19[1],stage4_18[1],stage4_17[7],stage4_16[13],stage4_15[14]}
   );
   gpc2135_5 gpc3983 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[2]},
      {stage3_18[4], stage3_18[5]},
      {stage4_19[2],stage4_18[2],stage4_17[8],stage4_16[14],stage4_15[15]}
   );
   gpc2135_5 gpc3984 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[19], stage3_16[20], stage3_16[21]},
      {stage3_17[3]},
      {stage3_18[6], stage3_18[7]},
      {stage4_19[3],stage4_18[3],stage4_17[9],stage4_16[15],stage4_15[16]}
   );
   gpc2135_5 gpc3985 (
      {stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage3_16[22], stage3_16[23], stage3_16[24]},
      {stage3_17[4]},
      {stage3_18[8], stage3_18[9]},
      {stage4_19[4],stage4_18[4],stage4_17[10],stage4_16[16],stage4_15[17]}
   );
   gpc2135_5 gpc3986 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40]},
      {stage3_16[25], stage3_16[26], stage3_16[27]},
      {stage3_17[5]},
      {stage3_18[10], stage3_18[11]},
      {stage4_19[5],stage4_18[5],stage4_17[11],stage4_16[17],stage4_15[18]}
   );
   gpc2135_5 gpc3987 (
      {stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45]},
      {stage3_16[28], stage3_16[29], stage3_16[30]},
      {stage3_17[6]},
      {stage3_18[12], stage3_18[13]},
      {stage4_19[6],stage4_18[6],stage4_17[12],stage4_16[18],stage4_15[19]}
   );
   gpc2135_5 gpc3988 (
      {stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49], stage3_15[50]},
      {stage3_16[31], stage3_16[32], stage3_16[33]},
      {stage3_17[7]},
      {stage3_18[14], stage3_18[15]},
      {stage4_19[7],stage4_18[7],stage4_17[13],stage4_16[19],stage4_15[20]}
   );
   gpc2135_5 gpc3989 (
      {stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54], stage3_15[55]},
      {stage3_16[34], stage3_16[35], stage3_16[36]},
      {stage3_17[8]},
      {stage3_18[16], stage3_18[17]},
      {stage4_19[8],stage4_18[8],stage4_17[14],stage4_16[20],stage4_15[21]}
   );
   gpc2135_5 gpc3990 (
      {stage3_15[56], stage3_15[57], stage3_15[58], stage3_15[59], stage3_15[60]},
      {stage3_16[37], stage3_16[38], stage3_16[39]},
      {stage3_17[9]},
      {stage3_18[18], stage3_18[19]},
      {stage4_19[9],stage4_18[9],stage4_17[15],stage4_16[21],stage4_15[22]}
   );
   gpc615_5 gpc3991 (
      {stage3_15[61], stage3_15[62], stage3_15[63], stage3_15[64], stage3_15[65]},
      {stage3_16[40]},
      {stage3_17[10], stage3_17[11], stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15]},
      {stage4_19[10],stage4_18[10],stage4_17[16],stage4_16[22],stage4_15[23]}
   );
   gpc606_5 gpc3992 (
      {stage3_16[41], stage3_16[42], stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46]},
      {stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage4_20[0],stage4_19[11],stage4_18[11],stage4_17[17],stage4_16[23]}
   );
   gpc606_5 gpc3993 (
      {stage3_16[47], stage3_16[48], stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52]},
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31]},
      {stage4_20[1],stage4_19[12],stage4_18[12],stage4_17[18],stage4_16[24]}
   );
   gpc606_5 gpc3994 (
      {stage3_16[53], stage3_16[54], stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58]},
      {stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35], stage3_18[36], stage3_18[37]},
      {stage4_20[2],stage4_19[13],stage4_18[13],stage4_17[19],stage4_16[25]}
   );
   gpc1163_5 gpc3995 (
      {stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41], stage3_18[42], stage3_18[43]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[3],stage4_19[14],stage4_18[14],stage4_17[20]}
   );
   gpc1163_5 gpc3996 (
      {stage3_17[19], stage3_17[20], stage3_17[21]},
      {stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48], stage3_18[49]},
      {stage3_19[1]},
      {stage3_20[1]},
      {stage4_21[1],stage4_20[4],stage4_19[15],stage4_18[15],stage4_17[21]}
   );
   gpc606_5 gpc3997 (
      {stage3_17[22], stage3_17[23], stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27]},
      {stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6], stage3_19[7]},
      {stage4_21[2],stage4_20[5],stage4_19[16],stage4_18[16],stage4_17[22]}
   );
   gpc606_5 gpc3998 (
      {stage3_17[28], stage3_17[29], stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33]},
      {stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11], stage3_19[12], stage3_19[13]},
      {stage4_21[3],stage4_20[6],stage4_19[17],stage4_18[17],stage4_17[23]}
   );
   gpc606_5 gpc3999 (
      {stage3_17[34], stage3_17[35], stage3_17[36], stage3_17[37], stage3_17[38], stage3_17[39]},
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage4_21[4],stage4_20[7],stage4_19[18],stage4_18[18],stage4_17[24]}
   );
   gpc615_5 gpc4000 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24]},
      {stage3_20[2]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[5],stage4_20[8],stage4_19[19]}
   );
   gpc615_5 gpc4001 (
      {stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage3_20[3]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[6],stage4_20[9],stage4_19[20]}
   );
   gpc615_5 gpc4002 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[4]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[7],stage4_20[10],stage4_19[21]}
   );
   gpc615_5 gpc4003 (
      {stage3_19[35], stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39]},
      {stage3_20[5]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[8],stage4_20[11],stage4_19[22]}
   );
   gpc1325_5 gpc4004 (
      {stage3_19[40], stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44]},
      {stage3_20[6], stage3_20[7]},
      {stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_22[0]},
      {stage4_23[4],stage4_22[4],stage4_21[9],stage4_20[12],stage4_19[23]}
   );
   gpc1406_5 gpc4005 (
      {stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4]},
      {stage3_23[0]},
      {stage4_24[0],stage4_23[5],stage4_22[5],stage4_21[10],stage4_20[13]}
   );
   gpc606_5 gpc4006 (
      {stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19]},
      {stage3_22[5], stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage4_24[1],stage4_23[6],stage4_22[6],stage4_21[11],stage4_20[14]}
   );
   gpc606_5 gpc4007 (
      {stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24], stage3_20[25]},
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage4_24[2],stage4_23[7],stage4_22[7],stage4_21[12],stage4_20[15]}
   );
   gpc606_5 gpc4008 (
      {stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31]},
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22]},
      {stage4_24[3],stage4_23[8],stage4_22[8],stage4_21[13],stage4_20[16]}
   );
   gpc606_5 gpc4009 (
      {stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37]},
      {stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28]},
      {stage4_24[4],stage4_23[9],stage4_22[9],stage4_21[14],stage4_20[17]}
   );
   gpc606_5 gpc4010 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage4_25[0],stage4_24[5],stage4_23[10],stage4_22[10],stage4_21[15]}
   );
   gpc606_5 gpc4011 (
      {stage3_21[33], stage3_21[34], stage3_21[35], stage3_21[36], stage3_21[37], stage3_21[38]},
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12]},
      {stage4_25[1],stage4_24[6],stage4_23[11],stage4_22[11],stage4_21[16]}
   );
   gpc606_5 gpc4012 (
      {stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42], stage3_21[43], stage3_21[44]},
      {stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage4_25[2],stage4_24[7],stage4_23[12],stage4_22[12],stage4_21[17]}
   );
   gpc606_5 gpc4013 (
      {stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23], stage3_23[24]},
      {stage4_25[3],stage4_24[8],stage4_23[13],stage4_22[13],stage4_21[18]}
   );
   gpc606_5 gpc4014 (
      {stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54], stage3_21[55], stage3_21[56]},
      {stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28], stage3_23[29], stage3_23[30]},
      {stage4_25[4],stage4_24[9],stage4_23[14],stage4_22[14],stage4_21[19]}
   );
   gpc606_5 gpc4015 (
      {stage3_22[29], stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[5],stage4_24[10],stage4_23[15],stage4_22[15]}
   );
   gpc606_5 gpc4016 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[6],stage4_24[11],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc4017 (
      {stage3_23[31], stage3_23[32], stage3_23[33], stage3_23[34], stage3_23[35]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[7],stage4_24[12],stage4_23[17]}
   );
   gpc615_5 gpc4018 (
      {stage3_23[36], stage3_23[37], stage3_23[38], stage3_23[39], stage3_23[40]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[8],stage4_24[13],stage4_23[18]}
   );
   gpc615_5 gpc4019 (
      {stage3_23[41], stage3_23[42], stage3_23[43], stage3_23[44], stage3_23[45]},
      {stage3_24[14]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[9],stage4_24[14],stage4_23[19]}
   );
   gpc606_5 gpc4020 (
      {stage3_24[15], stage3_24[16], stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[3],stage4_26[5],stage4_25[10],stage4_24[15]}
   );
   gpc606_5 gpc4021 (
      {stage3_24[21], stage3_24[22], stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[4],stage4_26[6],stage4_25[11],stage4_24[16]}
   );
   gpc606_5 gpc4022 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[2],stage4_27[5],stage4_26[7],stage4_25[12]}
   );
   gpc615_5 gpc4023 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28]},
      {stage3_26[12]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[3],stage4_27[6],stage4_26[8],stage4_25[13]}
   );
   gpc615_5 gpc4024 (
      {stage3_25[29], stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33]},
      {stage3_26[13]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[4],stage4_27[7],stage4_26[9],stage4_25[14]}
   );
   gpc615_5 gpc4025 (
      {stage3_25[34], stage3_25[35], stage3_25[36], stage3_25[37], stage3_25[38]},
      {stage3_26[14]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[5],stage4_27[8],stage4_26[10],stage4_25[15]}
   );
   gpc615_5 gpc4026 (
      {stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18], stage3_26[19]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[6],stage4_27[9],stage4_26[11]}
   );
   gpc606_5 gpc4027 (
      {stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[1],stage4_29[5],stage4_28[7],stage4_27[10]}
   );
   gpc606_5 gpc4028 (
      {stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[2],stage4_29[6],stage4_28[8],stage4_27[11]}
   );
   gpc606_5 gpc4029 (
      {stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[3],stage4_29[7],stage4_28[9],stage4_27[12]}
   );
   gpc606_5 gpc4030 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47], stage3_27[48]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[4],stage4_29[8],stage4_28[10],stage4_27[13]}
   );
   gpc615_5 gpc4031 (
      {stage3_27[49], stage3_27[50], stage3_27[51], stage3_27[52], stage3_27[53]},
      {stage3_28[6]},
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage4_31[4],stage4_30[5],stage4_29[9],stage4_28[11],stage4_27[14]}
   );
   gpc606_5 gpc4032 (
      {stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[5],stage4_30[6],stage4_29[10],stage4_28[12]}
   );
   gpc606_5 gpc4033 (
      {stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[6],stage4_30[7],stage4_29[11],stage4_28[13]}
   );
   gpc606_5 gpc4034 (
      {stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[7],stage4_30[8],stage4_29[12],stage4_28[14]}
   );
   gpc606_5 gpc4035 (
      {stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[8],stage4_30[9],stage4_29[13],stage4_28[15]}
   );
   gpc606_5 gpc4036 (
      {stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[9],stage4_30[10],stage4_29[14],stage4_28[16]}
   );
   gpc606_5 gpc4037 (
      {stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[10],stage4_30[11],stage4_29[15],stage4_28[17]}
   );
   gpc615_5 gpc4038 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34]},
      {stage3_30[36]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[6],stage4_31[11],stage4_30[12],stage4_29[16]}
   );
   gpc606_5 gpc4039 (
      {stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41], stage3_30[42]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[7],stage4_31[12],stage4_30[13]}
   );
   gpc615_5 gpc4040 (
      {stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage3_31[6]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[2],stage4_32[8],stage4_31[13],stage4_30[14]}
   );
   gpc615_5 gpc4041 (
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52]},
      {stage3_31[7]},
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage4_34[2],stage4_33[3],stage4_32[9],stage4_31[14],stage4_30[15]}
   );
   gpc606_5 gpc4042 (
      {stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[3],stage4_33[4],stage4_32[10],stage4_31[15]}
   );
   gpc606_5 gpc4043 (
      {stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[4],stage4_33[5],stage4_32[11],stage4_31[16]}
   );
   gpc615_5 gpc4044 (
      {stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23], stage3_31[24]},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[5],stage4_33[6],stage4_32[12],stage4_31[17]}
   );
   gpc615_5 gpc4045 (
      {stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage3_32[19]},
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage4_35[3],stage4_34[6],stage4_33[7],stage4_32[13],stage4_31[18]}
   );
   gpc615_5 gpc4046 (
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34]},
      {stage3_32[20]},
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29]},
      {stage4_35[4],stage4_34[7],stage4_33[8],stage4_32[14],stage4_31[19]}
   );
   gpc1325_5 gpc4047 (
      {stage3_31[35], stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39]},
      {stage3_32[21], stage3_32[22]},
      {stage3_33[30], stage3_33[31], stage3_33[32]},
      {stage3_34[0]},
      {stage4_35[5],stage4_34[8],stage4_33[9],stage4_32[15],stage4_31[20]}
   );
   gpc606_5 gpc4048 (
      {stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28]},
      {stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6]},
      {stage4_36[0],stage4_35[6],stage4_34[9],stage4_33[10],stage4_32[16]}
   );
   gpc606_5 gpc4049 (
      {stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34]},
      {stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12]},
      {stage4_36[1],stage4_35[7],stage4_34[10],stage4_33[11],stage4_32[17]}
   );
   gpc606_5 gpc4050 (
      {stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[8],stage4_34[11],stage4_33[12]}
   );
   gpc2135_5 gpc4051 (
      {stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage3_35[6], stage3_35[7], stage3_35[8]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1]},
      {stage4_38[0],stage4_37[1],stage4_36[3],stage4_35[9],stage4_34[12]}
   );
   gpc1_1 gpc4052 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4053 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4054 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4055 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4056 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4057 (
      {stage3_1[15]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4058 (
      {stage3_1[16]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4059 (
      {stage3_1[17]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4060 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4061 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4062 (
      {stage3_4[39]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4063 (
      {stage3_4[40]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4064 (
      {stage3_4[41]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4065 (
      {stage3_4[42]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4066 (
      {stage3_4[43]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4067 (
      {stage3_5[42]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4068 (
      {stage3_5[43]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4069 (
      {stage3_5[44]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4070 (
      {stage3_5[45]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4071 (
      {stage3_5[46]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4072 (
      {stage3_5[47]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4073 (
      {stage3_5[48]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4074 (
      {stage3_6[39]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4075 (
      {stage3_6[40]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4076 (
      {stage3_6[41]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4077 (
      {stage3_6[42]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4078 (
      {stage3_7[63]},
      {stage4_7[21]}
   );
   gpc1_1 gpc4079 (
      {stage3_7[64]},
      {stage4_7[22]}
   );
   gpc1_1 gpc4080 (
      {stage3_7[65]},
      {stage4_7[23]}
   );
   gpc1_1 gpc4081 (
      {stage3_7[66]},
      {stage4_7[24]}
   );
   gpc1_1 gpc4082 (
      {stage3_7[67]},
      {stage4_7[25]}
   );
   gpc1_1 gpc4083 (
      {stage3_7[68]},
      {stage4_7[26]}
   );
   gpc1_1 gpc4084 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc4085 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc4086 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4087 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4088 (
      {stage3_9[66]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4089 (
      {stage3_9[67]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4090 (
      {stage3_9[68]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4091 (
      {stage3_9[69]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4092 (
      {stage3_10[18]},
      {stage4_10[18]}
   );
   gpc1_1 gpc4093 (
      {stage3_10[19]},
      {stage4_10[19]}
   );
   gpc1_1 gpc4094 (
      {stage3_10[20]},
      {stage4_10[20]}
   );
   gpc1_1 gpc4095 (
      {stage3_10[21]},
      {stage4_10[21]}
   );
   gpc1_1 gpc4096 (
      {stage3_10[22]},
      {stage4_10[22]}
   );
   gpc1_1 gpc4097 (
      {stage3_10[23]},
      {stage4_10[23]}
   );
   gpc1_1 gpc4098 (
      {stage3_10[24]},
      {stage4_10[24]}
   );
   gpc1_1 gpc4099 (
      {stage3_10[25]},
      {stage4_10[25]}
   );
   gpc1_1 gpc4100 (
      {stage3_10[26]},
      {stage4_10[26]}
   );
   gpc1_1 gpc4101 (
      {stage3_10[27]},
      {stage4_10[27]}
   );
   gpc1_1 gpc4102 (
      {stage3_10[28]},
      {stage4_10[28]}
   );
   gpc1_1 gpc4103 (
      {stage3_11[39]},
      {stage4_11[16]}
   );
   gpc1_1 gpc4104 (
      {stage3_11[40]},
      {stage4_11[17]}
   );
   gpc1_1 gpc4105 (
      {stage3_11[41]},
      {stage4_11[18]}
   );
   gpc1_1 gpc4106 (
      {stage3_11[42]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4107 (
      {stage3_11[43]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4108 (
      {stage3_13[32]},
      {stage4_13[19]}
   );
   gpc1_1 gpc4109 (
      {stage3_13[33]},
      {stage4_13[20]}
   );
   gpc1_1 gpc4110 (
      {stage3_13[34]},
      {stage4_13[21]}
   );
   gpc1_1 gpc4111 (
      {stage3_13[35]},
      {stage4_13[22]}
   );
   gpc1_1 gpc4112 (
      {stage3_13[36]},
      {stage4_13[23]}
   );
   gpc1_1 gpc4113 (
      {stage3_13[37]},
      {stage4_13[24]}
   );
   gpc1_1 gpc4114 (
      {stage3_13[38]},
      {stage4_13[25]}
   );
   gpc1_1 gpc4115 (
      {stage3_13[39]},
      {stage4_13[26]}
   );
   gpc1_1 gpc4116 (
      {stage3_13[40]},
      {stage4_13[27]}
   );
   gpc1_1 gpc4117 (
      {stage3_15[66]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4118 (
      {stage3_15[67]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4119 (
      {stage3_15[68]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4120 (
      {stage3_15[69]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4121 (
      {stage3_15[70]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4122 (
      {stage3_15[71]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4123 (
      {stage3_15[72]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4124 (
      {stage3_15[73]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4125 (
      {stage3_15[74]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4126 (
      {stage3_15[75]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4127 (
      {stage3_15[76]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4128 (
      {stage3_15[77]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4129 (
      {stage3_15[78]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4130 (
      {stage3_15[79]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4131 (
      {stage3_15[80]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4132 (
      {stage3_15[81]},
      {stage4_15[39]}
   );
   gpc1_1 gpc4133 (
      {stage3_15[82]},
      {stage4_15[40]}
   );
   gpc1_1 gpc4134 (
      {stage3_15[83]},
      {stage4_15[41]}
   );
   gpc1_1 gpc4135 (
      {stage3_15[84]},
      {stage4_15[42]}
   );
   gpc1_1 gpc4136 (
      {stage3_15[85]},
      {stage4_15[43]}
   );
   gpc1_1 gpc4137 (
      {stage3_15[86]},
      {stage4_15[44]}
   );
   gpc1_1 gpc4138 (
      {stage3_15[87]},
      {stage4_15[45]}
   );
   gpc1_1 gpc4139 (
      {stage3_15[88]},
      {stage4_15[46]}
   );
   gpc1_1 gpc4140 (
      {stage3_15[89]},
      {stage4_15[47]}
   );
   gpc1_1 gpc4141 (
      {stage3_16[59]},
      {stage4_16[26]}
   );
   gpc1_1 gpc4142 (
      {stage3_16[60]},
      {stage4_16[27]}
   );
   gpc1_1 gpc4143 (
      {stage3_16[61]},
      {stage4_16[28]}
   );
   gpc1_1 gpc4144 (
      {stage3_17[40]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4145 (
      {stage3_17[41]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4146 (
      {stage3_17[42]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4147 (
      {stage3_17[43]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4148 (
      {stage3_17[44]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4149 (
      {stage3_17[45]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4150 (
      {stage3_17[46]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4151 (
      {stage3_17[47]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4152 (
      {stage3_17[48]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4153 (
      {stage3_17[49]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4154 (
      {stage3_19[45]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4155 (
      {stage3_19[46]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4156 (
      {stage3_19[47]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4157 (
      {stage3_19[48]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4158 (
      {stage3_19[49]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4159 (
      {stage3_20[38]},
      {stage4_20[18]}
   );
   gpc1_1 gpc4160 (
      {stage3_20[39]},
      {stage4_20[19]}
   );
   gpc1_1 gpc4161 (
      {stage3_20[40]},
      {stage4_20[20]}
   );
   gpc1_1 gpc4162 (
      {stage3_20[41]},
      {stage4_20[21]}
   );
   gpc1_1 gpc4163 (
      {stage3_20[42]},
      {stage4_20[22]}
   );
   gpc1_1 gpc4164 (
      {stage3_20[43]},
      {stage4_20[23]}
   );
   gpc1_1 gpc4165 (
      {stage3_20[44]},
      {stage4_20[24]}
   );
   gpc1_1 gpc4166 (
      {stage3_20[45]},
      {stage4_20[25]}
   );
   gpc1_1 gpc4167 (
      {stage3_21[57]},
      {stage4_21[20]}
   );
   gpc1_1 gpc4168 (
      {stage3_21[58]},
      {stage4_21[21]}
   );
   gpc1_1 gpc4169 (
      {stage3_22[41]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4170 (
      {stage3_22[42]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4171 (
      {stage3_22[43]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4172 (
      {stage3_22[44]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4173 (
      {stage3_22[45]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4174 (
      {stage3_22[46]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4175 (
      {stage3_23[46]},
      {stage4_23[20]}
   );
   gpc1_1 gpc4176 (
      {stage3_23[47]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4177 (
      {stage3_24[27]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4178 (
      {stage3_24[28]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4179 (
      {stage3_24[29]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4180 (
      {stage3_24[30]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4181 (
      {stage3_24[31]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4182 (
      {stage3_24[32]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4183 (
      {stage3_24[33]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4184 (
      {stage3_24[34]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4185 (
      {stage3_24[35]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4186 (
      {stage3_24[36]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4187 (
      {stage3_24[37]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4188 (
      {stage3_24[38]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4189 (
      {stage3_24[39]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4190 (
      {stage3_24[40]},
      {stage4_24[30]}
   );
   gpc1_1 gpc4191 (
      {stage3_25[39]},
      {stage4_25[16]}
   );
   gpc1_1 gpc4192 (
      {stage3_26[20]},
      {stage4_26[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_26[21]},
      {stage4_26[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_26[24]},
      {stage4_26[16]}
   );
   gpc1_1 gpc4197 (
      {stage3_26[25]},
      {stage4_26[17]}
   );
   gpc1_1 gpc4198 (
      {stage3_26[26]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4199 (
      {stage3_26[27]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4200 (
      {stage3_26[28]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4201 (
      {stage3_26[29]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4202 (
      {stage3_26[30]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4203 (
      {stage3_26[31]},
      {stage4_26[23]}
   );
   gpc1_1 gpc4204 (
      {stage3_27[54]},
      {stage4_27[15]}
   );
   gpc1_1 gpc4205 (
      {stage3_27[55]},
      {stage4_27[16]}
   );
   gpc1_1 gpc4206 (
      {stage3_27[56]},
      {stage4_27[17]}
   );
   gpc1_1 gpc4207 (
      {stage3_27[57]},
      {stage4_27[18]}
   );
   gpc1_1 gpc4208 (
      {stage3_27[58]},
      {stage4_27[19]}
   );
   gpc1_1 gpc4209 (
      {stage3_27[59]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4210 (
      {stage3_27[60]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4211 (
      {stage3_27[61]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4212 (
      {stage3_27[62]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4213 (
      {stage3_27[63]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4214 (
      {stage3_27[64]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4215 (
      {stage3_27[65]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4216 (
      {stage3_27[66]},
      {stage4_27[27]}
   );
   gpc1_1 gpc4217 (
      {stage3_29[35]},
      {stage4_29[17]}
   );
   gpc1_1 gpc4218 (
      {stage3_29[36]},
      {stage4_29[18]}
   );
   gpc1_1 gpc4219 (
      {stage3_29[37]},
      {stage4_29[19]}
   );
   gpc1_1 gpc4220 (
      {stage3_29[38]},
      {stage4_29[20]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[53]},
      {stage4_30[16]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[54]},
      {stage4_30[17]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[55]},
      {stage4_30[18]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[56]},
      {stage4_30[19]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[57]},
      {stage4_30[20]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[58]},
      {stage4_30[21]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[59]},
      {stage4_30[22]}
   );
   gpc1_1 gpc4228 (
      {stage3_32[35]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4229 (
      {stage3_33[39]},
      {stage4_33[13]}
   );
   gpc1_1 gpc4230 (
      {stage3_34[18]},
      {stage4_34[13]}
   );
   gpc1_1 gpc4231 (
      {stage3_34[19]},
      {stage4_34[14]}
   );
   gpc1_1 gpc4232 (
      {stage3_34[20]},
      {stage4_34[15]}
   );
   gpc1_1 gpc4233 (
      {stage3_34[21]},
      {stage4_34[16]}
   );
   gpc1_1 gpc4234 (
      {stage3_35[9]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4235 (
      {stage3_35[10]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4236 (
      {stage3_35[11]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4237 (
      {stage3_35[12]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4238 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc4239 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4240 (
      {stage3_36[3]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4241 (
      {stage3_36[4]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4242 (
      {stage3_36[5]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4243 (
      {stage3_36[6]},
      {stage4_36[9]}
   );
   gpc615_5 gpc4244 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc1343_5 gpc4245 (
      {stage4_3[1], stage4_3[2], stage4_3[3]},
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc606_5 gpc4246 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc1415_5 gpc4247 (
      {stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_6[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc606_5 gpc4248 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9]},
      {stage5_9[1],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc4249 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15]},
      {stage5_9[2],stage5_8[3],stage5_7[4],stage5_6[5],stage5_5[5]}
   );
   gpc606_5 gpc4250 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13]},
      {stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[5],stage5_6[6]}
   );
   gpc615_5 gpc4251 (
      {stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage4_7[16]},
      {stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage5_10[1],stage5_9[4],stage5_8[5],stage5_7[6],stage5_6[7]}
   );
   gpc1343_5 gpc4252 (
      {stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[5],stage5_8[6],stage5_7[7]}
   );
   gpc615_5 gpc4253 (
      {stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage4_8[17]},
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8]},
      {stage5_11[1],stage5_10[3],stage5_9[6],stage5_8[7],stage5_7[8]}
   );
   gpc606_5 gpc4254 (
      {stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[7]}
   );
   gpc615_5 gpc4255 (
      {stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18], stage4_9[19]},
      {stage4_10[1]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[8]}
   );
   gpc615_5 gpc4256 (
      {stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_10[2]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[9]}
   );
   gpc207_4 gpc4257 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc615_5 gpc4258 (
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14]},
      {stage4_11[18]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[4],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc1163_5 gpc4259 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[5]}
   );
   gpc606_5 gpc4260 (
      {stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[6]}
   );
   gpc606_5 gpc4261 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12]},
      {stage5_17[2],stage5_16[2],stage5_15[2],stage5_14[3],stage5_13[7]}
   );
   gpc606_5 gpc4262 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19], stage4_13[20]},
      {stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage5_17[3],stage5_16[3],stage5_15[3],stage5_14[4],stage5_13[8]}
   );
   gpc615_5 gpc4263 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[19]},
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage5_18[0],stage5_17[4],stage5_16[4],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc4264 (
      {stage4_15[20], stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26]},
      {stage4_17[0], stage4_17[1]},
      {stage5_18[1],stage5_17[5],stage5_16[5],stage5_15[5]}
   );
   gpc615_5 gpc4265 (
      {stage4_15[27], stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31]},
      {stage4_16[7]},
      {stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6], stage4_17[7]},
      {stage5_19[0],stage5_18[2],stage5_17[6],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc4266 (
      {stage4_15[32], stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36]},
      {stage4_16[8]},
      {stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12], stage4_17[13]},
      {stage5_19[1],stage5_18[3],stage5_17[7],stage5_16[7],stage5_15[7]}
   );
   gpc615_5 gpc4267 (
      {stage4_15[37], stage4_15[38], stage4_15[39], stage4_15[40], stage4_15[41]},
      {stage4_16[9]},
      {stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17], stage4_17[18], stage4_17[19]},
      {stage5_19[2],stage5_18[4],stage5_17[8],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4268 (
      {stage4_15[42], stage4_15[43], stage4_15[44], stage4_15[45], stage4_15[46]},
      {stage4_16[10]},
      {stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23], stage4_17[24], stage4_17[25]},
      {stage5_19[3],stage5_18[5],stage5_17[9],stage5_16[9],stage5_15[9]}
   );
   gpc207_4 gpc4269 (
      {stage4_16[11], stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[4],stage5_18[6],stage5_17[10],stage5_16[10]}
   );
   gpc606_5 gpc4270 (
      {stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30], stage4_17[31]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[5],stage5_18[7],stage5_17[11]}
   );
   gpc615_5 gpc4271 (
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[6],stage5_18[8]}
   );
   gpc615_5 gpc4272 (
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[7],stage5_18[9]}
   );
   gpc615_5 gpc4273 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16]},
      {stage4_19[8]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[8],stage5_18[10]}
   );
   gpc2135_5 gpc4274 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage4_21[0]},
      {stage4_22[0], stage4_22[1]},
      {stage5_23[0],stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[9]}
   );
   gpc615_5 gpc4275 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[21]},
      {stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[10]}
   );
   gpc615_5 gpc4276 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[22]},
      {stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11], stage4_21[12]},
      {stage5_23[2],stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[11]}
   );
   gpc615_5 gpc4277 (
      {stage4_19[24], stage4_19[25], stage4_19[26], stage4_19[27], stage4_19[28]},
      {stage4_20[23]},
      {stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[3],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[12]}
   );
   gpc615_5 gpc4278 (
      {stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[7]}
   );
   gpc615_5 gpc4279 (
      {stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage4_23[1]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[8]}
   );
   gpc615_5 gpc4280 (
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16]},
      {stage4_23[2]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[9]}
   );
   gpc615_5 gpc4281 (
      {stage4_22[17], stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21]},
      {stage4_23[3]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[10]}
   );
   gpc615_5 gpc4282 (
      {stage4_23[4], stage4_23[5], stage4_23[6], stage4_23[7], stage4_23[8]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[8]}
   );
   gpc615_5 gpc4283 (
      {stage4_23[9], stage4_23[10], stage4_23[11], stage4_23[12], stage4_23[13]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[9]}
   );
   gpc615_5 gpc4284 (
      {stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17], stage4_23[18]},
      {stage4_24[26]},
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], 1'b0},
      {stage5_27[2],stage5_26[6],stage5_25[6],stage5_24[6],stage5_23[10]}
   );
   gpc606_5 gpc4285 (
      {stage4_24[27], stage4_24[28], stage4_24[29], stage4_24[30], 1'b0, 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[3],stage5_26[7],stage5_25[7],stage5_24[7]}
   );
   gpc615_5 gpc4286 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4287 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4288 (
      {stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19], stage4_26[20]},
      {stage4_27[2]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[3],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4289 (
      {stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[3],stage5_29[3],stage5_28[4],stage5_27[7]}
   );
   gpc207_4 gpc4290 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[2], stage4_29[3]},
      {stage5_30[4],stage5_29[4],stage5_28[5],stage5_27[8]}
   );
   gpc207_4 gpc4291 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage4_29[4], stage4_29[5]},
      {stage5_30[5],stage5_29[5],stage5_28[6],stage5_27[9]}
   );
   gpc615_5 gpc4292 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[6],stage5_29[6]}
   );
   gpc615_5 gpc4293 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[7],stage5_29[7]}
   );
   gpc117_4 gpc4294 (
      {stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7], stage4_30[8]},
      {stage4_31[12]},
      {stage4_32[0]},
      {stage5_33[2],stage5_32[2],stage5_31[2],stage5_30[8]}
   );
   gpc117_4 gpc4295 (
      {stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15]},
      {stage4_31[13]},
      {stage4_32[1]},
      {stage5_33[3],stage5_32[3],stage5_31[3],stage5_30[9]}
   );
   gpc615_5 gpc4296 (
      {stage4_30[16], stage4_30[17], stage4_30[18], stage4_30[19], stage4_30[20]},
      {stage4_31[14]},
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage5_34[0],stage5_33[4],stage5_32[4],stage5_31[4],stage5_30[10]}
   );
   gpc615_5 gpc4297 (
      {stage4_30[21], stage4_30[22], 1'b0, 1'b0, 1'b0},
      {stage4_31[15]},
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage5_34[1],stage5_33[5],stage5_32[5],stage5_31[5],stage5_30[11]}
   );
   gpc2135_5 gpc4298 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4]},
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage4_35[0]},
      {stage4_36[0], stage4_36[1]},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[6]}
   );
   gpc2135_5 gpc4299 (
      {stage4_33[5], stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9]},
      {stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_35[1]},
      {stage4_36[2], stage4_36[3]},
      {stage5_37[1],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[7]}
   );
   gpc2135_5 gpc4300 (
      {stage4_33[10], stage4_33[11], stage4_33[12], stage4_33[13], 1'b0},
      {stage4_34[6], stage4_34[7], stage4_34[8]},
      {stage4_35[2]},
      {stage4_36[4], stage4_36[5]},
      {stage5_37[2],stage5_36[2],stage5_35[2],stage5_34[4],stage5_33[8]}
   );
   gpc606_5 gpc4301 (
      {stage4_34[9], stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], 1'b0, 1'b0},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[3],stage5_34[5]}
   );
   gpc1_1 gpc4302 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4303 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4304 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4305 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc4306 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4307 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4308 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4309 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4310 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4311 (
      {stage4_1[6]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4312 (
      {stage4_1[7]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4313 (
      {stage4_1[8]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4314 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4315 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4316 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4317 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4318 (
      {stage4_3[4]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4319 (
      {stage4_3[5]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4320 (
      {stage4_3[6]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4321 (
      {stage4_3[7]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4322 (
      {stage4_3[8]},
      {stage5_3[6]}
   );
   gpc1_1 gpc4323 (
      {stage4_3[9]},
      {stage5_3[7]}
   );
   gpc1_1 gpc4324 (
      {stage4_4[16]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4325 (
      {stage4_5[20]},
      {stage5_5[6]}
   );
   gpc1_1 gpc4326 (
      {stage4_5[21]},
      {stage5_5[7]}
   );
   gpc1_1 gpc4327 (
      {stage4_5[22]},
      {stage5_5[8]}
   );
   gpc1_1 gpc4328 (
      {stage4_6[19]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4329 (
      {stage4_6[20]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4330 (
      {stage4_7[25]},
      {stage5_7[9]}
   );
   gpc1_1 gpc4331 (
      {stage4_7[26]},
      {stage5_7[10]}
   );
   gpc1_1 gpc4332 (
      {stage4_8[18]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4333 (
      {stage4_8[19]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4334 (
      {stage4_8[20]},
      {stage5_8[10]}
   );
   gpc1_1 gpc4335 (
      {stage4_8[21]},
      {stage5_8[11]}
   );
   gpc1_1 gpc4336 (
      {stage4_8[22]},
      {stage5_8[12]}
   );
   gpc1_1 gpc4337 (
      {stage4_9[25]},
      {stage5_9[10]}
   );
   gpc1_1 gpc4338 (
      {stage4_9[26]},
      {stage5_9[11]}
   );
   gpc1_1 gpc4339 (
      {stage4_10[15]},
      {stage5_10[9]}
   );
   gpc1_1 gpc4340 (
      {stage4_10[16]},
      {stage5_10[10]}
   );
   gpc1_1 gpc4341 (
      {stage4_10[17]},
      {stage5_10[11]}
   );
   gpc1_1 gpc4342 (
      {stage4_10[18]},
      {stage5_10[12]}
   );
   gpc1_1 gpc4343 (
      {stage4_10[19]},
      {stage5_10[13]}
   );
   gpc1_1 gpc4344 (
      {stage4_10[20]},
      {stage5_10[14]}
   );
   gpc1_1 gpc4345 (
      {stage4_10[21]},
      {stage5_10[15]}
   );
   gpc1_1 gpc4346 (
      {stage4_10[22]},
      {stage5_10[16]}
   );
   gpc1_1 gpc4347 (
      {stage4_10[23]},
      {stage5_10[17]}
   );
   gpc1_1 gpc4348 (
      {stage4_10[24]},
      {stage5_10[18]}
   );
   gpc1_1 gpc4349 (
      {stage4_10[25]},
      {stage5_10[19]}
   );
   gpc1_1 gpc4350 (
      {stage4_10[26]},
      {stage5_10[20]}
   );
   gpc1_1 gpc4351 (
      {stage4_10[27]},
      {stage5_10[21]}
   );
   gpc1_1 gpc4352 (
      {stage4_10[28]},
      {stage5_10[22]}
   );
   gpc1_1 gpc4353 (
      {stage4_11[19]},
      {stage5_11[7]}
   );
   gpc1_1 gpc4354 (
      {stage4_11[20]},
      {stage5_11[8]}
   );
   gpc1_1 gpc4355 (
      {stage4_12[8]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4356 (
      {stage4_12[9]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4357 (
      {stage4_12[10]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4358 (
      {stage4_12[11]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4359 (
      {stage4_12[12]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4360 (
      {stage4_12[13]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4361 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc4362 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc4363 (
      {stage4_13[23]},
      {stage5_13[11]}
   );
   gpc1_1 gpc4364 (
      {stage4_13[24]},
      {stage5_13[12]}
   );
   gpc1_1 gpc4365 (
      {stage4_13[25]},
      {stage5_13[13]}
   );
   gpc1_1 gpc4366 (
      {stage4_13[26]},
      {stage5_13[14]}
   );
   gpc1_1 gpc4367 (
      {stage4_13[27]},
      {stage5_13[15]}
   );
   gpc1_1 gpc4368 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4369 (
      {stage4_14[12]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4370 (
      {stage4_15[47]},
      {stage5_15[10]}
   );
   gpc1_1 gpc4371 (
      {stage4_16[18]},
      {stage5_16[11]}
   );
   gpc1_1 gpc4372 (
      {stage4_16[19]},
      {stage5_16[12]}
   );
   gpc1_1 gpc4373 (
      {stage4_16[20]},
      {stage5_16[13]}
   );
   gpc1_1 gpc4374 (
      {stage4_16[21]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4375 (
      {stage4_16[22]},
      {stage5_16[15]}
   );
   gpc1_1 gpc4376 (
      {stage4_16[23]},
      {stage5_16[16]}
   );
   gpc1_1 gpc4377 (
      {stage4_16[24]},
      {stage5_16[17]}
   );
   gpc1_1 gpc4378 (
      {stage4_16[25]},
      {stage5_16[18]}
   );
   gpc1_1 gpc4379 (
      {stage4_16[26]},
      {stage5_16[19]}
   );
   gpc1_1 gpc4380 (
      {stage4_16[27]},
      {stage5_16[20]}
   );
   gpc1_1 gpc4381 (
      {stage4_16[28]},
      {stage5_16[21]}
   );
   gpc1_1 gpc4382 (
      {stage4_17[32]},
      {stage5_17[12]}
   );
   gpc1_1 gpc4383 (
      {stage4_17[33]},
      {stage5_17[13]}
   );
   gpc1_1 gpc4384 (
      {stage4_17[34]},
      {stage5_17[14]}
   );
   gpc1_1 gpc4385 (
      {stage4_18[17]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4386 (
      {stage4_18[18]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4387 (
      {stage4_20[24]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4388 (
      {stage4_20[25]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4389 (
      {stage4_21[19]},
      {stage5_21[8]}
   );
   gpc1_1 gpc4390 (
      {stage4_21[20]},
      {stage5_21[9]}
   );
   gpc1_1 gpc4391 (
      {stage4_21[21]},
      {stage5_21[10]}
   );
   gpc1_1 gpc4392 (
      {stage4_22[22]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4393 (
      {stage4_23[19]},
      {stage5_23[11]}
   );
   gpc1_1 gpc4394 (
      {stage4_23[20]},
      {stage5_23[12]}
   );
   gpc1_1 gpc4395 (
      {stage4_23[21]},
      {stage5_23[13]}
   );
   gpc1_1 gpc4396 (
      {stage4_26[21]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4397 (
      {stage4_26[22]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4398 (
      {stage4_26[23]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4399 (
      {stage4_27[24]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4400 (
      {stage4_27[25]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4401 (
      {stage4_27[26]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4402 (
      {stage4_27[27]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4403 (
      {stage4_29[16]},
      {stage5_29[8]}
   );
   gpc1_1 gpc4404 (
      {stage4_29[17]},
      {stage5_29[9]}
   );
   gpc1_1 gpc4405 (
      {stage4_29[18]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4406 (
      {stage4_29[19]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4407 (
      {stage4_29[20]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4408 (
      {stage4_31[16]},
      {stage5_31[6]}
   );
   gpc1_1 gpc4409 (
      {stage4_31[17]},
      {stage5_31[7]}
   );
   gpc1_1 gpc4410 (
      {stage4_31[18]},
      {stage5_31[8]}
   );
   gpc1_1 gpc4411 (
      {stage4_31[19]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4412 (
      {stage4_31[20]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4413 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4414 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4415 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4416 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4417 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4418 (
      {stage4_34[15]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4419 (
      {stage4_34[16]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4420 (
      {stage4_35[3]},
      {stage5_35[4]}
   );
   gpc1_1 gpc4421 (
      {stage4_35[4]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4422 (
      {stage4_35[5]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4423 (
      {stage4_35[6]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4424 (
      {stage4_35[7]},
      {stage5_35[8]}
   );
   gpc1_1 gpc4425 (
      {stage4_35[8]},
      {stage5_35[9]}
   );
   gpc1_1 gpc4426 (
      {stage4_35[9]},
      {stage5_35[10]}
   );
   gpc1_1 gpc4427 (
      {stage4_35[10]},
      {stage5_35[11]}
   );
   gpc1_1 gpc4428 (
      {stage4_35[11]},
      {stage5_35[12]}
   );
   gpc1_1 gpc4429 (
      {stage4_35[12]},
      {stage5_35[13]}
   );
   gpc1_1 gpc4430 (
      {stage4_35[13]},
      {stage5_35[14]}
   );
   gpc1_1 gpc4431 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4432 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4433 (
      {stage4_38[0]},
      {stage5_38[1]}
   );
   gpc1163_5 gpc4434 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], 1'b0},
      {stage5_3[0]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc135_4 gpc4435 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[1], stage5_4[2], stage5_4[3]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc1343_5 gpc4436 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[2]}
   );
   gpc1343_5 gpc4437 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[2],stage6_5[3]}
   );
   gpc615_5 gpc4438 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc4439 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[3],stage6_8[3]}
   );
   gpc606_5 gpc4440 (
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[4],stage6_8[4]}
   );
   gpc117_4 gpc4441 (
      {stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12], stage5_10[13]},
      {stage5_11[1]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[2],stage6_11[3],stage6_10[3]}
   );
   gpc117_4 gpc4442 (
      {stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17], stage5_10[18], stage5_10[19], stage5_10[20]},
      {stage5_11[2]},
      {stage5_12[1]},
      {stage6_13[1],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc117_4 gpc4443 (
      {stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7], stage5_11[8], 1'b0},
      {stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[2],stage6_12[4],stage6_11[5]}
   );
   gpc207_4 gpc4444 (
      {stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_14[0], stage5_14[1]},
      {stage6_15[0],stage6_14[1],stage6_13[3],stage6_12[5]}
   );
   gpc1406_5 gpc4445 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5], stage5_13[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[4]}
   );
   gpc1406_5 gpc4446 (
      {stage5_13[7], stage5_13[8], stage5_13[9], stage5_13[10], stage5_13[11], stage5_13[12]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[1]},
      {stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[5]}
   );
   gpc615_5 gpc4447 (
      {stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[8]},
      {stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[0],stage6_17[2],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc117_4 gpc4448 (
      {stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14]},
      {stage5_17[0]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[1],stage6_17[3],stage6_16[3]}
   );
   gpc7_3 gpc4449 (
      {stage5_16[15], stage5_16[16], stage5_16[17], stage5_16[18], stage5_16[19], stage5_16[20], stage5_16[21]},
      {stage6_18[2],stage6_17[4],stage6_16[4]}
   );
   gpc1163_5 gpc4450 (
      {stage5_17[1], stage5_17[2], stage5_17[3]},
      {stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3],stage6_17[5]}
   );
   gpc1163_5 gpc4451 (
      {stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[2],stage6_18[4],stage6_17[6]}
   );
   gpc606_5 gpc4452 (
      {stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11], stage5_17[12]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[3],stage6_18[5],stage6_17[7]}
   );
   gpc615_5 gpc4453 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[2]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[4]}
   );
   gpc606_5 gpc4454 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc1406_5 gpc4455 (
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0]},
      {stage6_25[0],stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[5]}
   );
   gpc615_5 gpc4456 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[4]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[0],stage6_25[1],stage6_24[2],stage6_23[3],stage6_22[3]}
   );
   gpc615_5 gpc4457 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[7]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[1],stage6_25[2],stage6_24[3],stage6_23[4]}
   );
   gpc135_4 gpc4458 (
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4]},
      {stage5_27[0], stage5_27[1], stage5_27[2]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[2]}
   );
   gpc615_5 gpc4459 (
      {stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[2]}
   );
   gpc606_5 gpc4460 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1],stage6_29[2]}
   );
   gpc1406_5 gpc4461 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3]},
      {stage5_33[0]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[2]}
   );
   gpc615_5 gpc4462 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {stage5_31[6]},
      {stage5_32[4], stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[3]}
   );
   gpc606_5 gpc4463 (
      {stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3]}
   );
   gpc606_5 gpc4464 (
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1]}
   );
   gpc1_1 gpc4465 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4466 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4467 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc4468 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc4469 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc4470 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc4471 (
      {stage5_1[6]},
      {stage6_1[4]}
   );
   gpc1_1 gpc4472 (
      {stage5_1[7]},
      {stage6_1[5]}
   );
   gpc1_1 gpc4473 (
      {stage5_1[8]},
      {stage6_1[6]}
   );
   gpc1_1 gpc4474 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc4475 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc4476 (
      {stage5_5[7]},
      {stage6_5[4]}
   );
   gpc1_1 gpc4477 (
      {stage5_5[8]},
      {stage6_5[5]}
   );
   gpc1_1 gpc4478 (
      {stage5_6[8]},
      {stage6_6[3]}
   );
   gpc1_1 gpc4479 (
      {stage5_6[9]},
      {stage6_6[4]}
   );
   gpc1_1 gpc4480 (
      {stage5_8[12]},
      {stage6_8[5]}
   );
   gpc1_1 gpc4481 (
      {stage5_10[21]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4482 (
      {stage5_10[22]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4483 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc4484 (
      {stage5_13[13]},
      {stage6_13[6]}
   );
   gpc1_1 gpc4485 (
      {stage5_13[14]},
      {stage6_13[7]}
   );
   gpc1_1 gpc4486 (
      {stage5_13[15]},
      {stage6_13[8]}
   );
   gpc1_1 gpc4487 (
      {stage5_14[7]},
      {stage6_14[5]}
   );
   gpc1_1 gpc4488 (
      {stage5_15[9]},
      {stage6_15[4]}
   );
   gpc1_1 gpc4489 (
      {stage5_15[10]},
      {stage6_15[5]}
   );
   gpc1_1 gpc4490 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc4491 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc4492 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc4493 (
      {stage5_22[11]},
      {stage6_22[4]}
   );
   gpc1_1 gpc4494 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc4495 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc4496 (
      {stage5_23[12]},
      {stage6_23[7]}
   );
   gpc1_1 gpc4497 (
      {stage5_23[13]},
      {stage6_23[8]}
   );
   gpc1_1 gpc4498 (
      {stage5_25[6]},
      {stage6_25[3]}
   );
   gpc1_1 gpc4499 (
      {stage5_25[7]},
      {stage6_25[4]}
   );
   gpc1_1 gpc4500 (
      {stage5_26[5]},
      {stage6_26[3]}
   );
   gpc1_1 gpc4501 (
      {stage5_26[6]},
      {stage6_26[4]}
   );
   gpc1_1 gpc4502 (
      {stage5_26[7]},
      {stage6_26[5]}
   );
   gpc1_1 gpc4503 (
      {stage5_26[8]},
      {stage6_26[6]}
   );
   gpc1_1 gpc4504 (
      {stage5_26[9]},
      {stage6_26[7]}
   );
   gpc1_1 gpc4505 (
      {stage5_26[10]},
      {stage6_26[8]}
   );
   gpc1_1 gpc4506 (
      {stage5_26[11]},
      {stage6_26[9]}
   );
   gpc1_1 gpc4507 (
      {stage5_26[12]},
      {stage6_26[10]}
   );
   gpc1_1 gpc4508 (
      {stage5_26[13]},
      {stage6_26[11]}
   );
   gpc1_1 gpc4509 (
      {stage5_27[8]},
      {stage6_27[3]}
   );
   gpc1_1 gpc4510 (
      {stage5_27[9]},
      {stage6_27[4]}
   );
   gpc1_1 gpc4511 (
      {stage5_27[10]},
      {stage6_27[5]}
   );
   gpc1_1 gpc4512 (
      {stage5_27[11]},
      {stage6_27[6]}
   );
   gpc1_1 gpc4513 (
      {stage5_27[12]},
      {stage6_27[7]}
   );
   gpc1_1 gpc4514 (
      {stage5_27[13]},
      {stage6_27[8]}
   );
   gpc1_1 gpc4515 (
      {stage5_28[2]},
      {stage6_28[2]}
   );
   gpc1_1 gpc4516 (
      {stage5_28[3]},
      {stage6_28[3]}
   );
   gpc1_1 gpc4517 (
      {stage5_28[4]},
      {stage6_28[4]}
   );
   gpc1_1 gpc4518 (
      {stage5_28[5]},
      {stage6_28[5]}
   );
   gpc1_1 gpc4519 (
      {stage5_28[6]},
      {stage6_28[6]}
   );
   gpc1_1 gpc4520 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc4521 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc4522 (
      {stage5_31[7]},
      {stage6_31[4]}
   );
   gpc1_1 gpc4523 (
      {stage5_31[8]},
      {stage6_31[5]}
   );
   gpc1_1 gpc4524 (
      {stage5_31[9]},
      {stage6_31[6]}
   );
   gpc1_1 gpc4525 (
      {stage5_31[10]},
      {stage6_31[7]}
   );
   gpc1_1 gpc4526 (
      {stage5_32[10]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4527 (
      {stage5_33[7]},
      {stage6_33[4]}
   );
   gpc1_1 gpc4528 (
      {stage5_33[8]},
      {stage6_33[5]}
   );
   gpc1_1 gpc4529 (
      {stage5_34[0]},
      {stage6_34[3]}
   );
   gpc1_1 gpc4530 (
      {stage5_34[1]},
      {stage6_34[4]}
   );
   gpc1_1 gpc4531 (
      {stage5_34[2]},
      {stage6_34[5]}
   );
   gpc1_1 gpc4532 (
      {stage5_34[3]},
      {stage6_34[6]}
   );
   gpc1_1 gpc4533 (
      {stage5_34[4]},
      {stage6_34[7]}
   );
   gpc1_1 gpc4534 (
      {stage5_34[5]},
      {stage6_34[8]}
   );
   gpc1_1 gpc4535 (
      {stage5_34[6]},
      {stage6_34[9]}
   );
   gpc1_1 gpc4536 (
      {stage5_34[7]},
      {stage6_34[10]}
   );
   gpc1_1 gpc4537 (
      {stage5_35[12]},
      {stage6_35[2]}
   );
   gpc1_1 gpc4538 (
      {stage5_35[13]},
      {stage6_35[3]}
   );
   gpc1_1 gpc4539 (
      {stage5_35[14]},
      {stage6_35[4]}
   );
   gpc1_1 gpc4540 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4541 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4542 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4543 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4544 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
   gpc1_1 gpc4545 (
      {stage5_38[1]},
      {stage6_38[2]}
   );
   gpc223_4 gpc4546 (
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0], stage6_6[1]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0]}
   );
   gpc135_4 gpc4547 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[0]}
   );
   gpc615_5 gpc4548 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[0]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1]}
   );
   gpc2135_5 gpc4549 (
      {stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage6_14[0]},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[2]}
   );
   gpc615_5 gpc4550 (
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4]},
      {stage6_17[0]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1]}
   );
   gpc7_3 gpc4551 (
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage7_19[1],stage7_18[1],stage7_17[1]}
   );
   gpc615_5 gpc4552 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4]},
      {stage6_20[0]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[2]}
   );
   gpc615_5 gpc4553 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4]},
      {stage6_24[0]},
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], 1'b0},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[1]}
   );
   gpc7_3 gpc4554 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4], stage6_26[5], stage6_26[6]},
      {stage7_28[0],stage7_27[1],stage7_26[1]}
   );
   gpc7_3 gpc4555 (
      {stage6_26[7], stage6_26[8], stage6_26[9], stage6_26[10], stage6_26[11], 1'b0, 1'b0},
      {stage7_28[1],stage7_27[2],stage7_26[2]}
   );
   gpc7_3 gpc4556 (
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5], stage6_27[6]},
      {stage7_29[0],stage7_28[2],stage7_27[3]}
   );
   gpc1325_5 gpc4557 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4]},
      {stage6_29[0], stage6_29[1]},
      {stage6_30[0], stage6_30[1], stage6_30[2]},
      {stage6_31[0]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[3]}
   );
   gpc7_3 gpc4558 (
      {stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4], stage6_31[5], stage6_31[6], stage6_31[7]},
      {stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc606_5 gpc4559 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], 1'b0},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[0],stage7_33[1]}
   );
   gpc606_5 gpc4560 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[1]}
   );
   gpc1_1 gpc4561 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4562 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4563 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc4564 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4565 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc4566 (
      {stage6_1[2]},
      {stage7_1[2]}
   );
   gpc1_1 gpc4567 (
      {stage6_1[3]},
      {stage7_1[3]}
   );
   gpc1_1 gpc4568 (
      {stage6_1[4]},
      {stage7_1[4]}
   );
   gpc1_1 gpc4569 (
      {stage6_1[5]},
      {stage7_1[5]}
   );
   gpc1_1 gpc4570 (
      {stage6_1[6]},
      {stage7_1[6]}
   );
   gpc1_1 gpc4571 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc4572 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc4573 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc4574 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc4575 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc4576 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc4577 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4578 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc4579 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc4580 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc4581 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc4582 (
      {stage6_6[3]},
      {stage7_6[2]}
   );
   gpc1_1 gpc4583 (
      {stage6_6[4]},
      {stage7_6[3]}
   );
   gpc1_1 gpc4584 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc4585 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc4586 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc4587 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc4588 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc4589 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc4590 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc4591 (
      {stage6_10[3]},
      {stage7_10[1]}
   );
   gpc1_1 gpc4592 (
      {stage6_10[4]},
      {stage7_10[2]}
   );
   gpc1_1 gpc4593 (
      {stage6_10[5]},
      {stage7_10[3]}
   );
   gpc1_1 gpc4594 (
      {stage6_10[6]},
      {stage7_10[4]}
   );
   gpc1_1 gpc4595 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc4596 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc4597 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc4598 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc4599 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc4600 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc4601 (
      {stage6_15[2]},
      {stage7_15[2]}
   );
   gpc1_1 gpc4602 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc4603 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc4604 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc4605 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc4606 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc4607 (
      {stage6_20[1]},
      {stage7_20[2]}
   );
   gpc1_1 gpc4608 (
      {stage6_20[2]},
      {stage7_20[3]}
   );
   gpc1_1 gpc4609 (
      {stage6_20[3]},
      {stage7_20[4]}
   );
   gpc1_1 gpc4610 (
      {stage6_20[4]},
      {stage7_20[5]}
   );
   gpc1_1 gpc4611 (
      {stage6_20[5]},
      {stage7_20[6]}
   );
   gpc1_1 gpc4612 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc4613 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc4614 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc4615 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc4616 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc4617 (
      {stage6_23[5]},
      {stage7_23[2]}
   );
   gpc1_1 gpc4618 (
      {stage6_23[6]},
      {stage7_23[3]}
   );
   gpc1_1 gpc4619 (
      {stage6_23[7]},
      {stage7_23[4]}
   );
   gpc1_1 gpc4620 (
      {stage6_23[8]},
      {stage7_23[5]}
   );
   gpc1_1 gpc4621 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc4622 (
      {stage6_24[2]},
      {stage7_24[2]}
   );
   gpc1_1 gpc4623 (
      {stage6_24[3]},
      {stage7_24[3]}
   );
   gpc1_1 gpc4624 (
      {stage6_27[7]},
      {stage7_27[4]}
   );
   gpc1_1 gpc4625 (
      {stage6_27[8]},
      {stage7_27[5]}
   );
   gpc1_1 gpc4626 (
      {stage6_28[5]},
      {stage7_28[4]}
   );
   gpc1_1 gpc4627 (
      {stage6_28[6]},
      {stage7_28[5]}
   );
   gpc1_1 gpc4628 (
      {stage6_29[2]},
      {stage7_29[2]}
   );
   gpc1_1 gpc4629 (
      {stage6_29[3]},
      {stage7_29[3]}
   );
   gpc1_1 gpc4630 (
      {stage6_30[3]},
      {stage7_30[1]}
   );
   gpc1_1 gpc4631 (
      {stage6_30[4]},
      {stage7_30[2]}
   );
   gpc1_1 gpc4632 (
      {stage6_32[0]},
      {stage7_32[2]}
   );
   gpc1_1 gpc4633 (
      {stage6_32[1]},
      {stage7_32[3]}
   );
   gpc1_1 gpc4634 (
      {stage6_32[2]},
      {stage7_32[4]}
   );
   gpc1_1 gpc4635 (
      {stage6_32[3]},
      {stage7_32[5]}
   );
   gpc1_1 gpc4636 (
      {stage6_34[6]},
      {stage7_34[2]}
   );
   gpc1_1 gpc4637 (
      {stage6_34[7]},
      {stage7_34[3]}
   );
   gpc1_1 gpc4638 (
      {stage6_34[8]},
      {stage7_34[4]}
   );
   gpc1_1 gpc4639 (
      {stage6_34[9]},
      {stage7_34[5]}
   );
   gpc1_1 gpc4640 (
      {stage6_34[10]},
      {stage7_34[6]}
   );
   gpc1_1 gpc4641 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc4642 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc4643 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc4644 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc4645 (
      {stage6_38[2]},
      {stage7_38[3]}
   );
   gpc1_1 gpc4646 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1163_5 gpc4647 (
      {stage7_0[0], stage7_0[1], stage7_0[2]},
      {stage7_1[0], stage7_1[1], stage7_1[2], stage7_1[3], stage7_1[4], stage7_1[5]},
      {stage7_2[0]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1423_5 gpc4648 (
      {stage7_3[1], stage7_3[2], stage7_3[3]},
      {stage7_4[0], stage7_4[1]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc623_5 gpc4649 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc4650 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc4651 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc4652 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc3_2 gpc4653 (
      {stage7_19[0], stage7_19[1], stage7_19[2]},
      {stage8_20[0],stage8_19[1]}
   );
   gpc7_3 gpc4654 (
      {stage7_20[0], stage7_20[1], stage7_20[2], stage7_20[3], stage7_20[4], stage7_20[5], stage7_20[6]},
      {stage8_22[0],stage8_21[0],stage8_20[1]}
   );
   gpc117_4 gpc4655 (
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], 1'b0},
      {stage7_23[0]},
      {stage7_24[0]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[1]}
   );
   gpc2135_5 gpc4656 (
      {stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5]},
      {stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage7_26[0], stage7_26[1]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc2116_5 gpc4657 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4], stage7_27[5]},
      {stage7_28[0]},
      {stage7_29[0]},
      {stage7_30[0], stage7_30[1]},
      {stage8_31[0],stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[1]}
   );
   gpc2135_5 gpc4658 (
      {stage7_28[1], stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5]},
      {stage7_29[1], stage7_29[2], stage7_29[3]},
      {stage7_30[2]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[1],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc2116_5 gpc4659 (
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage7_33[0]},
      {stage7_34[0]},
      {stage7_35[0], stage7_35[1]},
      {stage8_36[0],stage8_35[0],stage8_34[0],stage8_33[0],stage8_32[1]}
   );
   gpc207_4 gpc4660 (
      {stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[1],stage8_35[1],stage8_34[1]}
   );
   gpc135_4 gpc4661 (
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0},
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0]},
      {stage8_40[0],stage8_39[0],stage8_38[0],stage8_37[1]}
   );
   gpc1_1 gpc4662 (
      {stage7_1[6]},
      {stage8_1[1]}
   );
   gpc1_1 gpc4663 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc4664 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc4665 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc4666 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc4667 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc4668 (
      {stage7_21[0]},
      {stage8_21[1]}
   );
   gpc1_1 gpc4669 (
      {stage7_26[2]},
      {stage8_26[1]}
   );
   gpc1_1 gpc4670 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
   gpc1_1 gpc4671 (
      {stage7_38[3]},
      {stage8_38[1]}
   );
endmodule
module rowadder2_1_41(input [40:0] src0, input [40:0] src1, output [41:0] dst0);
    wire [40:0] gene;
    wire [40:0] prop;
    wire [43:0] out;
    wire [43:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[40:40]}),
        .S({3'h0, prop[40:40]})
    );
    assign dst0 = {carryout[40], out[40:0]};
endmodule


module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor2_1_486_32 compressor2_1_486_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4b11e8b49eff62d20319ed7a0dd18a53942235ab795fe2c8ec5bc41b507b05dd671473cb0f0424ea435faa2db41eaed39e30d0e58cb65fd2f9124384c90f59dfc27435d8972499cdeec4238dfbcf958a7e9db86f71cff6e4f0d4356dcca9726392d90758d941309971165fc91a707efe7ed6002efba79725de9c003ef202b0137ca4d91e85bb3369e3a7de8d2132bd717fc1fef1c7ade77ba31408ea47ff4e63d96c27f745b5f253808e69a0118e43c89fa715171ce30c757bae9c518e1c17d9aefc197721e408a4ac1ac55a6567dcc61f588d02facb43f7b89774706cea163605fa8daf2d77d819533ad955f1c5c5316f8f55cbd86627b91f81274ac94653953414654568fd6825f20880eb7f85661a237671ca28fc1dac7ac58f3598508e01e7320c25d0b20fc9546954aa53b3fa2edf8dd722316a07ae82c873093ea91cf859e00cbd4b6f1e4905b441bd18fdb1e53562a35cea99414ef29b731e54d7f6b667368776e19460a88c0f74e31652c1b9ff5847181f6378cad60a353f519db6411a5afdad64a3af48aff2dc8f3f12c8cf9cfdf80118c92cd8dd812bcc65a48c488d7005b6f926476b8e1c2109b387344d305ab8f58bea7d890f47eb21491c84196f4ad00e4b521587a36b75ae97425a2181ff12445bf3a9998e8bbc477a5bd78afd7bc1885302b88614d11981fd3e5764b1bb22b42e3a3ab83f1921250924eb76c8c556b0a8a4b3ee420c00054dd722e2ed28a90b93f7d7d98cf01100535fc5b738f9f8d5fd7154de5e872be9bb61e9f056d26478b9db522bcb96eef384d7351451a2e9b043354931b1d6d99e8fbff226eb6526b83a61440c71a1aa7e1a6cdc5f1446f52d99a932201f6e80a207367ec12666249df61acff8ddc800a959601dd5e817361df1ea44c8061ce4aea4551f99e9fb819df87029b160acfbac39fe96cfce460ecbaa172781ee626b060aeb8e78cb283756e96d2edcac4122ca26bb4fb4f5c7727ab73e8fe71bacf7993df497ea695d0c86493992a130efba7112c0ba91ae944766d87fee62e914be1c594d0bf55f9dcf710f91d72875cec3a27d079c39d2479b7eb868b5c02230e5c749024e2e29ae366898f7167fb4e0f68b2182c3da9c6c35dd69b7c7ceb4093c5563370ba83767b54e5c0d46710ba106df6a82f89ed09d7e3eef1e9818f84510fcfd0e0e6a76969e56f6b976519bcd7d18e588a4a64f2cd33da182f916afc084c9ac84cab6653803e61adde3440704abf4b28c877b578eb647d5ad8b7b2ce144f0d84c0d3d81cfaa3f6251b5af62688a095cdcd9ab8f05c13562bbe601db2d18e175229b2b1f82a3163d4952c0f76e5df4c673a7aaa68d69c9573dbd565cf02824e1f7201250e25b9d5ec98e381c1193bab47cf106e6117cf91e2909b65add8428c4fce68cca41865d5ad80f3af4e70fb326d065f5d4ed8c5743f415f3f9d2a64647e2f751b1940a6f58b83af2149395560b0df1ee174de6d659d12fead5f2d027a7470c9201dbff3ed600bc7e9c9d69dc030c52e3d14cf9c7127ed238fbda56e173ac94b1bd280d78fdca6f9297b3eab883e9beb17320e79c90e1c46e13192204b2839352c6f91ce4b10c54cf1ddc3f981a9128080e3f8b0a8700c0e5e5d133bd76cae97dc3d20bfa95ce32b06a768fe063f3af64a69c212443b2ba776b70b803bb93133549ac9aea28fb7c7dafe0cdb52a867e9eca161df20d5846f68b2ae71dbada3e6561c86ba53b293b23393398c85d5ac8a952e422bac0be6a756c95c98158b82c6ec58f7ccc79bcf3af4241ff3856eb20a4db11239f2509635f0adbc6bd19b9d883e416e09cb4216f37f3f82e2da33e005888acb2054a76d5ce21ac8556c90aab8d612c71e31f0c0dd94bb01f4fbe443af6d07ad76302ee4691c4d6f269e0c56df86386a0954ce3fb25616b17522447ff5c19e5b63cf7c9b1386c596684b53f380094469559df474e93dcc075bc06708d9f1bbc12678e7b5d7293c8353a238eeec9ecf3f619b736cf3213382088d880e2ccd3a39608ee03a6868598bb7c5e78fcf74b2f9fd26df73ca896e95c88fb5ea81578a95e49d8de719ed4f016295a2d5a53b009c1e0ed665992c59ab9d79ea31a9b10eb1b20db43c9fbfae43ce30382250a431512481c770780d8f051a467f58d37e1335c00f82ac8183d7e5849cb9b53cead40cc3a2d7de9e06dfd363b34ede0ff8c3428dd841d4d6ae6e74547a8dcc8ff953a11bbfa941c6365eaa7a2baa215d3af4164f321ea90c42d4acad4c083e1b33983445a7a2cfe86ffd7be637e39e1c2af4f325e4267cf1413ee7c2daddebaa6429bb230346c26a186d52bcfd9a0632acbd7167a4dc7881ff404390075954b14c1899f73db05aecab4b1ffbb39af911c11e7c18634d3f5c90122449789227f84ffde8a7b6204cbdecfdbd1a5f8452479b31fc6f410d753dcd67408dbc7c87c55a3b5cef72cd61b5c15027ee88ff38b72c253f7ad43659211c1cb332f4492391043fa73cd20c9df9d58bae02ab7bd016949b24f8ae0f701550f3154f8e8006c164d0a4f3cd900e8914512fea9e0a15ba689ab8a9bb27f62826b4bf0dd2f66c62be97d6cdb6dc673635ba7f2e5e7d701aaf0ab864c27640a093005e79e396bc3c9b93d07e8343cf08f8bdc95f7f935324e7164db395adc399555ba904a327290feb2687ef091eefc2f05bdda8192bef9601cc52e9e475fae39a8c3d848c04556138543d39125e4c3b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h17d889f7b42208182494795e7a3d2230256bf56f81ab3f442837c7f94c8fd414a66c197b6b394a3b152e2f64139eff450077b294ae5084460211bc63921d17d6d95196c0132aa41e9eb8b3c9eb474a48769bf85750f1547941ecb82eb631776810cf266ca22da12bd71fe36024e7a4a1a655f873cf3ebc40ed2425160a3dbed372d990fa86aabfc807c5cba14e3fc48b61b0231b131e68d2fc0169b5eacf57513096288d42df4379d29c95c66ca7c7e35fa0c4a09135a71ec8055d7a25922af773a640c0741f64353abee917093ff9f59e8fc3b71d417b3102d188eddbabdd0120345dd86855d19a39f93f4e482faa537f2a0e38a47e6396db8e280fc59aa831c8eee9d0344f6a7dcc108cda79e0899b5d1f389e905e7bc6f4e33695a251758869fc611e4d9e474059590a9dfbaa66df9d628ff5dd20f3be991919097e874aacd8c7d437f69705e3032ecffe8e04c0f6e277d984b667f025c202e6859efbb8098cea7c42b02ac3adf2de44b5749b76450d45e15c7c74c66c132cc2965ca5f4a3425590c932418a2a0c8c2e762c66b73a492c92741ba629b2233450909e40a8379be0e059a71bb5fa1e4ca35a1aeac25e35a24373c44bfdae7c1ee01669a55861942a55c94d2f4f9363edfa773a34aefc6e30b3bb6e280ea8f508333d714b2afae197bf1e3c526209eb098e8cdbd0fdb4beac103445c43a2baeec7d679c916027a425a732f26184dac571d81c23d506e512ac3566f77daaee50e1caf2c8dd20148dbb9e2cd3241fd734491f28ed5f868170e75e38d35bca905cdc56832109f8a4da97894e4ba0845ae8f63cc6cc2e31d67c4ae9726c035bfe474e0931cf081f5fbea0115813ebe7a71ffb78a3cba09de60dc765aaad2f589d23c8dfedd3e9b12acc617b447da51e5afadd5919dd52998a707cea538e6110873bafb898a710595bf731fd69cee8771f8efbf5b97564e867857a75ed459d213560aa2b5b55e7c1d1eb4f68b5d485dddd438f1d19110c0b0baf39a666df94d73bb8844f3291ebfc9691ed3833e92613251414c3186ea8378f0f2342c6f70c022252a14df0a3e16957ec898afb5999349de8483a7b7c7104737b80d02f547ee468083d18f5e1d3b3dbb086ba68e2fd2ac3a16f82a12f198f9568654316599d962fd12d7083e7afc7ead8d0a9af254686bb5fafd5b195141006ee7d0204cc4f629bf3988e9a6a7ac5d7846561f894df37b39f4a1575b69c1349fd3111add69ff80b444e7f35a6f95c8de8cc69c4ca630f0cab7b503cae850c68b3e4d5b2ab78133d00f61d0e08a8bd0d5f75fcd7730f5b7847cdd5ea5d6966373b8c4dcba23e4ee272c8aba633cc3274d6aafa8060c5aa731fae26d2dc051eae99ea3acf8d76e17fa791ccc78370b5cd57d15702f08ed86b66fcfc24084d3f11e8d95566e01b1d386a0f590af46e107f3622a9a4d5d111d5f8161986f8d56b312b0238e6f13a2e2d11f4c6596617907ce3f72af3ece1ec40956adef83abf74893ae7820e1d5ff273e72c5b394e42aeb9b389469feebfe2a5b9dbec9af0ed8e1cd3c572c431d119fe68792ea2287c8a3bde2440e00fab9bd6c82c8b3e28486646c9c52d40bed8c9c2b998d1c0e5d4f1a9fb73778c55d913802dd64bf84cba82876eede2f1674d09e6b3af85e592f8b5ba6c325ebd0d640d93acc06dd0f0c07fc74da9c716c1e7ffb11f5f2661ae1a26c5769dae4e2eef436cd8190662ca8c741b68ed2882130d80183fdac7216411c7beb801f6cf0fb5a83dd0d18a8133bf354677d4c502906724f9bd4907162d09efead3b0165d5bdbfce312a0a81694b81cf89793306c69ea8f135104c89a147300960018c1560b1821b6339c9e5a6c0ebbe5f1adea231a6afaffa7b175ddc790633a7fe6b7b0f94b16bc96d82f6bc5e59d0b8fef2e7f38c37cd4d1ae3f07f97c17b985daabba7c090d964ee09cf017701957c163d8d7c9216707fed71bd339df6511acb52bab3bfc6502a9e50e21d33e5a01f684f6e95dd5f679305ebe6ca258a69aed9db42f5116256d3d75fa903bbfef13f2304c1acf7dae8f05b1227f5d6c0122a03657a2dbb6362ceb5d9d7b3d12a9579018e7695481d0900679a7f889fe61be41e8387fa43c48b58231ce257cb664b67a97ceb47e1822dfa6fc1d7e53be746c55afb4b5617e65e6ea9aebb3fd8032708d147c0217f6b95de4e5d8b9746482155724f2ff5cbbf8c69285101f4963efb8d1c3ec7f8fe342d343df8dfbf0d60d5039eee514f97e39973aa575ee55963d417ffc5d4877294c4206fc9f357433501d69babe3c3f0080b2e6a3fe4a35f40997acea64512b8f13bdb9758345ae702093ead837c8a8bbdcbdea046f656783effb2403e16e45c0e7b70e338a155d516a55c1463e39e863f8eac44f313849efdc3092344466e78c28681da42975916581b88fb38fe3131c68c6fb4230eb2a400d880b7d06d783438148962c6ff8224584c710557a310cbed41801bca9da734e9a1dc596b7a87cecc4efcabf436fd8868636a35b8ff89cd42a039ba56da3e38ad10f30959edc2cdebaf8d4a0909622cf166d18c5fcbda9f6984e0d16da3f3b34888fcba6d2378d3a95cc882e702eca9bf1b495277f6685310b410659f1c8eb3b4f50c9948b4fb4add416f8944a83e58bbde24226a8621212219b0eacb42a29ddb3dbce775c804b75660828afa09fde90b632d4fc3588c7cf6b50a2b7eb1915eddef3a84b4a40983a9dc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h66823b4f394cdaf35be4e423a6497f8a474a4131c82c0b99ec6529e66c7d07a3a505bc2270c4b540e75695f2549ac154a08d425c42f63c6791f4c1727a302edb7a44c87ae09b8f244ae9c5fefcba78a3e11bb40bef4bf29a9c1b0e11eb3febc1d1742c5f83aeb5bf31e034f26ccb867ef2bf6a412967f834a64a745f9bbacc98fde5eb573da03e814af269e6cd5a351f470072061ad4e770b381a68017835f4bb1b5f8934d80d1a379c78f8acd0c2b06ebedd369c37210725a28150e48e8c5ea7e89c542bc1eb12e8840409ee9ae56a4169f9797210d703e37ca6db657d9ca0badd7e92113b94cbbd476c366270f42b49f4f6be623c9f1ae77a9082121f4e44a0d37fef855f78aa6866c1f91b948a581221a59e13f8a288f32443c0cb03da0e95b586c428120169fd02d56957665ac9ecaf1ceb8beefb692c726c6b23fc4b58ac3d70d9940fbcb2822cb6a17d5c5c53e71121982723bcaf063cc0e3333f33c5689dd5db83ffc8b30e3f05c1e95aa8acfcc4300c40c0863a9d12b6fe3407fb52a04346af625f14cf8365b00f3311b97d57eea1a12bf2b56b1c8f0889c43c0b2f5494c35f7cd0746e1c58008d7546495dd5238aab7179cdefda9c7c552ea42b6ef2254d003e0474d1b6a535058d41d0aa5235a968843742c502bb55611f86791333dc01f98108dd9f692454b798f4601146e34aec80314d77d70e4b3ff1552c16ddeee8e262195622d40f26a9d0b4d08dd25e0aa22fbae7f5adf8cbf9477db398f4680977cc888645c19d05ef4b04e950ca5bf6637bc2109d4d3b40c6bbc58cab02799c3beb3adef4f6705d1f930d889153354910d6c3dcca7838ebd9582e2a9dc04ffd6c8e0401680012ba0a1762a84de06d2edfead5af613f8de9c5e0b631e8ad932a7841fbf4b659890c3ef9c1f826dcd72c1e1b2b87f05c8a17eb4715d8a33983ad46aea6c165170aaa87e48c8d1e2f6e051d4f9f53442b05369114e6c94bdcb6d538a23cb954691388049886e69fee7cd69a0de0496f6ecff14480e7d2f8e44ba5f077da1df77ffcbd1f9690b1566aa0d872b0478554ef966417227b7e45150dbd832a93e411afb76cb6723c36c94242a54666662e344dd287579c161da5dbcb7cbdbd5ebca9c168028e6502d4b953c2286ddb034e877b120f9d39bd8f9d3a11671649cddc27af5376cb8343da1046e2bcdbc9c824b18f66769959c98ee0a86cb1574119a3e40d2d6c96e8e502614c9b1a1d62cce3ee697686e1f853439e21f5585d06960745c6587fe97678f2b2dbc65d0ce5da876253959f9152bb494d0603f315cb1c75ebdfd6a6290d4e5c72fd20fe72a80d64dbf35eba94a756ea3e9bed44b750ac40e1f68ddfcb3b27e34a4823674ba5d4240aa11cc16aeccaf24413f8ba8347ed08ab2748652dcb87b8eae31078edc091506350b0ddb6e2e00b277082a15fc918c610e96026772a59d5c161fa02d26d0a744df56cb96d91c729196e2b51f3a21e238ca81e9df7c6132f159a5ba9f1ae3d69d817a98a949958b9b1380a10bebdb9568ceab976d1094027df03f7ab7eadf71160d8e410797469499210a0fbbff29816a3cbaf32fb237a57146e4be0ee37d6b6340d3e91306106a4f34d0a12e9a251228d8250622617ea632bf05f0e42bd9599869ce598b98de8318b083be0152b3aa31302099ed519d01568bb4a202cb2569f31542f6b4dbb03d141930b80cfefe9a730b3f04fd6b30c04d9b814ea7ae3a782651f7635e71ed1a28893d8a0e52b170cdc4d632836c581ec25985ecfce1cc9407dcd5c9829d53ab3f7cb70f586ef3be0281f85d844fbcc1ae69d2c4affee08a40f324422b2f789e8ad1e048288b2c267d39e1c8676d46123e717643feaa78e4a45b67dff2bbee3a29b413a3e53c9f55e643509c02a09bbeea578aa67e02379146b870f9e6c60e3f8a47915bee81b93ba03b14c79888a1a78178c7d82580bd5f94008e662db35140bfdbdcb26f765e939adcfdadf1fdd2ceff6b4f217f65b280130a986a72a238aa8569f82ed04ffe02776600063504ef8c1a66a967713f2982be4f25b65da01fa620accba5eeec174a26e141dc50da0b1aa679ac11130f4e4520171f0932d1ad3066cd59f04a71026504de57b7ebc12c945a72e5eb761883167beb8b6758f52b8f28956a264076424651b326fa999b2bfdd16f4c7957fe88c1eee2d5d95306a6143b8a34aeb8c89ac6c72803ad3c3682a634e026fbe85ddf1b3a46b6344eae7bde81152a160bfba405e00511f7e6c7fa215afcfaa63169777315c81a45d4b723efd5d5d98911ece13db32b8bbfcdc820f3572b1d1b0cf136602f16226b8a0c71a2b06fc67df8bcd6423bd076e351f1ce1b6b85f803e55ee2aff13dd6403ef96963622331169d6ca2ef66a9bdcebfe831338052e5fa49e09f555c7d24a3a8ffaad744a9236d91ba210abfae7e1d611179058b45ab700f8eea5a1c612e8588b7025fe5ed005327093d30af04522f49a4d70307dff494ecb4030c56de54310cbe03bd3a0bc56a5b6ef2dc5c5f4f9ca8cefdef498aa3ed2ef2b394b02bfb88c5b2ef51579bf725bea8f61687342adb89f8e6cb4442d584a9b119cb602383c6738c336b1a404ead86a8f7c330976083381ebd70f7b6db78b97141704bd8e14ceba59c0286f612ee18181561e79f6626ea965bf65998819bb8d67404b2aad500be0ee18475636eca7280aefb6b82baad1b1356be1a9d481a90efc25d5991;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf3c818fd74ae9dd252c9ff5da9271587010cbfff9e94f7d977ba49b33878370e4bc59a4a00ac2c74097cecb74aef7c96fcd1dd549607507351349790e47715cde4913448f1f1ef72df4dc0b812272f513c20d818ba91e1bebce920b0aa4d016a93ff2251d520343b535b436073923d3a75e97598c12e23223738e90a20b575d1939d52bff4f14161bbb6bd212992e51b494c28a29b05f6682208625f6aeeb980bdd0d9266efcd2a6f60ad8eaf9508e1230624f41d4be9ff1158d988c44afb3144e5585a34ed8d47eec93e49ff340c592950c5b35e736af87270fa9def614ad7ac40079ac5093826aab432bfae31218a692072e9e2b6d49562e4b5c087c9abe365bbe293362788da42385f41212b4c9c97c40ad9d23d20d9873d1cbe4bfe293581d60b2fcc63ef2151ee677e7bdaa49ff38de63c85b890f7f921c534eee0f0a520c7810b146414b2b388324ba07773acfea45122a7f030af9adaa8370f2da577bfa55bb4d05b5e999205a3f5422d2c2b761f2a0e9c3a77968dac85cf50630cea4a17c5a7cd87bcfb9ce8437dcdc70fe0da8b1513055f37c70e1589114aa059b52457a4be0fa43ff115237349a26c07ce369b16a819ab9fb62b664821b3eab8ebbf2e88fcddaa729b065679f8b35bacc6df9855a070f2785f9e1c65c89a8fee49afd90c23bd4a08c0df1f5a8d513afa3f4792ade8b971e801cc83044a2ed72b02c96e4815445c6223bacbe4a73a421f4c3c646b1579a65a31666a7daa73505e8451c625e8dc76a93945acde3477b0e7995d2046dd9edbdfc22771207c0daa4382c60a71dedaa79abece5a572c183a248753279bc3e1ae3649d1669ea2af213a5a8edaae5c3735e809bb545b8f797fe26604daabae4309dbadcf6707fce4b40ceaca6c33716edb4a4c83cc318840f9884cf94e72e0679520a5f22b15924a8ff00511ccd0e426b8eceb31754e70cd541340664a5d794690434a16e5327d48142afa4ed27627ea979a42fce98f1cb267cf2e5d086ab3c2adeed8d1565ddedd321c8dd96471af5b174956be71ed1c89626cbe62c31cc2a1259266a68ca17741ddda4e4b7dc3d618fbbf1da5e23e326ad8c31739edca6d96101c1b1511a896982cb60eb932a7fd0ab62fee31460cf5b37efdb9c28aa9fe3f98a1764bbbae484812aa43c611c3036e5bf78bbb0fb48b21076cbfcb9a68875e6dcf3fe51c8f2c8a58372b256135b83dfcc1a4164cd994c570d9a716d47644846d49c9f674d1f02f32bcbf9dd55d13379df265ccf78b8073811842ac4c16710af7940d6eb8efff59401d66431a9e900482b581c1dde3d9767112a1a2e8eb0ffbad86a9625b82af1e2cd75bab90530b83f941790ca0b1a0a1dbcf781448952f97a797a2abae425a143d204ed24e412761c0177500b9f80f30a797340f18e906427c62169cd2cd0e3c3f4804844c9e332f93367a1662f0efe2f24b7363d2d41ff2503e9b1e48c78438e1d3de2f0a42fc3a230b03888ba744b43f3b59516fdda88ecc69e990a743f35d1fb5f23795da6bc63d7aa9a140c0d9113b84b9a46429d32bede825940288f0c093d103eb7ae36de3e6c96169838abd155c0332626edf2150702de9606b457cf29e08d968ae6cbadcf65f4a390e28da9686563bdf5a61263d963eff0e64b8b7703786adb339cdfd956ce1ff9fdff0eb204ced928beeeccfeecdf400ad416d6ac7611e74dda62ef67e059683cc0231309e42b16ab6e10b7ab19022fe94ada6721b73bd9792917111f933ce994b3e09a7c1475a01c9fe7e51af3fb438f2d6e153637666c5b99968aa53e142c09da535d7e1781d54d6ca688760dae8e5d235434ad4aa2880ef9beebe1f941dbfa55eb37f61574a54c57e4f0c8b97f0e8b353e6bda209eb471225cfc5b800c676dc333f5f606f2b34eab99ecfb3002a1a848e4b8cd11e39245200f01e8e35099e54f6b8bde97967e5d22172dacfca4f0fec0074de85d1a68c5cfb8c24c2fc6f2beeab8b6873295dba6d7015666b761639568c8ffba35f729739a5d5eacce7a34670d5073eb403f93621e00ff1ecabaaff40099859a745d389a46ca111427f3cbff7f2118ea44ee0b154eb3e5ea42c0e285d7292270f6e66eabcfbeab4c4c3a19650e8042f0abc08c695690d81a959ef285a94e2edd19c2134e6fcf68b2b97efa3cbdfd4da9be8858b2ce4ceec24444d379a4337bb8526959ea113c25d58e7904eee8df4d814aeac165fc07fb9472ed5d82e02c26bfcc61cbd8905861e1590d7ea82cfc6dd5a10079ab26d01f81ec3062e0fa697226798e75f646ad5481d79a4c9faeba0f17a74727f3df09847b3072c50137b5ffc1a6d2ad7554e3e2143fec0ac7851015589e5299f505fb202146a1f30775ea55471c733cf38ca32d3e72df76e34d5b1ad52d8b28726dfbdcade64b84e6d8d5ddfb094861480e5c72b4a62d62c4540ed1368924345eea30d14514615b374dc9e227fe794376872af72c698e85f8ab093e19ee7fab2fc4bdf93e669ad5af664ff0f075572d28d6aace75f87d96c816d5d9c67a816e348706a55b9fd2df3e3e12bbbf70ef8a688daf4e104574baaf55d9c6c7dfbd372366d91183d913383c2d27344965b07b6d28ae7f64e08e87a88aae56dcc4b998da7e8883c9a65cc3c58d862aa162e91a375917644be94ac22b58a1ef044c537b0cb5958dec47defc676232802454369008134da7b552dabd736fcaf765cfee908cac683c2390a79a7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h14eeb448d56b30b61f0a7f99c8a6314c035b65c309decfe7b153bc5992e90703104d0d07f01fec01c839ac6f1df11031b468714e043087fffef7f53290713715539a2fb02c7eed278ff2f2c0ce5c12e33350aa5659153802b77068083cbb4f3ac45b8ca140a6e813bde3abe274f464e858976272477e62b37b8a6a95ba37321297e74c888fffca160917bb71d04245ed6dd9237202f8cd513ed0e38021456089b8d40ceaf66ba3a5e74cca0681045e672f9cc0cc19c0a4548426db15a2c819c13731abd12f183715b269cd4ff4a15151dedb98677cf196c50895702a3a227b330116cc44dda6df825ca1ad5e8b13580bc60ec60f9993762bb9b7f294e6481da2f801393de9242edf2c819d7414acbc1d70ce0222a967809aa1b375c5b7c2f22152de4ec79d58f235c0a020a559c591317e9e44dac9714503739e1effca7d45da5f5998932d81b19f01832a83d49a76402b4a6ec1033c648727b2eabf4f8a65a6c914157a4b5b7712302021eb1d1bbaa8a34fe3efc0e2bd82fb31935d76d19258198f00900db0472aa55d7ea579fbcfd77413b93aa463960c5ffabd0b5e3a54a7f6ec7bda526a1ce7c1a4ef97e7226510a85ffe810fcc988efc1763e1fbecca38a35b3ab700888a05a4599df5952516a98f863cb9ab9f9367d58de9635ce764cad65af88107171734ad5a0d82fcc49b1567ebaccfd207ef586554eaa46a8935d934c0fde28eb43e2e1de50ab4142e03d95eb1937be3278ca95d38399826894e938a6c24221d621c52a434d485e54c8f4054606264694dca018ac1742b688cba16553a8bc383ee79d45372c05acf59637d4f913559bf6d3be2c61b5d2eb09dab2e9515d354b35734003d4486ad932e9963f25d8258bd01a2f0ac03037df9ecb12e8a62aa6755ad3f87991cf2ca4a4e9038db956572b0f92b2074a79ff8b8fc85cd2297fae7f153b02622ce63c47fee7e13a049e30d80de49399821a662f19d531153b399cd1ad4a42ed65bcbf0025078ba32e98f4fb0359c40ef2c87a7234ffd605c3886ff2fac15be4444bc1c1d7d22bf21afe55d60455fef2ce16bfcfb6594351ae7a0ff4eb4dfd30df4938486af9763dd365ff47111ddedaaaddaab3a1cd4eca9d533427fe43eb183f53e42ad013f802d71e779f97db85ffb02229505a45d4f2b27743ad2a24872cb0d123317b2b15c394c8d95e071d08b31d6cbb935865af5e7353f6fa16dadaba4df99399475949546a558e71bd9b59418ffd33da9fae09c06cb800dfc30863c0cb5c56900f1fe74cc0065842c62b358484d5300430cc155f94ced30d063782cbbd6422429660b532367a1badb5083937cf1c8ea37956ff73ce233ce8b343ee1aad9f05849a42e03af0543615de49f9164967a68a7480a54fdb87258a07f891bc95a8e40043273b8037c1983fd261c412689f2f5c86c536f28afdfe58f36a292f428fe22f0a0330c4a3ebd2b816925d8bed7dc7796f4d2dd560f0603be129bc76e68df53a2a6f5115d7691b5a6eae8b3f094ee67aeb1c4495c9d6afb372ea08580b8ae8389ff13b734eec932263105cec5992c9320b11bc8966891409a2fb7df431521bae0d1544b70a318ab9353275c3bf27710d6ffc595dcfee435d01764288e82d256716547caf1e229594bc38e438d7e3ec0c958caa71f26c20e0a9e58f67480dc0f489a3df6d4e2cdec3cec4c6dd790c4fb490b9e4cb1b3e82a8d84aeb8ef602acb8bfb533b5f46f71a91ba199940d8a5b2d73567c72fe83ee73f7dfac70245975e933d2b7bc25b4018e8a857c4f93db12165c02392c69bbd18df6e2a47de07d5540eb4f02a9886018f2ae5a06b7b08379fe2b15bdae4e1a66fb259b360989c57c4b30b29d33ad008d30bf9935a6cdf1cb1461e3ba71ab9df0236dba0fff5d44b6a2610935753f2823a453b4c2140801497a4ad9c6eddcc75aa4159a8d3af07ca9b79e9ec020f67c635d99c6055dbad370e84b84c6b6b8d781f45c5ab4222c0e54b5ba407497221e5daec4c65785b4457ac0d2488208565d15f24e95634e99effabc06f17dd8f7feb5ae4c9ba5ad9432219e8bd74af7353457e7767fe77e9f44ae232f7dbbc2d7fbd1734812d647da47e2d0719e924343d6a86fd7714282539f9ca7d3bdab1dc114c08bb037adf3e3b356c2397a1ec9ccb1881b59becb3d0e560107fe9d60985410a86a05128790ed191cee3525f474959ae8f879828958cb01735d60c141d99c6b9446abca130b422a3e143c4eb379771536eca9a2775d154c7b9321904ceff4d37f7ac2fe3a467bdf440d1e9b79a980cacb1d2ff811a968d7815f363fe0e5641f952d0699d331300566ff47b65e6fdf0d08e10591e015e9c949495b7d3f42879b9fef162a59f92e7862e92968b812116e49f95aefd9cafd038e72384f63c7cd972e98ee26152af3013ae02b09593d04959360eb95608ca87f031c23a09785b9bcff94de91b1425935e8ae2ad32e162492e1d54d67a38337516da07b1517046bbd9bfd75e7fb861594fc49ea13bb59bcbe305578d51d7cea3ef83ebb3ece83c90967eaa8088fc4e42ed73cb3c6184b2f5e6ffc66640e871e61d50dd6df5a4773e15d98291bf58fcd9549c5954c8e40f2b8cc3d40e0b93d47d9e366cb4f6eea4029ba39ce443c76d076fdf892528812b2d9c4b96a6ecc0fa7f5e13b7967c7b521e6e4616f01aeb6ed1a9e2243ce44fa0275e0d2ea27d976689e0d7e1d3a2343d39eeb40f0424a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h31c4da76f9299c50957d3c7ecaa96a259f051ea7831db4eac69d57287eca83325ec09de7ce2a49f8bcf443ac30b2f1674e08bb446f554ba6fda29b982690cc0b218f3cffef55ac3ce9429db9a5aa5a1da6c2c069446addf57455554e404edf2b74ef37337f742ad746ea0b1e007aad81a75179796cb2a7a28ebe78b85c9858beeb9036bf5e21421a26fa7586d758215c9060f97172722d67f6f36c32750e7cf10172a2d2747e1b55b65df1428e97d70a7ab639a13bb83990c61b99876a299c360d6004d7b2017a29c0881b09bbf83a24b0af77732413d756cf1816c675f13c63cc82d88c498ec4f61b75bc91b3834ee18905de1e1cc91451edab26a72d2a76a2f1d927142b2383aad49fce5213776ecc6287ba0c882ab120ad89339698966fb5efd71448da19424c853cd80e7ac92fa821ad155b5969da7eaa6661bd530bc6a3f50f142423fa0d477a23722e6c81f5d14e7f8d23093ca69a10a5df0d94f870ec3a447beb90550700d638e37e1b215f119748f29346be97fb46aa24fe906d336eb26eec52b8231a8a0da7266f99f2c4d4726205a4c27c7a146ea183496b1bf0ba39beb82677161dfd89eb19feabda7003393cb7022655fba194128cfbef0f793ac536b84d2af1112286353d649119bbbbbf03ffc6310abef6108e1aa03eccd3997fba0c3e1b2ffffcdd7b64aa7acf3c6c8366aae2ccfc0b186a017dba7b0084eb7f98b34e624a26ad8572642c878bae167df45b3bf0bf072f67d5acf2518f31733a8ecfba593918b907ebd85c1864cbffb1c56e47e2d9538097a8ed5a0494c859aecf3f748dbc82f268d170594e7d5e918ab0d89d2686ea3a82480b446798f06f1698b7f15ccdb895976ce94603719de0d6103a7fa2ffdf5334c2f7f5898e1c21093ad6cbdc9e5e7db18c2910b4f736726ec02927ab89f291ea09fa64eaf8c9f9b4ee38af6d8ca7c18efb1b7a44396ff3fefe287378e3615f78d6ebc17cf16d16a9dfb56804b0d6b78c49b34edc20bf2a86adc3922b72dee5350d89644fa385270d49321e68d6dd1986b10e1599ae759f4781d1ad066cfe1724e482f5b7bb3bd69fa88785beb1572df6883ced2b8bc6847a958d75ca606aed9c0e11014c6f9f3530a80bf1f4cbb296b790d54d44be08c6f92af99d4b37ff6ed0c24152105799d4d9e7dd7924d2bfc33a24a4040760699cf54f796b528cc8b65acac0922853f81c6a490065ec2eb6fef51c386da2f8fbb7a891c2b8a6ad05bfc4204f279911c620ada133badf5ccd6d29a94b3ee8a53c9a034156c26d6479c565078545c124e2bc44bc029a188a9811251239c43a55276f9fa00c7c892c3e5095a67ee89fe5c7dd92c04c5578b1d59abcbec235dace308c166504b202480f80e60649d1cb373f261ef8c086708a8f09f3b9de282448ac30dc245801b8373739797b242db33b4fe65b36d515cdb8c76acd5f610457e81f76aedbcf60d693f33829eb4e282c2a8ee22fdf3f32d24872cc873b33b541f2d59987b2650d1e1f5f6846ac5b5df683e29c9df9fae4901f2b89109c5715eddca20e1d042cd307d7e6e209ffb90278428282d111fec352ac9db996157f84065407495b1abb1ffc220f50700e4772c22ed0527cc576a233e705219a8fc037f4b873329c71190c256d35f78fa831783e33fb670801da9148a9d3e69edd90609989ff1fe3f625014dc8588cec94597f404adfd23ebeb19de9edf0b2cd7be56b1bb80864e4aaa466fc067351b6a7fba12f7bc44578fc06240cbdc506b9402586906d273bba607ab01fa20ba98115822ae34a7858b4eaa6ac0cf57d23f0ee61585f78850d07e6ff0ad4b0f81eec938f801a8db0b520cb2d0aaf866febf8c904ddbb15f395c24ff56f592669c120140768e5af28d892a63340d48ce1e06fa7435d3dd9af57fdbea1651288a646396f29072e0db50718786995ec47fed26a4b488954a60bfefd1c7aa71b13c2c3d9c8a77d393227ef1e0ee66cbde741729137701a2a0934d3104c7771b70977fc5e9bdef72d5d63b5a385c1be1165d83aa0adf849d9d9cf066109c360cb13e1509d73093abc33e653fd10bd5012b3cd4eb695c2df82daed75409e2f0fce75b3494bbce72e1d8597fb1aa609f6bfe73a75f5951c91b7c8627997976ebce3d7f102819a6299af876eec1be5b56cbd5c176eb3b0156b32983c98cf7d9127773bad15de57f95a31ec76f3ee6effa6696b6577f962f34daf37d9e7e673046841ab2c1e01e3b1bbd83c4760ddebb77b1eacd6b4bd10f8de8e42490f6b21b646b182467a7e11ae67fbfc57704dde3563daafc0bbc90b0b0475d63dcf9766db43fbc4a4233ff8aa368d9db44d468d09f4affcc6ea29f3c1ae40d22af6953c490b571ced2943037d669935ba0341d018707398e221166bdc0c2dc4b70b16138fe8a1829234d5414e33aa19d0aff0eaab7358f3ebc5954be0e224ff822e090446d84ed0bcee131a27a9c20a9c70eb727db0cac049d4eda78b0326e36b5c8424e485c43e477cbc9b34a7eceb46c4bccd129778a4980d9c8bf2d7bcf641d02c94f85f160638b417414031d81a0bffcdf03835691a017869503585673092aad201fd0fae03c2435e723ea9f65ba2b97b583f645380c4130bc5ba30a6f13379cea05a3a24bb66f24bc6c09b32d133391e5da9e498550dbae70b469e7c55433193dd7c44145f8be98b389dda21db363a6d92ada795a457b512036daf57d3aa6b192711f66cc05ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hdacf03fa743de6ab8fdae44ca719364c10bb8ce772349cf5525afe8cfe09644ab0f669b1a2a4ffcaca9e2635add36a8a9c2d0d485c33406670931de5292f323df5c94cd983d037fba8e582cec49e4f6539b5b161eed59eb9d79a5a36ea50d44b583c31b187948a841b0e67e540f721bde62f7ece175ff899daad4e905179a14baedceea455e49153f5b81daaeb3f29e40f4b60a6688d61ce777cc573cfb8fe6be0e61a5dbdbee652a188725ee7f46eb3a187ad283db267b874cdfa2c167350af67caaee7a296e5a8f2546089dae6efb62077261115fc2d9c062d7533cfe25e12bfb28203ecbe0f609f087296ef921b09572b4a668ffbddb7570342076be0746d0a736871421f3c252b9e5120385060c3b00973657f93a46599534206f41cb91cfd1deb55f8b7355f87f09fbfb58fdb3eaee78dfc9db1c20709b13c38bc9d3234e94db3b83fdf560cc336517da5de66c8ab730eba7d9253d5b2189feaba7cd06a699fdd0736415e641a3900cdc258bd21d6bde7503aa1e9635455b993537768682f4252c136aa6728f6483787dafbd60f8a1f280affc87ffcf14c94fa841d1086c47f41dea407d26be3e57feae4752a229efc8e926c30811d80969ab163ba0c4041247cbe8c7661978e6f7f2827a63c7bd390b98165281757ee28ee4b000458aae081c19f3264b413d1f21359ec90f2bcb9bf6a45e528d4f41a9c1e577b12472e865360df655df6b1705462cbba0ff336cd95c8a6d5a9a2c3f5b940c25aaecd3c36fcfa3206de377935b8a342897dbde34b59c27c66179cbac1656bee9c02d1cb71b0f069ab8583873f74f69ba17bc95ebed6a3b84d90a4bc5c5d93be56d754c15bc5561973efed725fe7d90ea3e0fbd931853518014df6b0bb525807d17be0aa5ed3943f04d5a89db974188f363ed41e57aa81383a3778fe4675638acf5dfc64adbdda284450c00231f48a081207672db151110431bab26c29ec1a6d7e93aa7ea72c935c82ed4960cda45db489c98af0e6d065bc321626155f63850d55750c57c00a3debc2effff0e8b817f04f7a952d5b08d053fa067bcee00693db36b2340bad0683b49244d39f29345649895b291ce2c916c9e496ce0e3f0875eb69068c362af5e7a20394112d64b1a94cb22ce5cce5f0f69584a83a9eaac16d2dd410a2839c0ac2b0dd88bed94edbb943ef5dc3d51b2db2983aabe2ba64e9d90b559ea2104133395b76da0f943561c337bd24d79e17ee0a0d7810ce6a90aa4ef8d18935d2f55aac34e9d58fcb48c30002e5a08d20c8a0d972daa40c17063515e8b17fb84765f385d4102da8944ccf2a39af2e80a8faf8f5d84faba1ab362c801d9f0515da4b9e919803118c52f29a3ad5b74ceeaaeae7ab021fccd3204b69b8b14cf7e4c76d37027ee60d2e851e823ec40a4074c3086749725e70ec18fcf5db67fedcc06f5842ea5d2d01ebb5a816c8c30fd7d00a5fc098bf555e8f5519dd936b7703d50a83bd3b79cc60e2920900db9d72b492717592ebececdb42c81bed6974bf52f94c77ae4217501f85b9008518a46d87aefecc84489501120eac3159154f3adde4f070dee0616fa7680f12afc3306539296be6f3ec37d00eeb149995736b06f097ced64182da6944ab6fcddec64a90d4eceff670a68a7b5aae54a5b8c8f67ae2f3e89f2c0da73f0de4f3ba24b235d174fb17b65d0ddba716499b120dd89c802dd4afe135fd8698071a64c0d7feb6f456ade94469234e75e094611ef80dd0011fa525d6a8c572d35c378346f56fcb33c4575e647c24b74156b615a5dfa83566b5ada250df29e1b0c0131f0db53a8fe483f46c1a2e743878ff12e7b95c6a69ba4c3702791976e8ca4dc4e688382c0eca0fafcc67b3bf5290034172e35cbc50cf0c7b2e9eb330cc6ba7f2bf12994aae6c27810717965376b1ce719ff0e2480389d5b068841dd113d42a62d86d718e6eb74a967aa5ab0c40592463f70cb7aae15af8b0f28f19bd45acf59de6a0942060f21ed16a7dfc8feb6694ce2829508b0764fea612481004ea90caf740da7cb531739d69c6ddcd1888b9cfc94f104c30a46187f9d73b250e8ef8ffd1933be0b8974c9f883ff58cf20d4be43b6f09407226509e9f4dbb7d228cb788965023f0ce871f1d6c231350191a01118bc7d7cf32e28dcccfba50aee3ad4b02978eaa49204157b3d6e3f2a0094763a7b2c5ff22381bb9dd94c34c83fd85af18cb8395dd4af3720f91bce29cb4e75267309d5e409a48cb7cf32c9561b47803c37456746e68fd69730a4bef7aacb411debefd9323319a655ed437345a06e4b4afdc24fddab531c623747d2daffad917f02949c8a5dc454cc4a19716d0131bd6bd9a194d4c3f043beb14af8822e32689a948397d2320e15bbc797b70f9bae904fa31a54dcf894911b5944d6b0b3cac24ab160685a03fae6c95563c50c09c5a4bad1d0cd668b9e93f571b1bf5fd95ea71b38049a6de7f4aecba64d206736dac9b03e079573cd83c06219159ce953af7966b241727e820d6058cf3c72b770febb751840c433f00f127e66dd8c228131e253f207eebbec3e575630d1272e2d4da0727b55f1ea4c9f22c0b3dfa8e4f34c31191469cb3b2afa8ca27abdffd591e51b651d5e584e143e7226b65961770e9e6587b96a230eeb33e88f1c3d4033aa2db57164079310012dbf2667c7682205bc655a9d5c23ca6ce3bfd6075ad5c705e5effb3838906d1e1b842d1ac18aa94e1298671cf72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h87ab3f21c5702e839c6094159be78f080ef32c5ee373b6b4f6adddad05a2a4e0a7482bb64f240ef236c904f48a497ca3a01610f9599c8ddc5390c7a57e775cd1fb85345198013e3ac316365174cc9359a734e86e91ce1f8942dc2b5f689728ea32e0fd74144383b55c11301e81215aa53f319d7d13eaf19c0057aa1ccf94b59feb3d98610659851947e874d3bf91b00cd0bac3d01c7da6e73a3e01c533c945f393470ad40ccc6b22774a5eb5dee8165d214bb7fb89efc1064b3d0d9c7df3c610af00ca83fe5275f7967e028f99f805e416451a3091c3f19985b42cb88fa4c9c1d3e4ca23c4a8554f286af4293c5cfa33a2a69ba42cdf5e96bdd05e04be40d1f05ebea3198161c604bb4a6b0ede8a64f698d34a71fcb9987902f149c0c4bf2ed92cad696caf186ed170a61fc01d9312c88807c83e3fee016b76af6eb53e8d302b7df4120410cafcaff62c68ab0bd64be9d75ac6e0b386631e05c0e0f3647ef5dace03b6f204eaeb0c7dab5652e29246896ca6b882362c4f6e58b8d8273ba1a72b2d0fea595554327dba319e251193d001d68e61833cc5770857f2a11e0553a060b4cbdf6f4a668a1cd7dd4f90c744a419684cd351e14899af368ccf929c3bd2b7b38eab343ab702202d5710034bd4217e8b6dfb005ba5a76ee1e302d05db665fb746e90b29e8d3393019439c674c9a58e8e7c10dff34fc542135734c9b38e885136b1588e96c1afbac9bca688e0f413b27357dc44d3e9453ff68678e6f7e8c746fc072f5c422c061057e338cc657533737cc037c076aba60742f017f161d54956a23c4c68e64653cc3c39c6663fc1792735bb386751b2ad6f61eec1da71d0685404366e7672dab911889021e4689cd45a591ba2916057eda38d666a3b017d93041d2204d95612887a8e2bac49345d337fe692f19918d7ea20758fcbe21ff58b0599d0bc4ad314d78f19f4bc559b6f04af3ff9e2b935abe5416e6d7bcfb2a7cc64e3dc9ac80a007edfc28cd60046c1208c8845c6a7137b61a837716fefb5f795855de84d64f8efdc4715ffcb2c2624e4af325f650843f5ac1c9f452f45f3450a64ff5ac26c795ea145a84538a7fcd1240a9d17160560849ec889bbbbbe7f15004c3c69691e493c48129b93e68efdd65d3630777ca8e525162501fc086d47587dd3f7018b0ce9a47fe49ceb6e580078bc7b1eb0ddaf2285f446b069fc2e4f838eb257cbb2ebff4b20708d708bf4e6872ba51fdb257eb35e71951d92d57dce7aca62709ff690e0c90b6f7a4ed58374ab587566251e6d9ae51198011aa35ef42c7cfeff4afec252e5493ebdaaa356403f54ced8a83634c02498247d4a9ae8d88ced76d22cfdf6d4b80d570e73b0b1faccaf5c239b05c6591f11da00f4650e514aeab0866428a93c7249fb33d433220d94469a6fa5f72564dc81df058bc4f75105503d5d4643b42b3da22653c67c06c9e348f310e98a4a8ae8afcc200c8f66c760a666a55782fe6f7164c02525cb9f1216c1af52033a9daad9850306efc867615459bda79dca0f25b56c4a7be158c14a9fd44255c58253554d7b3acc10ba78393ae8696352f708bb0e3219b2afd9dfbfa7433d321cbd156d3881aea65a0de4fc51dea84a31859d882ff1dff40fe8134bc3a2efa956ade4b706c9ee134d8d3630bf8cc690dcbb1b7f5b33cc0d2096d8517c50e4ad6d6f07f7902ff0c25e0fef586708f68aee5c8015646be000e893dd8269ab7a928817bec7c84d55f3276708fbc44470e7a1e3a2f5f258124b2f96af5d62a16b8330d37e560fe311fd9181cf4ce280b65fcf5d5212e3edf1b11f4c2940198ffc84cd7f177a71f4e8a1c500fb4eb0405e68d9cccaa7017fe44a6dc4f09bae110f6c7a19c346bb38aae50ae79dc6c94681c64d4bff386db059d9c639fbaea7326468077711ea07c048d5a329b8fba94eb9ef25681640fd9882982335e74554faf5a021cebdb5978b75afd787b3380cab886e6a040bf955a9b4c8de6091bb398688dac90bd70918b6667872b0e4e51b385d01a3299f92bbc156c5dde185f7028e2bb1aa31c03bbca024c32ca12f73b7ca2c39e227b3a8d8addf13046d170bf8aaaa23a9ab156112296278e79b606cb1be0d80a4f89fee3f015ada25ff0b8e4aa21be8abd9443566c4e3f12f559272368a3b9a2a56f3cfed9df144ce1beaeb112a25303d67699ddc08171d57b1c99a05a0df5aebbf77a6c1f37d1c194b065a75501b401a00734ed986597dad1084835eb54e9eba62d0322d540f78bad702268fcf8fd745062d75aaa3e71ac36b734a0156cbca90f5c57b2e01678a7d4192ae5bd92b680332237c9ba96e35f70e6514e54590db7d3b8b2bcde91ef9821b5d931f860d7c2fecb2e3b246ccc99d31858165924baeb101e28196f3c17e089e7d8b2a6d59ed95222746606be7b5a4cdab807b65e46947f50fc318d617942e11920136f4716532287d20d2ab3af9de7c89e237d9883193e32d1215ebcd946b022412c8e8b0e36df9bfe663f2aa58b88bab876d7ad3ccaa140b3827e6620caa1cbf90100f6c62788b0c01444203cf5f0ea0f3bebf0d3a1f5b1d50aa8285f7b0c7e4a719a68bee4031d9e69b074ec2ea3fa315c4d212818ad831b6d60a9fa971502aa1cf786aa68b213d8bd3b86a0bd79d4c27a65df12f973651870b282d0576865edf75ebfaf0629510ff6976e128a1f434d50d78aaad2307dcc4a9d9f2593df92578f2fb05d398be30b6d7670e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf68f3c63ffe5551aaddbaaa0d7616341d126a38a72dd5951c4a7fbca51611292bb53dab054101ad76fd90db8d0e3596e4a4215bdfbedec7581b654e73685eb1e6a6c54b2126df881763ce8faf99972a0687c3d615076cabbc960233db72bc409ee5eef019b9c45c299e49e25e98ffa9b24e879971fa53cb08b87590a4737c77147bf4271671a4e4959e4508f14c92fab137b03336fce38084ee1ae961ef1c6d8794482955b11f62ea11d9cb2982781d555c693127a2dfeeb7825eb19ad1f6ed1159e35e3b6e13cc8aa31780a878035eb9f0f231aaf47a4b83740ffa52215008ed4812fb7527ab2202e3509bd44de4607f40a2f7e634ae764dcf3813f3e765704f9e144737d1b0ecec821c73ba2251086df622d6655844159e3dcae40ca18cc6028b3dbd620e2a8685c7dd49f20683f0a0e19268e148dee295829ec4782729ca468016d0a40826cbf214e2597f2a17ed1e6c1fab81c0eef2cd2900d2782155d02b6211668fb0f663ae0f7e5e0fc9994cf5f17cf4420441920bd70efb3d6182bb54b9bbb863e4cda7a0b5959c400185c977ba51006e98d1092273dab37f5736ce41964cad40350ee12fe397ee1924f27520bf6b503214dfb04637c70a725048e1608c99da5af254ba0812c2ccd8b0431e7ab417f4fcf52179a26e5d497b241266bd178d016b938e3d6b3041026c7cb820b46809c339efd6aa64cd39d5b0a754f1af302fdbb2ea1148d31854a6d78c41fd8db763f8acf5ec9a0ee6b93a87e73b007af924dc06bb6a688c1eb2dc12a25131f44574505f707778220f5ae367fdfb380365d049b6c7f9b1b87933e1e2de40bff5980e32b81d9a44564764a2ab4f70f96067e509ad0185b807431c3aa0720111e7989715bd9afa7a8c9a9e7a988b1d0925fd65d535eb6935b051272b5d5efc5e2299b31b46adafe80d32f1fcedea786a93d6a3cc90daa036ae8bead19f24755d1a3033b82df5ed3ee250cd00f740817f61e51f968d6b10bf8dc8c513c30649853576698a64b5adf744aa0e28df7c9a12a5d7fa4f68be858f5c4a7c7344deba4e7ea2f98d52f4de83337a157d1ab4cf221c3cba26bcb8c28f34b693f2841710588078e45c9ce8aa9464be31ef0912482d8f77e879da571b3b639b92ffa45b11f3240fb7d72acc0277b5501a3127965b672575555a1bc62c960c87307b340d0c18b199c1f052e08ac924b0165d50d0cf2f768a17ebfd37e2abf8f1f39a33cdc429a9f2d7e38082f0ac2c958bbacaaa058a96e1030b86438301ab44fb0a24b9f3f9163e3afeb4d40e9f8912ab28a87ede30dda4eec2fd3aa6d29af395373b210b2cc30e0353e5488bf06148c76fbcc7e42dbb988711b2c5cc90daceaa83f0008e2cf41fb5e231c975b0a80489cdd6a3c2d9e845cda6b98f8df552d8827cf235195d6f54795d0030197cf0c7b60d4c822cbc37f4c75b694862741875b1bb5ae740283f9221decf2d441861278086092ebc9955990f63605a0c478c5846cb86d968c87c6cb39e3c7274f77c502b27265f61827762f41fc6bcb20997939ee41e42b06a08b77c09d832b6ee7bc386cb618b0edaefca470db9e673ff32eeed85649c1d32cdf74a9f8ac10ce4a3347d8887c49bbc6ac2fc9930effa0196a6d40ea5f88f1d8b53f55f61d9c8dde2c393579338caf7b6b508da4d07c0401109e0a49aacc9d55f741d048cf61217cd5f6802faadf6d884e876f9ffafdbf0d014c49fc35352d04f7684e5709ce02e08adab735ebae6e419b7a98b347152a655329882fd1da43132dbf7741c8df9d320a2e82e3db42c3984ded7b4864729b188bac3dcea331cbefc09f62e06e7b818146db63573e23d074fc6719badf3346176a22034a8a5384c6aba04c2d93e405df6bc4d1d8012298c920f6f215473de5cd4aefab416c6414d00eca7fdb935f5b4f6a83ef0bf1a773b643967856a3c5e4802d3642f30a7a63d06e0dd54ca2c82930e25c193ac6530260bd0fb18d36eaa6d3ed6f5d35db4387952264f26d5a20254e2cfc0cc7b0b99df75d0b8a716f351dcdaa2e83ab87abbc7d088fb85a855a74155f91d394ce2467fcd381814236cfca2a8ee1efedf7de8c72af788ce485d38a32aa8d5b8cdab2ca388330218c618e256e02555d2427b061b329d763437f12d563891f9c90fb9c53bea060c99e6d1e1fd2e21f597a1ebfe81b2727071e210113ad807e5bb6d766e732776113fb10951c0801b0a2f594045affc8c0c768118b2240f3d2882752af52d29ec5bf4a5df6e0530ae2a86d1274d8eb0098f0057a99f2c5d4975a23462d0df411838b00a9dc75fe9480306349bb2329503a2c3561b61e46231785022589abdb667cd933bcd4158b2889bfa22fd4786bdf6f3af7681b5e8bee73ece698f41986d1b49de58c7f28223f4a12c43d4091b21aa1bc8c62ee4279059b506385acf8159c909aa03e0621cefa3982a767c432c95bcac046e7f5ce7981f476d8593797dce8b693caefbb7c71e5debae22aa1663ca2b387e8ea5297d6b245ca7e4f890d90d268cfa91b7dd8d75af7ad7b270c659424a47e71db349d05f369c8b590e0304d7380e92052f3af5079d323f4db6ce941ff671726d760634a14ceb23199acc0e0a6feba10eb4c750771f45b94bb583886fbe291c084149b7398cd043a7aafd8fd245c47f0ff2036c83eb27fa77ea4d0276525ba9bc7d76e121c388fc747ccfaccf2ccf9e57eb107a645ff18f2d7fcbadca348590ee79e58e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1584e398fc02746b1c8cea6ef19520bbfd91d3f19b377102aac40bfdd209f7f4002eb89cf7a5435db00191478946eaa06d08a4fd7014ae818082d2fd65bbb8f0e78c93d6d60c479bf8c4ffdfc9084d0ecf3f1c4730245478d93bce8f50028fbc1d3938d9be2d9a98a9c9f6172230057a02664411d9c4df8a42d9ee016fd0084f5110d2f50d19f9632a52fdfdb3d0d262e16cfdd6b40934201f624d8fe3628a6bf19c5e214f203d57b0a22e8c7f1ba52ed2790401bd4eb99f99df1f665054e092f6bea3e7398fb9199a902f25d604c95941ab451fadedcca3b62a97e6a8d4d169045aacdfa935ed0c907ddb0cf33b190cdd8c8e138dfe136465e999b0347b6af6450f28e6192e7432ae66943d43370d56d3111d8d5285cf229bfaec4be4905bc24835e286e53e59a4e4a5455f27e3ba009b2384e496e96c2b4b171f29c4ccd5734945730628ce7e6c41b14646b4882fcc0ee2743380e8a19e13ae89b277b85ab8444c9724134bf52ab05b2dd46d7fc4eadfbee8ecd1607990bead0f8b6d8c5a129c2e3481b905749de7f343eae8848b378790376d89bb64d5b06f6725881f53afd7ed528001217aea3ed41ad5c91e20a512278215dfc4ab9d74e7285d06b29cecbf7ab51f03d9d6e0ebe27a0bed0519e9f69e66c894237b6cea564a13eb903f8da6347729116b6b641df05f3c013767fa9975fb72c88efe4893cffb7568cfabdc44935397c7e5da53d15aeca298f102315f0ca1cf891090ec4251fd6ef44c7e23a6a822fc714455dc51344190a39c7299013ec0d1bae06899ebd52d2e9e0be7639b6e2cf0dcfa672d42de86a03b2e867a5049765f74e1480accf0a33aa543df8f91641635ec1b72d3b97b3abe2c5bacc68b2078543aa7620964c80ea7a32a22b241a1998da5246cb0536f3d3e10756ac589d2d5ca1a6c9168ab8aaf99f502320541b1e3201b0958c4da4e9c32daef35322a03d02fc5661f707357d0bc02b7621b187847a58be4e242a8d5e1ab0f67bb6d50649f6f17a5dbb992f4d8a38aa698d46a9cbbefcf68e5e2fae2e7a478292d2aa99daf5362f41bc479a7a78239296b03ff3f618a5d62a27ad440beb015748b344b421b22e1701c3fe3afbf6da5c13091b0c986235a732509d6610dae4861646db16e672664ad8eaedcd304297031d9e49f6f0fa76793239409743120acac23cce6d52dfb01146a642ce078225f8ad8a45e2bc3dcdf719bbc81d3425160e888f602f9625978b6cbfe136ed50fb19fb4944018720f47fae916e24af46a5cd4cbdec96a1e43589f397794f0d0a924b19ef8fc7efd3162c6ca38458eeca72c0b76132cac61d449365c775acdff814c37739ee68c65fe917492db4fbffead013ae3b9956b0101839727d868728df209fdf62ba13be81e11b7468d6580834a5aa6f0a4363c122e09f4bba02ccc2f80e55594b41cc34419c5dd3b026b2b91f11fd64904894cd876ffe0ce8aaa6930acda2d2a271102433e4a40b02802598a5fd22441f81fe876067c36de2f47d624f13ea2d10197be683b1e31ba86db39ed6cc81ee8928eaf5d5fdef93538a5eb9e65f451acce0f436df87ff424cd9bab5806d8ac83a7f46a261a6828da29bfbef5c74a9b814371205821d09a32e8a3ed181b6e5a6f92fd5b6d93b018b32191377e3051f7da92622020a7751e185b3dc7440b901dbcff042cdb9597ea5fd20e49403c0738229aadc9756b680d1c6c91d000a73768db069ff3449332221bd9dfd55a8d179d571ca1cae8bbe7c3599d06778ac2e5d4329536cf7888caf2b1e6d0e8f5fd16b365e6155dc88214378b04353790c79e11a11943bde35b42c70ef041312b3720a343a2944beaf22692da3fdf890fa8372f394cede4f11f1a1033260e0b714644cad08900441baa308076e3a6271e48586bac65d35033fe1f9a8d4a8fcf8f5a04b78e42cc4d12791b8bb701d7c4c9f4230e8f5cd4a84324b318043e694a2cea25ca79c6613d5334ee1b0ab6b7ced6023a2728937309d1e0e0314f1d2d7dc96adf60e4f5e56c192cc434d1eec6ecf3efc570a9f1a8e413084e5e4ac4ab7b87f5bfa2db1feff6f38a68729552bf11fa644d524206ce0bf72455af66830e64ebcf1557d403179873f319ff4815db7a276bb1681e3306bdf029bedc7f661ce3df75a296176c99f0d6893383b98efc67d5e4b4ba663aadc8a64d6874f806e24a743976ebad8139ed39da0e0a5d99c6a8f0b0c3b2a576c123c2176f9bdc507efa691ad61942e6bef2d0556c6508380f17b6efbde9ddfe1454307ee0d5f1d0850bdb0423ffe15777e6a022db4392fafe207a18b8bbc2f6176f46a85927a9872d467469c42b0c9d3da13197f6edf02948bfe59870730c81570f4cccdeabc06b3c2693809aa30d782d54a36c8ff87ce5c845b2b92d08d4472095c1312c5746179771040d8e16bbc56c33820c044a801a5d82f5ee08c5c79d84c014713e0075a2b0d790bca4171ea5b60827e28b78dd1b9e160c39997f0cee0e295757c9222f93bbf817d0fb53c900dd405fa9af2c85e39ec733ee4b6bd28a356876b261681d7b9251a63d4893df4176fa688fe70c326e26395c691771a0ea37a2ada47346e73604f2b0e6fee39f137e3cd5968f55cef96ce920e30b1c0e3a4828db4a3cab00f000ade233ed5fe617c55a8fb140a59825053db7f74d4ac241b295694fb2325b187f7e630885d779365fc8afd0974174f768a913378abe1b1e0884ad0234f7d30a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3f6a80d251b73d1592ef4c6df86498ae9c76534f9c149f792cc131096a59ae96c719bb2e1aa0e8858e114fb2c28b7c1e8efcb8b527960e185c3bcae3dbf600afb1b272a7881af565328f4130ba9639b989d79339029836831832dd2b1354a740848b593cfab8e7fc03f01cb6f439326b261eb72c0bc8fa8a88a2356a2a1b7818cece3fe4b82faa9e363840e7cc18d8d4c3c4fe41d5cc144f908b99003386f62ad52397289565466f246e9f1b6e5bbb28cff1aaab5e4e8c60b8c7e8e6a1cd2951ee0e58d55be0d3e1d08ac1d397ed4619d986c8f5b479289cb605738c45ba4819b41d709e2bb33f64c64dd7b935d8e063ee177aab1185c70dfe783f6b5b21d49bf7ba049632f1b70d0b978f5a1b64662bc949c81a8d1f3581e8e70a18af72abb80939b215cf3c6f18c5429be9d7e121a2fd8bedfde060ddaecc5a233cc1ca92d7a3adbadf020defd59107840d444a34e270b213e46ab259ccfbf44e92db0236b3fed1218459bbba273ca52d8d17f29007ea6d67aef82bc743fd367c4a4c5e0b4db960be3c4213d44a561a4c2e20484113a6afc41af6fbab6f7d04c34d2247bf0128efbdc4aa674138a82fcae59a8f83e2669fb212e58ce66b14ef6e92d256210f88a43e08f9141c172fd864f6e394c26b119dddf81f912d50cc9cb800534df6f45d371c1eec1aef53622357bf0ca09e15a30d53c41525868baf2b53f2c493cc178f83078ff41588a0603dbf0fa2b272ee71d2dee7258ab19a7b7c99415a9d0cefbddf67e365b7fd9d7f5b2fa935cc5bcf004d4a967d62c38a4260e00850340ae77765a4fb3ce157fbd40e149187e2feec42583075a22563e5fb0c99d4354ee45285450f5a01db50901d03f872075aa4cae6112a5ef476ac66ee05796f22a5b894cf0fb80431059108efcbbe721b9c4294d186f2880a3c9c2bbade937225d1d383ef225d0c8c4eafcbc47115f99c703eada245569311c76fbf19faf7699268797038c2fd903d88e682c324418670c98659c935316396a3f95eca4d0ed32b1588b7a07a795568300836b1d330256ff3e11e1632ab43fbe433c15c82d9ed8a3a4d993dcbba258feaa10ebe01a047b75ed942e9f669223e77ce5a7e6954829403d3eefa4aa24e6bb7710503855921878cece8f1c05aa0a37c70e003804276c43c0b24c2893ba574918179fc07fcf99879c1c5d24053531578c321e3586a74286dbba212f85ef7562b0482df6f6ca543677d9134b81caf00bf6867519d324d4a9354d8c0e43375420a7a07f6ab11deffe63593d8267af7924033e84e6250d966b3fd78876492f5cbd002a92dc4474121eb7a0ef211de60b8832cdd7305cd2c25d11218012d34e616b5448ae61d3433d39ebf532937f9cd248af6c1c82f82ff8c609a1ad1619c2df6e47d5db6d84256a1c71894441eb6e9ceece24395b27c2cdd3a9fba952d1f438c04df77bd012b3c1d2fa3bade67c8c6139d149e7d58e049ec81c44e527adfbf9c1d911801a7b33010fc1f0bfa54e4773dd4cc7359e092d51fac8687f735885f38c2b368232169943d606caac7f746b14944ce2ec5f1830eee654a977917663b85832e1154b15bf6d301f73bc77dc30f35e813c95ec7509918d7ea2bb765c44406e1764764e30fdb4c7f0e664dfaa10c3fe813de3959e8de40ee67c48e48bfd6ff13f32bc6fdfe66d5090c2701e408df73edd2bce74be572ee3fa7febae8d65c09e9ba146f635a17964d480c7e973ec39b6f1ec5bd2f73dd9b2054fa3f3d72864dce7ef6a5942ce63f4ad5ef925b19e26d91b6f5e0c2db7e68d1a0044e75fc3575ccb4b7dc8c44da7d3932f4db7f4e5cd05e625d4dc380b98d1933017921764dba144a90cfa030f180ae8cbaed8c2a018795b263bccfa6493df602253a4dea0ccd076a9f6f0a343b408df82ac0f85e55a3e5d72568f967bfc63e7ac9ba640d83ef097b35c7ed5d6cf4d6ffb2ea7c83f97548fb389bf580f8d717cfd9723e6e3dab50d2773abe54ca7edf45e75821def1ef1b49e24633d87f0f0384adec61abf199812f353fc9a7e7daaf2dd5fa5a912ab585984fa9cbc18d47bdd910106f780aab6864050348a255be5e29a1bd15261e9f70803829323bd7cde75e1a7cc6c9c50df61437aa8a5311d84ad72408f8b576cfc56cb3c6797ac93a927015cf0184e8fd11edd4958d6be9b2449281af07f1061cfe7b824e84a7ae50d79a134b5bb966889b57b402489ecf815f18960e86e0c7f46aca1f18c941ed4a75a4e81addc7d8130e1f6815d2ed230d205585cde853ec81773434968e17717a96cbd672a1003aa6fff195359c2fb092c3c6516399ed98dc928530b3fe1013e07ed743be8248b15a4439217e81b5f2b4fbd2d0f97f91a6ab10fceff520525e51773bb1f1905abb035a16e5bf2520739d0efa828a12b184e33eaaaf45d9e9cb15b7fde138223a61c9edaef929948e392a781ce54f9c0f8ba7516027fd33de98e5456415dec2d9b39a41436e6625bd6a1d20847c09a2c7f8b41e57c190b0dee9c2d15a6d32346e448006ca71040a47a8250f27f427480be6627f9588195d492b4cddfa586536831559b23e317fbf9c8086e71e27070a27b8acd3309d5101cf546f42e7aece6325d87240acd6fc104c0a6a73e5325798eb74d59aa801d83a9ccef9bf81e51e471113326ab441901607eab11b3440cec4f062d97cb18130928902da1a6f7ef4b2b91930657bccffbb63c79c6c1bca5dcfe0c86f213bb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h64e9c215de01f8ce78d7ee538a7bcac17b8a39b610d4017d3c74aa105ac8d99e6044c5fba16df4bc0803d4e0fbddf9bf34d8e57d75c80cab075404c712e5e5fec560d7c35e87b936f27a383360e9258056b577617144581f2cb25a2ffdccd2a31189110071a54bb65022dc4b30bb856b9c2707c28a95341cca31917f01c06a5d18acc9853ef60fa35da57aa8307707351513fa087eeee3b07af62bd656993801c319af3006469242ebc7fa86f4b4890738604983e24cdaab023f6dc70f760722c3656297465fedfe1116e00d0af0ada88e5385c8de714ecda556128e62518518e965659912d28b6c181b0aa2020d11c89d984fd345d6ed1b01933e49d711de657fb428bdbf1ee7e429f8033bb86f9429238c391fceb4deb632cdc785e728e6137df13609b50eb63253a3c752851a9581d125dd3d923461ad01cf552e5a305b3f7491d8b17c5967458364191c217fa2610ec789ff69feb4a23ad52cd337ab334511a197225f0a724312a91953c1cd3152e9be94bb230e477d347abefc188a79ca0a3e2a05030e1b6812ce508ec648b09debac249d8f830bff495a29ccc35dac4742a040c4ef3fcc478b33a2b2a195cf66d360d34eba50a5b2348690098fe267e46103de1ce55f5271923f670fc472ce3829a88058abbb8bc9b2f6fdd76fa184a9ee197990bc97e5b3432d5a8d0cc0c85f6967bfb855eb740f2f123a6d2027839f3516ebc564ee58fe87170941bd128a4d9bf8638556569f3418e6a1d4c2ce8d312e42105619a41631cd3ed16e3764c0481883e4d402d710baa9a4fce61d1bfb4edbb0a044e5efceda4eb29b7af192ce8798421eb440faa13889ad3439e36f3b08e27369714a19029e902f443ded0ec395e8b258f9b65585d222005bf2fb067a0de6a46d77c39f2f2ed094f78e6c48d930353b8f353bb008138b45742ba9c2bae236fbcf8af976c9185d86fa7e40e67d83e52c2ca9aa167eb2e3effe2bfba0b18d586fc4a609cb4b3eb86aa5a744ce8d18dfef2df1262c280055e5e57ba5b86849239e7e8a7b04fcac360dc83cb67ce304d0a42d6f5ef53abe46b72fa0f4ad0c2b0eacc2308218110a9534609b0333dfb76850f6d3e9eda92d71276c22ebce7066980d06241a0459a2adc2c6aba4dc6eff413e16292e8d25e96d012d9b030bbd01899f5185e5565e9c2268601d918896cc02c7f132f05f0539f4b5e3f800ceb3ae7e4c52300285a6d63dba9136337f2017f51a56dd2e8b8d11f592e5a7170ab9bb5f7576b39d3dcc6f48465cf99436aa2153c9c08dd6af6032c4b8df2fad97a833c934b8a5c140c915eba8c233e394711ee067585f21677fb9dd93daa66f0b2e71e55e01716d38fd5e5c7f37d1e00fbc14008b3f46399a6c9be47ec6626656537df58b4d51ab46366c5c34daca325a589e8215c9bec15f5ad4d8ae74deba7475625d90678ff3dd90a68877b88bd50b2dc78bd885cd8723127259695dea0e6b4357b971c3791ce62f199b50884f27f887d87d88804102835cf9283d9e99feb3b020a6da1875331befaed390eda23e90058f710be5b6aefea0d6d25c8b3b6f1e2e75928d176ef91ba6f25e83d8674175e0f69fbad44c00cf4ffdb8a09520c1a604b359a38e6c9ab9f90fa64ed58cb299b5d1ed6f3e8cc218e523ccc38f47c94004c464da20bbcbf72849ca6cd8973fe6c2cfc77151c33bbb95e182e5e61a72e243a4d7ed2e24e6036d0c9c9d2b410f700e6436ccbd64050cc8b9e55e75cd24bbcbe000a4df99da5b8f650b7f824e37451b740f2b870090e467b3a5f435e94c42a63bebbdf7a47fc3fdf293c1493b8f3ace9b77fb2b3bc03a4e2b68bfea532e3208c18e6797b818c18c1c69be52491817c57f29bbe1fc0e0a68263ac5c168d2e49fa671586508ff9392ffb6b075b1621be2e9c10c421706e6d8802fafa0b401e9757670c9a9e9f92246cb56a3e39353121e9f527d68fb54a0c05015db0021dd24cd8e2aae0aebc14ecefc9c8bdfcac71e0fdede0a5dc199ef765a016be5c9800fe5c013527b3fcd800ad2a5318d78d2134442756b07aeabbb2d611db88786a776f4c6d785a35867afdf94baeffefd0a7be0c08eb02ff5ae8c30983546428f68f0eff09b609447fec9173d20f3f860c6d6d1d60083234e142123c60c38dc6da03cda2a7aaab1ffa5a4a95f9513d2fe3cab04d60c5236238ef453baa1d70fa54d2d69aa36b208f9d5fd709c56637772865b73182fe1390a2959c327f2bfa21a7daec3ba3c6ec2a37f9f52fc6c64a1e572f300e5919f1aa91bc0cf4c215b016aa34df163157d6315baea2bd6cefea38085391dbe1d6e159d3c77af1e769e2961e1e99dbd8495e2ca75416fb080ef7d91ef3f6f16be80dc2feb6fcf88e57d616535deb18127e1e7a494aecd7dceb32b95e7e93b1b15608314927e57b1dbb8a5625f97cb3f70e76dd4a44fe148645005bdd076c7bb9ca7fd5bd9e1ed7444a5164d0192f4d4f51cba95247e25880c6d9dc1b428a039ce7fe179fe66b5b3068694416f835d0ec79f074601c2b5c385a5f2afdad252a73ee21572b00a46e9ae39a1d4beec1453a004ee8fe28a7e9c3b81a140751ad8af088bc9c81ada7ba551e1865191b3b44788c67f2370e6adf695ad0be004b86f72ab9c429bde5bb2085c407b554f40f259742a80d65092ee7b0a36ae34bf23cc6f2b5d0e6b95906f66335603d5a1d2e8a516975c388f0acfb944fc8453ad3c373567e3bea9edf30ecd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3ab90130805dd50520455758835b208bdfd6f60072ed75266048a3c92b70afcc98152268da2a03a7746e0e62f1b98333ebf4bb1c4a6c969221f5c9eb6af469201433d956d04d33efe6c488243db7a282d79e69dd802f5d958bfa33d7a77e6ec641572e0c57f63a3db438e5d14a295c89b44b45f4484ea2b6ebf1836ba83a025de30e8fd26e7f6fabca38a33e08926a0533dcecf150f53e6e36ae1dc6e12d1683c385a1bfd706b36a18a70ec7a12384aadad729e9ebd7f45730bebec1a8dcd6e07c968b25131247836417e84c2c339286f44ddea95319ed35370c76bbf2e6a626e3ed4f0aa332a926389655b1dcbdcc8c3167540d78e495be7c66e8fe4aa6310c3b43441e88e22da847b0968153b9d7443b24c5bf09dd9b28f85c48158224489e5ad33f7811af098086c22b66cb968dbec4426b6306c1711cb04ef2c3a5b5a346bd486fe50133b94384621e8131c87caee4ab7dc4f7bdc73a014713b87d690bd77688aa99ca4aed27f5ac80722ad9d929a45f5f1ebaaf3f1c9e38a23f5e67024fff8c9382ae275907ee77c1db321b49e304acfa6f6222808d2192bf70d2876b42639025c96f17b9cfd730a815cd7a004df8647ce80edffd138395fa9db1db3e43f7ee89cbb1064594618a7293086f8313adf9b87ca4f12a34df7fefc5be58bb303954d7bb07ab026947bb4a3c2a1a0c26564a2c6a1c8e9416a50c2eced9816a3f20f6c6aead758bb0b60901b107c21417a0607332e518e30a529f68e8657a0f5cb85322e901fba7187902635d5481626b1023881d8748e8c1c1dc6f8e39a47edf3e58dfc339dbce6b24a00537c8729583f9f569871406617d38ec79742f49dfee8c1626d3fb1a6e35305113251369b661ec2214a723e849837dfc164c40c51ebbb192646546b90aead3db426d1c95bc563dd6f6833ba6ce8707eb2bcabdf81fc2264f001ca3947c159c1f5e47cf1e732b530a259a7f9fe3a2d7d8d4c5f031265c5b0bb3582b1ffe17d7425d7631bc829994efcfb1b4ae7b4779617f811f20e54c680166a1d906fbd2bc0d114dab7649a18909100ae55adc495c240426bec9d59605135afc1906f123b0e77b7a53ece616282c60c4cceb0371f3ebd0b5ebfcc2e74e2106baefb154cef95b1581289bae95a386ad6b3080bb351414307b34048be69ef484581e5245513a5244bb00ff53df838598e064ecd3e9efe080035d119dd894c962a6505d9809060eb29027fdefa1b0bd632e8984bdd991ac2efce4d924934aa02b4c187cbdbc4b83463938fca88b8083c91e21eddb2baef709682d85d3a7a55fe90d32c3ddecc3d0bea91e4ab5e26dda4882c8e050aa09a0dc8410f165c6ac6f6358aa6f74a4c83841f36224e02c324d8763b10e204d09ffe67ba572514c75e9504e20a66c396ccb9a0440ffe4c07504386cfe2ade4082e2d263dbbd76bdccfb9d24f43f136538074a9b8459af54b16d528d1f14853aef90dcd104a54617ecacc3eadad5f1b073ce0cc945b0b165b9705d51661d19f72a2115f6a0eabae342a98e0debaba5ccf4de5dfac14f736cc226eef199447807265bf391ccc358e0fea6e5525fccd2cda1b86a7144ef42c721982503e3f6e14b67ca712c54142af209e0c09d2eaaa9f1aff62852448b3776f1a274a96787bca1fbf7aeb3967af45be74ef2605fb0ee43ccfc0040436b2d2ea923914e88851d74a29c3262406e27204125b5f2789cef9475c05e9cf21412237b9b9c5b2e8eba5f115207a5cc47d3bb763c28c34ac3a8b1b65a5b67c5f4ba384679a6f230ba7b0a3dfe073f00dea1c17744e2ea274edb226741982d8404f014d7339fe9a72a6ee95030fc1d8bd1ad5a07395a3b2a993bd31de68e834ff43b4385bff46dbffe13c1c21f3116e13d694515afd7f1ea92376b63c5c2f9ef70ce7ce70a5309d954bece6a4d64d615950e3a5aaca022b895ca05dc15d39c52e4ede2d0ec0099bdc04920efab65012cda0d93de7484bc40090b1eff9a07d6e9fabe767d8ca39ef1ef43c585557a2139d6720e3cdf4f17af4b6d1f2eb8bb6a75418cc529c604a3d52ea03cc99368fa09210fa71312256abd76933b4d40c0f6033f183c54c934759ca5485c4a0790c226779a7f11156317b4099280e5f916e659fb0be32fc329da960eb43427520a14c9ef1fb6a4f54bd672f5233c6c582bd6ab543f521f6a698dbdd62de82399988e112b687386884d8bef5e2f3fe41e633562d6c91569ab109560852b9b5207ebf8f5b694d7125fe0af0e0e353413321b32bd5f891523fc7c1669e6639e55a0ccc5b235e1abc8b42504d53baa9444f9c1ef22b5e2691480ec7bc19fe80cd94c56c508c26f131ec4f4fc7cc6e920bed6703e9f988e0e83451ba52e7ca406a71b66169137dfcb624d740ad1976b86036e1dc5d4d249293a86d3cef2041e18cf7d539b5415bca5aac24830a23cbd9ee37e90f7fb4bc65317aeaee6707854a527a86be76ca0041bf188c00c1dd84be64b4721a7ca1e6533af21d141cac945d5cbe4efeb887a68fe06fb1e5657527c03cf0e9c47f3fb622f01c2cb8a15368e8e6983e07e0d1e8f4a03d911a103ac8f0365471e939c912062a56ef3b1e9c198c760159b93649c78bf7af01d73127b5d5413886efe120dc5069f60ec606363534246a7a1fd11cd47b454f06e9cf081cf5594d2d83f2903659ef711144ff311ffe6201d0406cdf0610ab611d58db1b5395e418e204847a81d539d26265b04decc58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9d7c8ce081a45a68b05fb1a9432e6bdcef1478b668bb8d6373e231d6d10e487df147fd5b06da7706d7a8a54607af459967e37c18b861fc38022e3a52d915852eaf8bb781e469b61470625758a4c0f33c48452c2cb4d8d85379d6f68b53ef929da5dda0258e4c9d8dedbb6b07a46c72acdcaa945e1e0523bac26def0383968537c88648270e6582c070f6f0d2eb512a5e0a5f763bcdbe16adad87483edca7b2ecb26efc670dd8eb47d0ffacbb42b389f1cb65f75255e71033af34254c5e047a7d7800caa6d8d71d428ebaab4958b60b84a90f859061955bf6873cb607733496f3f88794104b89cf301e7de0b28f6b8d92418333ce2bfe78f033618cab63499246b51f0d0a75bb9750901385171a893de0470e323ef4f727f8f407abec5ff8013413f60bce4ae6524a983951a61132185dfbdd0d0cde581e945f3c0f51e4d07ae62ca0a2a626c27672065368a04c87fb87a167be2a10c9e6e9a96167427f5f95ff00c6447483298e1e4781ee4ef95c365fdfa0c75b8b83ef3e2e61ee88ffbce68a4c6bc37806e2a32d8b9083819b6e40c5bd043994abbe713e8a4ee4962e0c54bbce59bbabf59d9fa829467700a7a24e4f8b39d44e4c5c1b3343e217acf17511890e38a050cffa440d74d455795c4bbc3d8dfe1ccec7c37c765c966604e5457b8d889f3a725e95be6b3b2148c7f689d518f01fe124de747e4508d8ece8937a5bd68ffcc9ea3932a7021b909678b65f5c4ab255f20ab24bbc5d95fcbc35adbd72f37c96c2b0246eee89772fd8eef949eeb7ca33052e33827378a88503508e58ca5bea2dd9650a86aa29900e01584f277a67db3c0a0484f598020c97806a4a6be81040dda94f860ccfd5dd7a24ba950f31a40cfbeaa0b708465c3174a06f438636139a55283c91e08139b6f58b5a602c08d15efcf969104d7db3aeece567b8467796ec7f0144acc4bb808c20ef752bba83d62bbddc5413746b4285e102be8368b57c4ca83b5dceb5d650ff9044a5295a9d6d92f7de744259d35b09c5dd7f489f653fbe7ed1e4dba2f4f8977a8b8c47e4be92ad952a24ba85d3c705aeb0f1a4018ab44f9d882962607267241a576da0dc5cdf5ec23a71cddfe8e69b8f7211d169bdcca9467e9aaf70caadbf2e49d16156cc951ca310a2fb1b12b313b4ee213915c7861fe7920a690107e43bbd51c91e68f1c6b10a094077b1778738fb3d5b04c457636962ab6622f52384e93713fe0f28ed3d20cdc9fd3a74ab9f000d12f8a9c3cfac98af66a47e8692b99010c34909fa32ffcb2717b23059ca6620b96d1520baa81770e65e74ea32641ef82e82a7e046a4711f9ab418c3a7838a76cc9a87a57d9bc226fff4a17a196e38b513ac78ace21579d1188ff125c374a19aa7fc717a20abeb4a28bb138be177160860f6f26c9696377a84a954e53503e08850d8da4a1965c0992f7bc7da1e7007505784993c4ab013aa1468ed74fcc839bee8f30f00563815a2dac2166c0f6405132ecd6fd8a085d02144fb41de2a67944032f3aae44ffc14d12103345a2729ede70ad1353fadb8142c1dd7306b68c9d3130fa09dec831dd7fad56a69f3e81e2c236b76f658a07dc576fae35d29c6363d4a1b09b16c71c95c9c53fdfeb2e0be659981d4f8f043da44c3ae908dcd51526c1400e0db1c82d3d17e15eec3dc48e6c01eb34bd58512f38c63e9bd62bd448167aeede65a7025d3b24affbf1dca8a2b01184fa58f56e17afc5f8babafd03fb53b259bd2260b3b537da715e8c28b4fba0b6a10573e50ad359ce15d8392affc6a7dea3f4cdd19819a854ed6b68a4420a57b27350d4b2caffaad0ca9c958ced835f47e70e9f3b74c6ffcd1aa7a72c29da0d413189783ac3be29b1bfaf3a7e86723f66034dff1829eba96298fd089363b2c912a521f4813db4cb2843560f68ac332ae52768d4467f288d2618180caf2acf56e15c7f304f60cf65bdfd7c4c7df59225d6fc724ea04518395c9b3270b39a22b25a57db848432f43b7f57916d28c2c62436720cd1841ec96220e410f67d03caa3388dbf3cf701ed248ccc787f9a5661813fb2322728e09b255377748ee8cd403cee108c52e20374f177d824dbeef00cf1d11f5b92deeeb6883b9564378550242a9ec9156dc20a31c2b2a3a547c96ffab0533cf9e3e030f08342563e06668f9bae20ab5c8b49f24007928fc4f2020decaafdab110c5df11905830189f4c5d1e10f0a4ad07f130a1a86ef9de9adf49e186f3cccb84d9c5fd2bda0a319da49f7b8ce93b83439397bf463e0ef9ce4a8a9eab97090c74d3f875932be095897a8db8e8406f2d41a8102d3c646b0678a03340ea750a54757d49b7ef7ee3475baf7290fd76bd25f7e3dfa189d5eda6612579a8ad3574ce854d2ded8cbb8be7eaf78b24b2b395af44f8dbca7abd1c4d640c49f699636ae6dca9d34bd3b490ff48c71c06b6e69c801e8c2eb1c55baa73cd28dfab9ec02ceb20425604025255da8d7c7f4b4e4b6c97922cbf68af345e61216665e3f59ad2ea4d00f5936add45f3b368e8b8d86f4c712174bdc712a7880dc87429c251166dc873302fadc83049ac3629009fedd3e4de93703c09e151246a103b2acfb64c47a0c878c7a76374fdf246e5a4a88ab69b9625099d293d7d9d4fe8ac914683e862b8ed6123aeff80db014e0ae1be9357fd7c4d9af4b5e848d8b1bc427a7cc21520c21b68ce6153cf03e4eb1312b42e575c02fa1ac661724023017c344819765a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9c9bf311320ff290cbe40d4a939bb63459d184fc05e0f50ac2f85662020412dc3a5976e5a8f8c04df8d941558653a66fcf2e92faeb3341ce511c83e3144632481b96c524f403af79f60597e481150d9ba603ec08bc6525ae89badd349a8e74e05f89803b857ec98ee8aebd2c2a0482c3ba3e4e2b605e8062650b399eabfae6ef0bbd846d42fa500482b41e1ec28926b5b2713404827c433e80ef3a073400d9045e6ea7f674ec3d3c1766e358c7cc4c0319133409ede9435393c8a18bf1216cec321e8caf0c72264e47147239af77d9553db06a80700a6933d3dff9b6728c591bac9de37813454c53a3bd7822487511bfd7419b27ccd3dc4fab4719e7523a4b1deae3b228997184ed9e3291575785112fdfa466159503a5a3faad5e3c95b3528de69fd0e09a698f6ee162aa6f4692fbfb26909dd1dcf833c5cd85ef1c096442fcfd22eb15c2be6e63359930f95beaa4fbafec40a9f1015598a11c6a40adf76f267d190add089cb728f50d430d190108850f31239dca9a39d898b1d4cdcc14abc998d97f2d5ad08ca9c2970e723a4cf178bd6849203ffd20b6d7f5156c9fce15e6ecbb36302878ff84eb7a3d66b7488b7427c6068e7768486cfb6b0261addb39bb3ab9ce02c89d41202159aeedfb1b0857e3b5531afc663009e4196b8e965c65ea4a7f829d3dcccf0c988ac69ee9487194df6de4a82bf56f440457a57c28f04642652da0c43c6905bcfd94990fff48adc3e4e3d9d8b9d7b3b09d5ac461416bfff201f454020a58fb1458e78d4f310d5eea49b399f459be17d5a5c62e39b2c1ff2154b45043dc496b68a2b9899fb3139abb7f4ead687f409dee6bc513caa85ff09e3c6815c0b74c38bafd71079caee17e3d361b460e8501b7e51cbf994b93cea04577016f211b27841581bcf7628fa2983da71073fa49d3dde58e87b029b56c24b48e63cbb2cd186513f0c5dad3fb7576f1afd45e76ca560d875c565dc96d277a645246340b68cea1884be744d9bb899e2d65dfce8aef7caa695ad248e81d50e63801d97c8986172f4ecf0d5c65828127dc496f6be256108c733f27c91f5c98efdf1a203b4dc9f671420123a66a60bddbc0bd3801d7888612bcc0cc67866f209f21703354cefe61b49368667b675ffe8375379a80316bec29c17d5e33e872afe65da2d11779662cec74516f3321e89a0ec43b7d1ba03616ca9aa713fec16dd4a97464a7d34f5513988b0779601d48b6b7aa5600f514b2fe10d4ce4ea977227fc0d266b4d8496e917a7f9d6a32dafcd015c019f4ef277b457ff98fb995473aafba3bb087839fb2a4a28d37333a37d199112bb029b23d2e95c7e24e2b49264945688ceca9243e8539d3c4d72e0a1e0ed640c8d9ed13e0b609f7151473bb71222e8905cb8668194d6eb69890268cfa11891caf3db6c55cca0aaa7ffef15e5abf90d8e2a8c5b3dd55edb2808122815a54c3ef16a903fbab988343ed4b6dd919a3fbd7fb70b90d802266f2c6d3e5c3aebf65b64ff7abb253dba49d88e29d620a07fade974d4b0e94b051076aeff294d45250020833174c9fdd471704016008ecfcfd7f7a63ac1fa095430115620634aaf20048b8360a6dbfeb7a7de68e33225a198aee351ca241db95f355fa214623c01e2f60f72ae5a4f01979870838a650871c9268d4af11005df674196c5bf40074b83f8438dfd279d2f4789c7370044d3954ddd34335628456e36904553cc5a5740ce11733d04d464a4773211321be059c45cbeb472bc4a461b976f9e74e93d01177b7a9f12aee687136b3a44d6bc3d97c30e9175fa61d0888c936cbb8ed620a81e82b7377ae2fba5f651350c516cdac68bde7b83581497b23e129c308f9ea05289033921de2868dadd456bf33483c4e80089ac80b103fbb11bfbeca384a24f77c59341324300cac73f429d9441529e49b2df26631ad40651fccedf81d0309aa9ce74b66162df41d0bf63834743040ad5f107fee58ca65a96aca3cf5fcf2516cea93551543482a33e65488be9a1a93640067e211d94517a10f69153468d4a559c24a618059bd57c52c122a230eda96e2330bda4ab5cd2a3b34a8a4eace106d5931b5f3f77ca1c850e3f99f2940c7ef3e7b97e1f0f2fc20b210ab1fc3a72ac0fc50541c0f615da68b670222304daee24d5ed62d37b0342ab27af1eb84339713d74a7f7ac41c0b4f9c66526359e9f83c09f7fff8d30c4b1e87cde5e3144096bf5214b951ad662128cf47d07766313516a3cbc0aaaacf85ec93f30db6215808468725ce3a471ed868a0845a890adf28ba67fab17277034be2c30ff819cff3b60cce941a4f453398e49b42b37135f007804a96eeda6eff95ab7a758576a57c437fe0f1dcf4fcbd9f53455bda017d09e9a08d44136924afd156d1ff664c85916ed1fe05ef3ea6f8f63e968254fa0bae9d8006c859f4679705d76a893de33b6b0e282d22c643ea88cff626e99829c70a3e922aaac5fd44508245f8c297b9dcef956383101238e8d212c43fd1a2bae426d5b464543810cf1fcef87f710f4512149abd998ee8fb6061fd3fc9c3da0442f41f3c7bdc3d0f0c7d21a1f42c20d61c4107ee28400ef862590e35545d8f1be6c2b75eef973d9258f59c008469b6fffdbb1bb4b9ece516acce8600a0be0548f47ba2c0144541162627c03fd40c3f8abce003d9cd8ab5c8ce95b80f6eae0252692b9db095300d858e1f0ee9de0b2a261552d592a1e59da1a7a1888fcbc34602137f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc6b43acc885208d1ca10eb0a8a9bb60cdf1b7a042a52f59689e198f6e305aefd0134c1a77e80f0b97e727eb047a416ca8afc9886aa05cdfcabcd43d9cfadedf94def8d31905341a635c1cd631a16a22c3863bc90f09c1c9422977d308f425beca10e5f1c9549e6eb20ade8ef6ac0f18af426f56c3812854bc9f459664d7bc48af703454b87afe9704f18537b321de8e580df9cd68ad292713f22d78e7f6caf4b32fde12e88992587575f3a8301a6f5477857773fb8764a0552d4f023deee9de27c5a42203a73788512558d299a40ff3986f1a61ab0c1e78503af63ae08a66cd87acd06923770b394b8a22da5295027f20d88e01ff4bb5ad1acd64e12f8782f270d6178f3aec4e9f97bdf183ae2f4c156428e80a34887975a3119cab16251fd07c0dc831925c404e0a22ca278b9cc6c4d2a90537cb9b9c285c0a08b4a5b94fcb144a2de11a7a3ae1e90fe72417cc7fe5ba51e8ac8b4858cd6b135f4ac94b05f925465d1bc30282f777dd0ef05f3ad8bdc5bbbf97e4318a987e57ec743bf026fea3e3c56395bac0f810430c70281f00461309385b9c7224b6a50ec2cc56cd8ec4f3a346caa75b9f5ba944201d3d8cbfbc11dd4eddf4534bf728bc00c357b078d0c732bb0695e7cbdbc592aac6990141ddb44a5a406de937a19aa72045338ec3c3ffdc1cbb0aff9e8e11c05bab89d45f00e05a9a785b811f0b3ec9e0667c120d169c9f7169fd1e19f6a95756e3c4c22b70b6f4ccfa1e9416682714df65a1c365b982b56d81aa243d9e84d05252ab10a71886c20fff21ea72bbb9ddbfb73da4ff74c8d60f0aed8cc560fa1f7f919c9ccad2eab8c444c174a8e7fe8d7503a5f7264a49c01547ea7a64bbc6f6ed4a9a988d7409398b4c76c2d3cf65de51ba09968610e644fc2fe4e1cc65133b5c9207caed23816c8ec4e98bb622921bac93ccf7842748444bcf25087d8b5c3b92a0e07ea7bb7d9f97f21b157c611e9113c74977db459897401ad6d75bc679a8c38ee17ade60244715fdea38859c958378e23a72ac66e8e30f01519c5f09f1f0a77b77dcfcb4e1e7d4e96991a41d1734b6b5a14e3ccdbd1d9f8cff8a0a883769604661902c0a993fa3abd59c0e92dcb820122936ed14dcb1664186407820131fe5c5fc4d42d030a5433c6d8a53a254a6070b838330bacc61c64fd73e4a094255c4507d173a4c3c14b500d743650e78da605ef85356abf37a809268e3a062ec96e3fa7aa2fad947be880c16e56dab3f60115d75e2ecb82bf5401a3a04f076198c75cb0c80b2e9ccaa3d165dc8c7e96d02501b70954ee5b4eee55ad191d3a24b4e6c3c41137be909cf27a987f85175ca34f1c4607003b2d7a5f603c95ee71454e182090a3325a22f1ed2b3df6d4848f41c08a1201cc773fa215ca241cfc71d1c57826b91eb6d1c2b8d0ccaaaacd15f826013f590f6e3e686f6d331c06b81638baaea448bac0aaae01b903d6a43aa24248b45b5916d2161d5737fe01f031216d8de99f75152adc16113012f049ab4b6709233ec108ba08f3ea9d7be47322c270cde065de2cc1f5b95a052274ddb06083320d0b941ff870c41a190941ad664bbe986bfd9e7a619c523346fec6b2d3f4a8b55fb8c635ad2853a85550e40712d730d4e07e35b892c16e9b19948295a69bd209d3915a9a1b70e47ba21bc78451fc7c9fc9029a7797606db687070f02c0903721e6bdff8b7b8c796ac8255f5f1ff32e76468e85d695d3668b7ee7479fad44fda55ddb3e7e8c3c2fc4b76366a21e515df0bb46bff6a935b4a41cee5713d59e44f66d779f7037d3b06e358f11bdaa0262c3565bfe9ba0c5013e428da1e8453b2234b21f9e6df0703a080baf43b15a90fe9945790691f0599884f2c56433edb7db33259dc423d1e11ae3f0ab01abd5370f26566e56594eab8ca594542e7f683809fe644e288ed8dfc1d986ffabe76bde66d9553e52ba27baf6ddd4ae1eb270852cfadf1d7bfcf829e411e13969c9f54f1547e1bb52bc453fedffaa095e59e2d3728958fa571c888d8566a1688abdafb43d4bf68cd51a97fe404e242acec45618ea5d1f64c36f7f4b886791909ca2c308a62b385a732c797ec442f4d3e35f2ef87aebd893b7d19392dc7bf42f85afa461c446502307daac7a6cb7b6d67bd16baaa0d002279c6d4fb95f26636e07c05d3a19b28f200f3376d3f58a952c02a6f0323c6e4e2e5b3afac9d117be681e6ba4bf2714b45ff4aa1eb263ed506847b377071692caf43ab7dbe9c5af909d4e7db7962d02a8943f681f9ff6470ab1a55950a48364db25d143ee5fdc75c435a3dc572ffdfedaf1a90df8f4e9a15e2a4a7288f532375d0014486033b2f4b66b739d6bd0ff0e26858542ecd8b347d9ff35f9ad6e81e338d4268c1826c32100bb8e5078dd1287889822d6712c071e0dbba8f1f143e6bcc19cbb51766936b5c0c2db64e0dfb074de8a3826689f4eb1e13c069a207f3e21ea934e7663be35b15c19c020f70fdc757e4707f8d4abc02edfe427458c7c69caf848ead0db16b27e04e77bcb765791c0d215245b3ff01cdbdea7d38b7823a39da4379eaf31d43451b7fa530634aeb1f9ec13dd982baceac61674551b820e08cc7464c0972840661e043826dc9d313bd11771e41cf6ae534e443e564b7862b8bde09c6ca642a418656ca9430450918516110a5c63392c9e0a244d4abfa73580a65e37d0fdf81ffa90ed14c150b49041d94b9451ea02184248c7df3b5d0d6abd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha446910dbc4ce32a2703364d421fd3e8edce743d1db657f8442d5a44ea987643c988f53bcb6a3bc2918f921064dd01e140a92cc94946b7e00d47587b59368e18809877dd96e66186167525b07b6381fa5f04003b958f1610b64014224c6bd07b20fcad5ec0076ea8a526c5c70fdae1c8e8f1b9e3892adf489e015453e520b6511f9354bb7e949ac70ae55829af1c632229b65438330c03bfb2301d7f305f50d08d00463c6c9e2c23a8a762b4643a5625fdc2e1e118e4ccbc646c8f8514cee54deb972239557e6dac618ebd2afa47effd43f5dd8c3a95f4897a2282249086af8393fcd2db7ca0cc43a25e27fa1222d10c38555c251f38ed225fbb050f0d585be6af130a339949f0c59c5e14d1f482324a758d0654b7a3fc53381511dd6182d5f8fd1f87801d89183a78566ac7a5e61e714ee92ea4a0fa95231c8f8a4889092681096c8cde681eae292ce770dbfb4bec422b89d59d14f83e3f732bc07b5d60b9986f0098233cf508fe9b0058769fe79a00dc0e39ff30dd7c4f4ce199060f1dbb7df5c222fbb18d7298325b98943cc4bf7cbb9bcb09db0279cdc25179a2d71ec8dff914617433280a11b1ff891fd081a2ae4fc0ad297899dea63c882f392ff6fc9cb616b0e9cf425c7647a8a4128cb019460b2f862c33bf31b190d251d9e83941373a0305355e4ace30c0cb58c85d6f5f021eed9a8b5a73e32a6a565c3e9ca665485ee23a30d12d28fd0be53773390dcd8d463f93358940fabb0637225ae2fb8f53aef5307d71ff154ca2283516268fbd8802b77bc45157acfd3ac17fff240266fe7fe9d8d012abdc6855e918b6075a86b8149aff9f0b523edd301eed713d5f7eec14d95a11985df5d742ba3219a4edf1ef3cf126c998ba0ac8d22579b066cdecc0062623b3657c27d0006a34eb092dfcec351c74e533d5758e3ed7ce6d946c86303af669b10220796ea0823e672139899f199e157594c1a6a1f31148152f08ab0c5f2d04074197086fac6a64ce85863f56eddf426d473feff037809b69cc8ecfaae805b9c5eed1953307a1eaf3f1da64f02e65aee228c57e1884cab9f2836a2e8e41b7716e5ca6b768a045476e9e9093624258eb8365a819b53bcb52a14d20cacb48f000525fc066d3312ea5c925cde4e7ffc981fd104ac14b15f240afa4c0c0f2e1dcdcbd9bea5b38124306aa6bc2b0e6374ac10adc607a45e914d066460bf52ad74884d63ec5b7ea06b03eee3204b4ec3485270b6a2b19c8ad308a3038afc74cf89cfd21cd05803756b8855091a3319a7446a0dd7b4e57e276708096a005fcfb62b40ff871fc4d3bc1fd1cfc717dcf7dd38ed5ac165ad71e859bd6172683de9da26881bdce702938ab8c02433dcdbcb7a82fbf178b3c39db2e4a77e86a67b87ad1bcc9a25394bf7b965d451529401b87f2dba83d14ed5a13416bf02d2f0554a9a92181c036284a7039fcd133f1f379129058623ef40bd2e2d2f5a577139a5e956b1cf19942bcae441eb8f22aec8633a518df7b676cf26dc78ffcc560f80fa23a0cf74ca4b303aa802ed8f51a4d9b263649dda8730019757c440d0731115ed8ab9aedaa9cba2f69e3212d3fd8690e067b91b8b4901d60815d153babfe12e5bc21e9680f11b615834c7b2a5931c22d2f52b377a283fda6f9f6c0af3cda85f3562264659aed69a2e9e9b1b4de6ce64df7690bdfaf90a2ee6e41720d334d6f81a311f503de28793a74afe7f5e447771e756d2d2c10fc1d78d20b7436bc9bfc9c56cc3ebdc8f44b746f87e7ddd973e4e5b0615a1cda7d4dd9d0c02d1d1d711ccea9690233cc27e011902c46c4de8c29ffe6367b59e6dcf9bfc053db479bfbbed658c10f70108626cc0ac67e2233ef1fc9ef56439de4eaf8b6c746fa667da9b0e09d8bf895eeb8450264eab19e64e96c0c7f7fd7555884f1ea0ef8219db5b3cc0ae32aad1c2c35d2fece7e076828fa4bd69ce355fc77df3bc1eef269f5c0e2939a8143d852024d0884e87908f0d48090fa8d500427eb4feff524f9b7b802c7a30d596e991e336ae69b513c049e73adda642871cae078d790b93b61eaf57192f898c27516f6cf22380d4c4ebc3de2a57319d886a97e0e67d2c060f7f33a4a4584d48747d28ce1a4b7a2975f8d8d8c4452c5eaae2fce5b00765eaeaf36c9270a755cfc803738a7fc59b20e0bf1187a84e6b9a58acf6ebbe0c4111a08994c0630b1a4e91c8e63c62981f5dae6dc1a4abeedb11ad6a937b99f9493eaa00b2b60baeca52ef7e6424e0aa7979c40d4e030795921492873764cbae5161ad0040a4bf302ed4e098cdb1c114ea52122ef95b8bbb59594a62011254eb35f4fd05f1a66f425f0c15f69b3821cb2f844ee10c16e476200df63f4063e5d7a377ed059dc300af9027630c274a5d2feff1f63d01cb5baec92e8bddfc361e7296215b2aeadcd105e49e7f8b50d7a7a6f63ffda9c5c586760d5e89ad7d2d6e8102d76bbc6b3b90c9e4d0a77d6d1957832ca0677f303e7859c39b98bbf257126558d02bda2132597ed72f26599bdd26156292dff193756f0339c3ff003aafefea6e1fe52e6e41c30310fdcec3c8a0f2ccbc9a2735c7f5e0e43cd4a5344c700b7955c2cca90253946621e18ae6dcc272ab9d228aced41c678d3010c128aa93458fa57def5207759335b3b9b9915c038d08d61e6a5fcf6989147e7cf72a0f907279ea1e87c91411213df65f8881e38e02f96f4af2e1b9143fbfad72acc093cb39b84071228;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc526a18d8fd99e1406b407b9d5184ffdbdb0b339863fcda31b30d7c9a82b2bf01fc99196f384e2de0deccf4010a27ddf046db2f8e3e22b533eaf82d814fd629c41427d54c5255425ea34d53ebd31dce66a1cb8b4e5526742f0b264eb6d9def80b7ad91f876bb59136f22a3294f427c0383b6686d883d4374bf137d8eb7a5fb256ee06de63bbbec85a8ca494ac9b60691b7340f181fb599ef485e27528f4993dc6f7a00e7426964ddaa22b6184bd85c7bca8046ed5d70f7a841d6b86a2b3b90acf94767944fc431f2eb3a08a3220bfc8d6ea00e1439cea58ce2d98a89707d3596f170820d59e0bcd1bf8bd5543574914470d8ef684494e300816aa9496f6f4eb4e12357bd2a003921411ed62b53d4bef2f7a7f864eb1b876fd8510eeaad8bf3478af33928ba5d93b4b999ab484abfe91b05d221050dcb8a943ee2e2503cf7c40d02e83f8d5ae5515d2f16fa3767a6778306766d56dc098d4d13511ba81208f6f2c8cf9a9692eb00c45b1d15677789054d37ca78f7022204b773082d93d9e8c9cb5978a0dca4c1d045e81110e2d4ef573443e8e39ef6b26b43ee33bd2297965f497e0c262c1fd25e28e66bcde049fb5bfc93bb0919bb9ba9790a65fdca219f3ee957e337b81c3576caa0dfa5e5dff7c3ad7a07d274db7323dee6dad6597fcd20820d081362eeebd1d6e089ac597187f80a6bd78d75946a9847595e97a44495215f39be011415268b0a7ce17a173ffa835a72002509a6dbd06319f3e1525c692834d42c1add9e217228b08531d3b87f1193882ccf9a61e54b75aa02b78850a349b3d8e9e3878354fc2115bedf79122a161ee67cb760002cdf6ccc5fbad3e57e84d4a7d7f485648a6a24f3052efa037a3fa93fd9959584dc96349a864c48da60143c89c30221574fed8a85311bafddcf7c2bd62f36bfd431f3d47a3cf870dcbdb3ef8c234a00e63454d48f468286a4f62d8918531f63b0933057d19a73bf289777367aab8bd8cb2c8a491d4d6a1decb5b5401b9f277c7cc9ff7b30fdd5a021153a2aa8900ad204d566b6f3dd5bc8dc2d99dc0977fec97ce5f80d1029994b45079d56861cf560265026c0509b37468b4056b1a950253316fa6c3e1428093badd4f6261e7d42eb41ca0fccf264c1c7f66b57bd2cdbf9115fe8a46d3aedf8c4c391bfc9cfe8a6955e2cf086f2be31b1ad44240d3088ceeb44d6aab10f78affb387463b8aada28e6e9908b9e5eef047930b28858d83049c3a8948e260be54eb9e833640ebe6e8d82d80a15f356c62e0023b91063e9c1d08848b87c929f40b7efe12806cbdf8fc098110b60afefd09d5b66d9cd045853454b7dd748d53656117b102c4b951b13131e1b3ccbea8ed7a9ac62a7da3af3f5028eeddcc14937049f51501cd6607b9d4e4593e863915ff575a4bc7d879988b0cf29426b011107cf101b57c205ce7637971477fd6d6f9e346a9061408e28f33863db601b53c16616aecf396d953f78b0f940e682e6f22732c65117b51d50f666db19d03e0e4a753b860be0396fcf88db2fa1f4556d0037f403bf13e5e0d4258e934bb6b9f54123e9529febf243abf8605140725e642fc31069f24e01529a70e7516a88e77eac377183d9c6cf2596ea60f79b773a33b9643c654f993207d4f6839af77678399e43cb78786a51ad86f92ffb52c3c779c04f76662db1bf3c0331f4c83c94feca20d8b6f610a22f59644fc991e64969e6d6583a5f33f95548b4b9c0c13dd20999db8b872797d1dcb42e87c6baf597b252ad28c906076d3e11a53031ffbd8aef51e6719f6c17886a37eebcd04d075319bf8a5583bc508402be03307c0625bc89ac6e2a1a480b282a0ba28b377ad161336f6d77b42d67580372c43b20fc7ac15c6b365e36a3b4872af8375b1245fa9cc3ee6d1e29fa9371482bfc01d694291b426846144c210349c949032127f93dd3705f7f3639651c533a8084b897161cc8861f497b67912680a5d2b70ccc529a17dac01f6e68af04d678476d6dbd956f58aca613dab4dd4e393974124f007515c3ebaf1c2a8ed267355da474b81468bf6545d72870557b0ee0eca76858881210db898cf03e607ddeeb6833abdbfe176607c53cae92920b51550367d19d54def57ab94a128d1b3de3c69c9c8b11ed424b038f1cbecd9a0d5287013069712e382ee9c8e35d159e2846f8bc881e79020a0a68eeec7458af1076d4992dc659b6db36cc9c43b796d62af42e8275da1865d89a47eea8924a61d3bf92f5c8dbed108ed422bd79bfe85add3933f7bf74212b1daa19311b5be6d75bc13d58fbbe06d4c47340aa25e59e732b3a929e350342f210e48f1b9f499015d38f1b30330270b9d4d635a3ab7054b00889e10a4f65796182ee5ce064b700f23aa5b96371c489b327f5100f5c3d8af950557d77c1e3ec6e37d022c0b639a31fb38a16aef6c55ffd060aaa9dc1505785fc94cbfb4c26917f0b5fd0e606f523b0a6ee2f0f71e33d74a5bf4f4e38ce9d145fed5b632467e998d8c3ffd34f2e87f58624be5b35d504deb6877599a8614f718f26e8704bd45f4b6403980afaed25c90970977539af2a3528d6dfa9574c61a46abdb1be9e1d118e07a344962b4d10f2ab958dcc6d9622281e3c905f964374a006593cfebd357e0bee148a8067885d24a3764960120b9794cdc18b5a9a0783f0371117a069796294ced3dc14d2986fe045160a3a6fba1e358c61bc1d3fc700322c582fc46d7d1b489e6be0911810;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9c00172cb427eecb95235480991fe51cd54ffb58f67967b8b28a72352aa8371c4e99cf50dd7a18445fc48d9e19fbee2e9c1b215b7186bd8dda3f56305f4da7cce35a1cdcdd2b4b2ceefbe5dcadfa98806e54025344669da54f02e14d4f314e04895742f6f5c7ac21dc05f20779dc3a159b7b033cee57b041ba82639031e04a8b42f18f4fa1a700bd9710f3b213e43c186bd61cd8582ac35240ee749ca3c71c55822e543106fdc071bab41821f826f1977c0a0eeb5fb7cda22ff740d17b36d6574266c71fd00683a385dc01244a3e59e64fc1eb67718b69766afe7c80dfc558126a64542f5a19b39546e6d05c67af6e1c17f4a30bde4fa10aef1c5eebbeca874cc3cf244769398b6c1d54469ab9fecba006af880c5554272e094183d4cd090f1bbda9d565cc0e678cea957ad451b7622cbbb07db5db01c9f0c6dce4c5f140a8909e44ff21dcd03600aee64fb7603c6d8a2a8e059af6d38474a6740d741d4477d82bb0b8aeb015d1563442b30a7357cc1a18b5b8b30db572593d111a2778160ba92e22345b2cd656fc551a1197a01bf19792eb76551fd90034fe2847d7ad8b452054c7a3d49ab2f73b64e81a28c80e88cb87853136da496d553b1ebcd0be0d50e879dd0e7367ff6fa501028e829b808427da288d2a86b0ef9f049d5c980d80e3c433e8868663a15d409cfb606b217ac2a2acf2eb8d8896d067333ff04b3526b879d623cf38c6d8f8594bdd9f3f0ead588f153045f1437f08a93af3ee435f866daf2930253d67f42a6306c2117017a8ed9c3bf2d53fe364e09a1a585825e23d17d7d4c2a3a354a3130e6c46810c6012bf469a200b8736730889bbdd2e00484b2ecaa558f2d96f8f607baecc0d75bbb73a0c2bf78ff8fb63f6f4ef08e76e13d441166c6f4e92d2099f8ef3c0802003e0b36df445793570027f19e77113428215d880f1bf2fc476bf1a47c70cd3a13fa09084314ba40fa9ca496461a9b0e294d221e8131145cfe2a919c7ec7da90e6430741e08c2f3e7475b159708ae737e3f6a9d41f49201ea61f9bf41f7a195db534bca68e57c864ce12ec686afa2ffc5c3b12c05bdf50a800713d46a1edf4140f4de08f44f7be586439ae6384433857bf76a9f74d8b5f8f5dc7f5a830d6713ac1aedeebd0d2afd78e3d2d95b004f0f3bb0ac0d6d498ef323d3792bf918de1e34fdb0c491723538bc78144ce1515371fa3c532f7baa6b459183976c6de2feff26928c78ef60cbd7c06193dfe564e9e61a5fefcf4add7f80bf22f8a5495a3b88c11fd4e56c82774dfb25fe7c74e0154634f5706aea646f2c4d7c31f73b2f4f78d62b6eaaf45ff01e43d81f0c58338b082ceec5643363e6ba69aed42ea47164cac1add6f44f0a00fffa2090129c12303ed54c19c69017c7c05371f5a00193fa9d253acc7e7654f9a5abeec783eca967331756557cd9577dc3556229bb930044a65c2e75db07f3e1ec647a1ed1cb0cf3d6cad4060975d1da07b125269fbd6e5077e4d221fc0b7b5689cff2df21b92bc32831dab6537009481688011c5123205eee042187aafd3cb95266dfee99f02ecbb64ebfaf6c733750001e2254196b28f03062460925e4ee7f65ceb96f5f4c92993a60fe250e894fd2d5666c77430ee3fc23b9672a83152e9c666b9522377de3b675cae10f39fbec4a6af2a8c5b9e38899f7b20971cd6e446bf2b131346687bbe4e7d404c561b8d684af3c20ff8b717718b8e7947b38bc2dacabda97e822ba2379a449e57fabc6c7d0e647c37f9cbf476e35df8f412cd7ed5261fc0600b351ea197baa00b083bb60d6ac17908ce03ebd5014ab628f7263e3c4f97aec52fe7eea07b8560574c16d8391d31ca9beff0c7d7fe5bad59fa807b37cc10a95691cfb33477006947e1cb4771c42e38a953f67a046b0859a9d8d9d6c6c35adf585fba97b05d7b4c20b6f21d88b8418aba16a5e775f93bcf9fb828ee45c14c2979a31530f39d6217d4d444960d07999f325a3675d0628f5cec4d2a237d36549e0d184d560165d332b9f12bde6403315f81d545c3778ffd83f8f50d275e7f6e8a9b0cc512fdec61dd85483a6f1e36e23f2f62a58b2ae117867b956d375c94e10455eeb44869b37134148f85da22850ef10b958269ca863912d9a16ef870ccc84e5e6f42dfdf7caf8e615103d25ebb368ac2f28a1d4b06a6a8f01bb938fa8255e3c49b5143dcc6333a978846655d9f03f726b7861851c2e617b53f6454794c874eb5e6319adcc618c2767e4af01e658d1802c18c79828e545fba2229869d9d1e805e9996e3f83ab04c225ae06ded8821cb08e8200da188b4d19d5528f0a722275c630bda7051ce2169da628d46a08e0a1dbcda76b5b9b381c868cba912c5b6914b21c5a3ab1afab9c225f67cd66c549743ef36417bf7fcad6b2127b80e2ce4448837a20e0bd30ed32d07ddaa257e001abbac329be80eded61f610199a9dd80a629302e8c56533ca632d9dd74a177b87c14252a0a6930d6b9e0d4c0c0241e31ada961ea3f22f8f7c4a1c04e3781eb3ae80f454d9c8a31e16038cf044bddb5a21402707e1c8c3b6d4cd9cc1a79e82db12ee350d76331903b5254a5bb006c7fe2335a005066f77bc4c865d43eac92313094b7ff4a4eba88267ed2686bd4812f6c80e4c41736fce936b6303ec7520541c4e91d1aa9616431df8100c84c930507c721d5f4aff3af33434ec4d90c8bc46399ebd3981fa50a79de87c51213d9f305a7da4e1f263d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h322c84d9f39cc30676b5bf43b74953170309f201bbeb73a65a06bc75a4c31555ac994dbdcc7cddafd260349f10706f88413b8843234a68f3464bc540954ba5e2d02b68591cb130f42f7ad5322286d33a9893aa206308883765164bf4dd0a907776950ac1bcf85693685d6bfa869b6d34b8830e5a05428b727e9977180fbe28f8ce54cfaa9aad49281b48ac343c209e795371eac7ae630be1f2bb63e3bed55b0f4d51c60419e5d05dee0328302ad81f31c4c81769285fe05ed642950d3af488137ff082d7b7cd3557e951e538a73f3e3cacfd708f9912f92c2a3c818016d60062ff004d3c476789d90c254b91ff3a3bf1c7ef40dca2f1145556f1271bfde8cd52f89e566a01ab680ae7ab699e77c6b99bd155c4e8404bb127384278484aa15f9ca131b48c19ad51920956d7182a4fee10d2d8edcb8587905a48fa747561fc358fc8b1ff20e891aa2ae89116f2e9b5f3ff1b9ef16f36583a7d77a25ac32952bea7830ae347de6ae625ae48221cf7dbabd141b301917b53f34575587264b5d5dd9d5d49081b205df68b3fbecce1b6590d8773e68e665e261457b082277b029757e9da841929b7bc53e032f63bbbbec58163072a8fbe45e9f30339b67a91268613619f4dccb5d5551176de4f259e5d10e9f5aea4e3dfbf4254ea676216479c8ad85adf2e3cc158c8ac7f3470722da4a0cc7fb1a622d879b95d32efe9b5029d5cd993a34587b097d4263a869edbd6002a9f776c2b7f1e1ce979ac778a1826f7faeb97ebd99c33961941d31e5774fd98ab167b083597c863e2c841f0a54e490bfeeaee779c55130b61e66abb142fc8b341ebf12a47b516eb4085683d7c041dbd13c3c119bbce17a1406a77b700569fc02b99eb3c533b690a73f599393c86b914ffab41a51172c9013b402f6ccf81a39ace50ce724c745724057cc6c533dafc6148a9fb7936f94c35962c4207237429ce5b523eff29516ca99788d28fc74af0b4276b7bf23af1e5503f9abb15663226d67fbf46d248fd31cea02e77030c8fd58295409c8b59577fc9e7add2883917a8325cf616bd09ec17669cb28ad339d4a10554152b39be364a0169239b7d1759597082e0bb078ee14066f5338f0599621fc1a0ac9fc1a791549d444b37a3f1f674957310bcca324780830091e484cba8c984ab4b4d5036270f497e73025ce7d18e8c1b5035e722d10e43f7e130986aff4553c49df61f620cfc64c1db668f3732b6cb151288edb33556b9e1a015f9a465675db781d9d4161bff90b741d039730ab37f03b10033d12ca1e92cc5ffb8fce2fb98cb4a65e73130c42a347c12812b84ad0e21fc644c17ac02ade5cd9de9d26853d429353094533b45a88191281d89cfb1fb86d44a488b31ae12db9bf8a3f1e3f68101410c3286307fbfccf4ace3e4f5ed1ed42809b9b2ed5ca06d2232dc97963b5271b4583b11e1c61f937b33cbb174ad2ca0411b5121bf16c1bca29c3c14c6534b983778346d2eb6c9fac7c069c9819c5377df5ef9dc1b23a851b53c732c646e8c649c6ba705d8edff2de72becb9ca542f31fc902c47362be13fe5ae6e076bcadfba63cbd3b5e2886e8e350ad1a2be4a5ccfbdb78a6f21e60d6f34b0c761b0a501858d7b50c3999f5ea569bda25253209c252f4d612f43327853362d5c6f16d80d97f23107611625b391ada54dc835d6bbb168f2e4d575e654252981bc150e74e43c2abf19098f77f2543e49d9971a83a91da90a758f7e754a9620a3b86aa356b0d897180ca10af43b9795553eca0caac1e515ff0a02ac1cf3e3291411d253b31a24d9d9a40d4cce6f2c80ba2a3c99c43c88ef813b4a5fbe47df6618f5791c3ea6f0a2a3a5de394cbfe5f4d91bea0d3fd60d3e599655d15d3f2a8cea7e96115252d01772a1bf8e027668a7e8629a23c678cca307353cb7e5134c177f060d751e6a24d81f2fdde0ab523b7f83b45d7f0e805abf26070878b7c7afd3c6c6291a64555d799e4dd0230464748a2a822e6877b700f9f039a7d1e8f6aa810d5d8a6b5d3fa7607ba29c393ca9e8247e1bbf8b952058e6f48930d6c082db2d8152669e6bec7c34795e7751bd35e7cbf51e26f741a6efffb143a39207737dbb20d5e10425ef3415a15070d164227e26ea342b0fbbcf9102cea980ebc0d98233930ebe259b6e2d489b63a3e62943a42d6fe91efcf73dc6f0a5a824505962c3ae274a89c5cd01d2915dbc14a70b67224aa986e5763638eed111558a5da73119eda453962497967cd842c411332b835fb746d825edb662d81948ae9e95a366db1efea8a454fe9932563bacf4ba2b197853649b37cd7d110d5f7acefb578f2f0c51e4fab770c170fdd9647edb4b5d448cb6ff5c726007b9334afb9011beef89596513b85fd6cee3779ac0e05ef86d7f080d656b2606c9943636191ef58274e8633478d84af8d7a9688a864b1c35d8bf53ad5945549b25fc41b8977cac81f721515f3e78cb1b9b2d6f6c3a78098f58c82b2498d7c5a0c0ccd54cd0c29e192724a5d33074e261fcfb2fe816869de35f15221c0c10acfd3cab4cc4a25e3ab49e125ad74126af07031e29851301aeb84a897413c318fa249ba23a88ad413a1f9c1b250017ee307e378f630633e939ebdec999cf84cad64c0812668befbf67ae2e159d267c9fcf737a7e0341d6a91b6aec4ab62628388392938d59b47360c77821634a29e11ae585c529f6bb6ed6611e7b1f172d1f988c1f03fa99be4f25c0a2ae9892bb43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h69be524a662222d213fc9d5ddf02f3a221430e824ddda3f8829d35f36151a0d45e072ce65191cf89ce22a21c1e3385d0b1af1af7471c26856ee0941d00676ff83c542406ce2b4032db319852c50e79c768e9de33b27c7091b5d0beaf753e8460b6e468f0b2160dd48643afd3614b9b2025f2b3a9110c9725ca41eab63531d3dc9aee94fb933163edf54eca6d7f1cd19b44bddc016bbe13eb248c61758722f301fba920a73f20f8df18755725f4d5024591326f07b48e2c21b7d523063c0fe4969f43988aff6cdfef7ca76601af32ceec12196c097a34b33775c0371e6ebdf916e5a9c135a3c044b779a530c81c1ed0f000e8282b6d5e61a8a3b106e095d4eee122df2df95939dbb58523396ebfec78b45336f4dcdbc790dffbec36bcff922f6e60f8dba1bfe97e60b203ead157e33569f2ea70be9d1ec1a3a25815efc8edc4c852997c1ff72c67e04937af16bd663dde7c75788cab64d2d5161ca2ff8839fe30c73b3e2548a53fdb73f241a3443b538427eb47ba46fe2a23a2ce4fded5044441ca82aadca53792c5cceefb054fe25781c665fae869b5264ef9df4268751c8c1fc001b2f96e11e5fd159a3e798c39e2c5122bada21a3d0dc403bdedcaade9e6844a2f70025eae1ec5be4f166508e44a8deba8e4120c632a17820dde5f8d6bc6efaa63f423bb9b26badd273e4e9c20c3497fb7d6f30b6d39132c52ee120da398860ba2eff1134722fcd19d75b2d388e53afd2a56243b36818bf32afd04e0a15390b445750ba989f95faea52d12377aa55a1de68fd9a109df63463c7f011415211e3d84a0b258d525df8b00592f13d4a4f6905a1e9c35fb863d2df9afc99d718652561fcde34fda133b92be72b9eb97463c84716be457e1e06e8713fabb8ca8a7d2bad59fd00386a402fabc241d4dea96d814817797c84023dd5e9f854856888b9988068dd2f02748670c39bed12940e1a2cbac5ab56f154f9dd4601452bccfe0740e2de7617dff9c075e94b636613ca090cc3daaf407522fabc830b4719656d23e5c69f4b70aa8b15f940f8e4ab75c34f0d3d3544df8c2086112c1eb02c34b97708879128a1d80489ebba9998ce5c0c7712e3ff743689332117d72cf68fc7313c3498e9f001f5808d6a483ca0b77706e81b67d9612bb81f06c168d6402fcc08fd2e203d5f0b098f4cdc925ab4fc0ce6739b0a092669d5807c5f5998dae2a46adda080e04174931f6d41909ea2573be6a00acfb4c583b8de757e780e949ef667b19edba2764f017a03f276ea647e858f3d99c3494bf6d2a5f1e60d9586551e3f72c00d105c09e10d8c0af3e62a373f60c603b5eca004e974936d7252156519bac23c8056e2e6f7611ed372ba1028724ee58258ddee706ba34af1bb97714848e1d7a4b42cf99384bc641d3c2cae187887eb84eab4978e378e6f2330c361eb1efd4e42748230035534857a4433e791756a58a7ebf45d7a1673f7419bef199482169b85baf974b9290624d6b5542cd7a718e290180ec5085b61d1e0b5ce48d03213ae5cfb4157006615c2fc263dddffedff645e1ed661f3d3fc1e0b70280f5e3cdcc91c403a91869e9e719820fde410e7446fb2c4817f6606210e525270d7573a857508f0c6bbc0185cac6678fc0a427a93b2403c25d48e69cf37149264bfa15070eeb83620358130eaee358440e93c34c91eefa065c61ee8a10305f3faf19b256b5836eb9f06880ee608815ba68a4600fa44e650d597659d33ed83c53f2426363a33957acb5a8a2ef81f1b5bc0849212bc16d68e370bee96e32b9a607e44f092dc60b397175fe84cfb5d669375a45a2aa306b56349e309f7aa88daf4c7e2cade6514c3aacc8b6c93936b14152eb7c1f7b2ff68d5ad4dc4e2790c4f35a2ed0c9239c28f3529c23843d50d715ae5e05dd17c83c8f731831dd1ba012ba4cf6021c6a43fb75a9426bdac7909acc9dcb7e0ec85f4647e666b4172255fe0a8df26bab47334425743467df30924e2412c8dfd585add7e7ce73d6b9db5db71d22ec85772488152061e96247783cd7b2558a251ee538fb9cbb8f6a40b9d6c5db11ee12ab52799554585c05f84da5fb9e2b629cd91b1231e2735dc24ac22dbf0481172de0a4abcb13c485de401024bfd8f9f2138ec96461d4eea2369509f87fa44c5de1f1bf6ebde5b34192cdbb7cf0d53cc7c4b0bef4ba71a2a6ed327d0953e3d049aa4b57d32a8136ff1552172776c2b99cd2d5363377f47f15edfaf4e9f706c7eeedf9a6a905bfc7101fd5a9aab23fb0f8808f346897467ad485afd398664ebcf728df1f7b51712547894bd60b9545a9dc3fda278acde0c28e113f3d0cb3e29f698cbf7f5854c9b24910874ec23f8d38b517cdaf8b7d8ae659db288db172c7e3d84c66481fb8ee48afb7cb0209c86a68020a3c0a9d95c3b2338bdec60e55ae4f1d75c387db9417e5076ac4afed1fbc9c1e04344fa3626f5a178c5ca4a7a76fae36d4e48ae20afc891abc9cd6054befe94191e1392ac3b9bdad392c7fb93d957538c2148ec0ef1b87585814d5eeb1674e0b375b2029cd8c9341dc08c5c7ee922405d10f9f8a19d7b6456fc26ed88a6bada76310bb3db0ec3d4bf910a9c426d85d3bea0e3fac065b905224c39a315a2836022c609f29601cc9ef99e260f337947667d24b2617c4763caea02a51d20235eff4b2dccede77a517f747b187d78c4301c0509009ed8d6727526a2785381323d7b2dd32a4534938cdc52dd06c6376;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9619fd36ea5d1349ec372909af48ae18829bb736075ff90d431c9386f67fa59ff98331e20787dcd3107fa01bd18acb38ffbf4f935ef25622f949f23ba006beda8651770317925e04d9df386770d6a44f5c9392c3ba8b23b4f0cde2ad34186fd07ef94f5c1f232782c642ec7f8b4a136cc30510bccff0d5b2a36ea08ba7fbc1e164c2f4439e3dd66915d062fb22ed368b037dae7b2ed0d0ceb633a880b2e6a82d295e419e084c3845a3363f53b394ef0f33f1a74bcf81fcb3234e989f892c714d4445f6f91afd5a32537a77df12cec172e1969f2da84b2f1e54874d39047328dac4bfb10821ab6ae8b87776c16b81bc4df2935d9abbbfa9c8409fb4fa124b449566baf3cd19a407b1670202dd2b6fe83c6782644e112c41ac8b47485c5a5783664195a604fe0e4138729d144e49a02f1cbcae9860aac5ed167b9e38b2b607e101ea8cccfe7a7a6006672ff6646e17b54aafc37d6c9fdb2e5f62dae717a4a39a1a8be041ed4709a9e314d481d7f46d3841211ff06bcf2a44d17084c8c996bd5aa76f47e2902ea41adde55b72e99b56d9c3634654089d2fbc2563ccc055e04101cb2d23479c0a084acc449a0c118a95a8468d5246d5340638648655436de708d04b1bfd66ea7a57fea2b02379fe4d8503d6c35fc16bf98577ae195b11ac94b900b01f10b6c3cb69fbb1b5977d69b153077c59dacecdb0bd99c8a8778079c8b87de27124297d5d4a2bcc509a26ea79dc840e7b9eb75e3ba3176ccc9891df4eb446f70045df94d9461b7e15de8210d6c41bad4baeff74f920340217c94cef092aef3e8256c95614cd2434560fbe00999e3553856220f7c0a832b78506ba170b1619b97eab7160c856cd14fe27ccecd7319fb9afcfffd43bd37cf7be3bd21f6e935584df4c98693a3e6726764152aae5267f1574dcb2e5ca65b3bf0013cd4f08d6c15315ac4a912becff1d28ccf040d7785687a7ced1dd3113f210a43261abd1748a4af2279d4b47cfa647ffbab4fde4b75434d59a7b864350c0cfbb63e0e8e2e5f8be9199b4e01530568752ef516e9cabf6eef100d54804c4a1894ea6b4168f8eebd7d470920b3079fef729652386c3e0c0da2c55d941ac8b70cb742cc7e5b6f336b26df88d29ac38eb1ecc14dbfa9c0a24f69785a2ab00527d3b803af454476f3b65edfaa3d81e780322c3d09d4fdcd820ae5cca70b0ae77c8e5a5f1ba9450105104cd035a98cedc3629f7e0111a4d417511a54fcd06a525e0d70e2fbe0c5a5dc0e8e84f06293cf67b0acb46ef03c6fd5e01e4855ccd53fdaebb87a77a33bc7785d8adf2427b33519f316515ebd8b2d89e48fa7699b31bee3aca09c2f9da60806941264469d8c5b0d1b96c1f8334b3fd38c9c4dda82859962badd99a79fde20e36d4ec0ddde563336b925d4ff324bfd5b226e89c08b26bdab62f90bbdb12a97fb91e2cfcd4b4615b65cb8b82d4b7eea22f17dcb44bf0aafeedebe05c151d358ba46371bc7fd8b9f28111cc6e8a03ac4cd48171ccc4d03a9bf4417b53bdb821b5177690a1e8bb3086f043330eef74afca653621126f312918941ce204fd71086d32116a56478fc6b1ac509ad1928dbe2c0aabf9f33bbf78ae7f9ec2bbef143cf855d2b25b4ad2bdade0447719e6d89b72335bb07c1bfd7b82da1f9ee9e908cd0fa2c140d055b03099bd5f0248ae72863bb77620615187ba127959435841aace88bb6af3b6e7fd568be378a07cd92dd7b8a9dab534970a3b7ad0ef51f5f60ed2daad7914c8e7e6a7ef37d1b336ae38051eb0151ebf1c50aff6121d336c34c93002207dcfadf45b27c3c7ab27547cef073f784305a2947d47f309ab4f37f9c4dd2a8cc2183c6ff20fae75b967f610ca14298d150e1e3be232557013d87168f3c6cff6049f1c4b505230dc936b3b58f7dd7a705b1a298545784ebe0d7f6bd61abd1cae45b5f145e8d62df75ab355e5de9a1d638fb4e390fc2ff3d93efda4da797c984d5e82973259257f2af437011c6605fb57bcdf13f62b83dc714a53e2b9f34a3bed223947d8ce7c78bc65c86b770238e6ac4b2314e893c58009e0030474981fa676979100ed40bb8fdabf11e5ea69fbb0471929c03d0b4e108c31335f8c55a253704e01154ac400401b6735a551420e0bc04b32eb63e724188130beb5681580392714d22059c6c7c6b7c68dce67805d4d8f9e26165f0e222b25de38ba020e8b94660e49122fa70ee9b74b7200a439f2ed36a70f342751e76a080737551b85ff337b53ef9f5b8c317634293ab3b5f5b53fe2294f932b41eedab8ab9b563931d68066bcdf691dd808b1585ab948f91138307d4f00c084cd894d9fe2716b157a7da3e4d7e6c99234d2a04392d089965791cb89b0a3580c6a628286b494136b76eaf4b7eca6e6d89f2f755865cebeb367370c5ed05f3cb36c708b69731ca94c7f6e3e09bda70b614e8940b0a797082e58d61687cea5e1845a3674d559b6b85b1814444c61683a52bdf1e975dc33d8aaa77adaf975869b95eb195cc3d0d45a0fb29665100d6a07a8d299078e6084f3379b9ff348210bee1e37b1b36de9a4b4ae537e9aa335abd24c2cdcde0d2c781a8b468dd6e6890ff1e9d099d08cc19c8c5743601f20a9a88731958d9a9781ab88d20a99e9f3b20f3218e3355cca62205a8fbebe671c1494371d6c8020cf2582e57e9d2c73b6bf0487045e971811b390ce69786a4c4ab5cf30a7ae9270fe4d5035762c47b6ea0e8b9086815ed84ea5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h51f6922a7779df7b4a1f8c206ca4c9168df9189f1308da2aaf2594f77cdb73f431ed65ce2b6c2e6fd96ed92232fb5260dee16fcee8160425611b74d69e1e9ef4500212cb08e97bf2bc857e580c32e8e3607aeb188e8ba126cc9b445da7eda906d11e0b57e4c9fb427d2587b96aabc5c1a088a5361dd6a85108d565c0ffc1ab61985a734b139e3d236e453e189eb63a240f38541c2ca2fe67a61e28bdb0a9a90518d88064b704d4c29f74ff68c22de5f8acb0a788af8582d1a36de7af799608ae16cb33cb5043b1d51567eec2ccabbd01246a35fbb04db4a2b31148d0cbcc690df1f51bc855d34eb5268f77853c1519c21f11f8b8c578d584db3b41abc98cd319d92f38bf503cc7e533a95a5b28ac14fd379ca56b842688f5414b34775b169f12ae33a32e08c5f8b7ba4486f143c0ab30c525d95af795137783694667b286b9053c216a8a7f3da1475d80461f6adb1bcc67c3e491da2b282def3188dac9cbeb4f50dc4dc2a3d255277e3953aea0c661c49b6911080d03a9309aac94650a8278ff6980c593a4477a9f62d4bd792665564bf9dea6192a8870c7c39cf6afa65e92d77c891051021ab79a35749de5750c6cac292b46f72d5e7688625a77a3872f9367402c55207ec12ff4a2366bddc9b9c4c40d94457a75505b554580063602580acebe1143cb7c9439859e0f99006061eac0a223bbfbd286437d8c4a6560d60f6a944ca5f78d1a4323af5dfbd50d76491b07963e582717185707adebcf0e14d3b00b8fd79d0d10df07c4b5ad18fcd66d6cd85e3cab67823ab22a10bd61c50eb015c4dc8d944d44955abb4a3b12e25b9381f9051463941cd287fd55d2ba110fe5a17fea285a67a8376bac1691b0bd2e1023a2d6ec15a3aebbcf3be90b009d4239ac35bf15eb1b64e3bd10737321f5b11bb6db77e56e6a7bdea6cf3d6d863ed9c143d5387c9d35bbd4d13144e3286529fc17cb93548a09e6f2700e67ca63b0b2e34c07b3f11225d8fd07eb270714c16564f664e085e6b9c11149d8e6d0532cb6dd2db3c04eddd3849eec676ea8ee036c1993a8244a175103e8fdcb6e8255edd7fc11fb5335030acf547212ac834cb81760e57b1f939847cb8844348ab4955cc760651486674b956835c13edb1368d26d2680a402058573d3edc52903129a3feaea1e54fbb3d7c23a1c59ed8222a962ae45da38706c65b271b5e87ad3019a49570789d8ab66bdec66b035a652b2f67f8156337da8c8cc11887c990b6b444ead292ee30d3a467ed3d1b8bab1405e816927cf21261a966e1eb9098a969cc9e7033f66d27e994d38577a51b52d356e9f6a001c4d939e5bf2613634a2bc1fb91daa412ed46319673c77b1e08d8a8e8d1f27edbdba41b8ff9d7ec8a836e822950b3034743dc89da23c2d868f3919f9a1c4cc6f71cad82ef36011665b6a7b82adc9ee842f5a3fb51ade383436fc9d2ec4725a3dea015af52907fdc0da810f100e5c66d72c178e5b03dcec496bebba3af32411ee84c8dbfd767084c557c8a98ff02443cfd7a0214f49f62f3b6a2ab60d8dd46b30c106c335a3d188bf3ae6b654e8d7bada47ebbdfa3bda63ac87512ae023dfa5e5b82890a06847a6d55a8a5f2b02b9df3a91d8bbc318f4e12a66290b60363570b5a65d76521ca3656e6bf1dde68b8ec7543e2ea6d6531e761eaa5d224dc1f7312582315884c4f4e9b7e29f85ce98e7aad1a88f387a8548c6fc81e8692a9efd83f80e9b6df826e7cedb959c22cc73b106b0c1163b6ff684152e7af2c2688015e23d3dc427766c779319c38570c6487771359d240a30de6a65b0994785503aaa73a82575f02f791dabdc4b6ed03e5c34ba049b5616017e9d2b8128261e5c8139d9abab25fda6d7fb83c78d4182032823f702ad3010322f1fb090f6fd4cbeffaff889fc78eeba8df2c80f748f76fe155306a6ff73aa843b25230ff5737caf57986d1d354407f28ee18d35b4284c44dde47073d171e054d3810b472e01bc6770f20b9b06be7e4a9ecc27c062eae760bed0babc82361977117effd97c8fd4e1576627fe4eb6abe6f989b547ff187320b4924504af2670a64f35d3b22c82d0ec5960b20870cb7f9dd2df145c67e1296d85d6ecaf9a4e5f0f38fe9d9049082a35256ef00f0b1444c78afe14a9f5f222ffdf899b2da24801deafac814ba636a62ff1ca4fef5cbccba704fc5c8dd2a46491059ce997a2bf744f62d54e8b4b0b40609f19e68b8e4d08edcade12c736e9c07d9894814fbdd1d0c07eefbc4a5ca52c374570496d9061d75cc8a173a71168fec407d215a8a2f1c64cc7db1461206a592a4321ea7e0ba8d3e706f225a9c17c8dc22565e17cb1fbec0751904710b39f2505fb18be4683ba901b5f68b9d130efc6dd03362c9e079d50f65e01cbbef72efb2d4524cfbf01a30e57428f2c039506e6a11af169705809c34db8627abdbaf43cd704112e80fb8d13981e84458075f8fbd15b277b77111ec63c8c22d512e79cb8345fa4328e07d583227828c8c7dce73e9f43af192890553047381a0d04d8b64626b0763c48a759ad98f8859cff609d6350c7a41418610b08c4fba9aa33d017e0826098001a60e955752b59ddb7a24cd1e064c17e3de7bdf31ca47fcb05c6fbf4b676a411a34062b7f00038c00515bb14852011c27b9aba00e354a0c5e77c20dfd124c391be7686b6f0994a475e2506dd8cdc2f15fb007ee8a8564f1b61ed2a678f9562641ee667bf8dd1c195775de169;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbd6a51337f2ed7f364c02c580dce1e05da079336ebdb68250920b863b93acd92eb9f47338965ec197db0a7a4a9d6ff3a5720782c5b85ed214b118242a16a4757915da040a264ee4d259b6ff6e64e6275c8471ad9f559b90db6da6264f27ddc0a3109e47a94737fb74f037f310688c99a54c3561bb0270a6a129f55acbd86119d39df517946bcbb9a6e6297aa430d461b14b31cdf57f1449902fd41e6bb48bad6f9928280ce5b3835ff9efccaefbcf34ef324ea59b17cb733a734c9c981a933cb15c2d4f886c31459f4824bd39cdfe952876b08a445d776f4c1b6a07fbfe821558e2f36b77d34367465eac11069279143a8db70675a3639551667fa5a688f13688640a8b9652285fb8d934d0cb798ddee9f3710873b5d7dd454a7174e096eeceda53187ce3b7f3e0cd5e4743197aa3e1b9d08106c1c04c45f5696b6fb8556d09c214a17767cc953db9ff2fdd7d26967d17858db4a37c234a5b83ff0ad1352f870424899e8f3b4dd5be864c1b2a87ca644c88ab8d6700bdae8588f44f7220712a0a7e5c0429325755786dcdcfbae879efea3751a48a7082724cfcc117169b48a07742df3a20a0eae81463d1fc1ad324ca6d7f7be3d9b0a0fbe95bfcaf436aa210c4938ebd9e76059cb335fea10bcaeb580dcc2c2477ee2961fdb3421fb8e754579f1b889d49aec1ad75507b7aba1832c9a4c51524c41aff34c5976ee1aa566387bf119e89a93072edb05e21fafe4ef187e273ad31bf944fb7d302a7ac62105e86f824c86168791a5751e16edce06ff27bb07aa42b11200f80260f1d395419776d3f82d9a3ff085b74c4afa501d374319bf5da719afbf8de6b4245308dccb5a9deb97668fa4ca54cfe0b3be110008535af3e64a990807597e70d0f6c59c2e93ce2d311641949dcaee7ae7f478ddca4a59c4df8ae31e2553f302fea683ec17562133b3d16c029676a25aaeead21f0ddd44861d74a103256cc9bae31c5fe24137f19639d4f9ce16cf46f9682e4e3eb686d070bb40581ab21750cc08c26022d0a8c1aec2bebf02a745dc4e37820a17c73dda0a57b9b73636d95992326bbe3ca798b0feb450c0efc6d5628b259e002ed3f12e49c764c919520e8edf9400a0f063044a14f5904ff1cfdd28a9bdb606e5d3c7d49a92ab44094345321cb6c6552b72af64bd8dce2d1e423559dc2c6f035f8e66f165424b62fa7ca3da7488cba06df322d4378ecb9b82ef7db7d4d11c71173a68510db873f3780aa8c5299a6cb41ab781ef06e71282e5ddbdd87c77f0010b33d2a0c0cfb129497bc42925d540f078f9a377049e3d6d92fd9035022efb0f7b7c064d9124367afd1a2bd7e1a676677feb7a1dc962062f1867f403025f9008213ef0e76e6c685d0e87c90d4e5acf1bd2918081810159374df46a945833ec8e77fa6c2cce792c437fa61baa9c99b9d195ec7df525c2bb4cd26d6a7e1e09726d5787b8af9eae07145a487b37435b58fffd02582751dad9efd6a33ed9ea8975fe27198a63df0d201a6a916474784577d527bfb6a65fb4ecc7b15896d4063e35c3fd09a69441f4e0452c63b271b0cc250eb237918fc4119f4ca8b3ce5f905555f36d43b8b44376e54ba46a413d1bc0a826f7e99d0a5952561f9983b29bfb49a7d5bb6dd9c8e8e340bb318b6c60048e94e975f07219860355167b0c162694c83a62ba914f440de100d57003154e1fce3c6abc9af987508d83c355761f0cf7219f044b0a6b34fd1218d714b18a329ac3c65e63c44b0d5ac64557cb198ddd8154a6abe8299d5e6a4c0880903344f28356ebb93d15d9900e708fa864fc5060af8853c5b1ef310026acd344cbb45b659113ace3890dacbc256a8bb39b236c3531502de6c1123812a7008da84e0e9c12aa5d0ffcbfaa3bd1cd07335f8d7a58dc1b2be4fb017705bbb71cf2d766eab835a36abc96050f7fb6321bca0920ab659d6de2a5622d88d6903e265cbd6988abe910b157ab301d9e20eef88f5ecfd8e199769f30c5ad5f1525e16e613220e2f599bbcb4bcbaaa441d5c7ea46e3c09f8a25ede814a16e51b3575fa5b4a335c9d2d539dcddcac0d40a48307eb1b1dfb9bcffa08f9ccec6a887175c9ffd918b3c3c67d6d04e34d860601983c36337ba72ac6ea73e44880adf9ab5f194ab91f6bc1d6ce113d68836f2c1c45b4eefe93aedb9443f734c42a339cf212c4cbc2d74a16ee204200027a33f9c67da08f317b078851183ef2d0a28b9586a53dc14be58754ddd67a4f0350ee42521cb3ae3a8fdd9d267d27c0ada13e5fc17a487232b00b3889fb1bf8dbb05f1ea2cb820da26b4c1c9262ee982175a47bcdc063264932edbf7eb91a2d2187e45d3bced18830e51f2901d0faae63575fc6497dba28bc4d4a36befcfb18535029c84d5af27659d79a0c234bc3ba0a11f3c6df3072d4702e564e036fca8fdb82001c3ff388f8c35d973f87c27a6a7b7ea3a4be7d7a99e7b7e270f0e2025a0f4061fb2c5cb0b23208ba6eca28419c3f4f9aedb3898953fc8c581307f9a5e3bde513280013abc619c950f9611cfce3d7fbda9188a94e9d5dccaed6c750febb39ea9d69f71ab7a50f9d1ce5e1b917ae8f1a64fb49059c072b1022c24ff93da8c4e1cdf9a06168bb0e91a3d650eed6b062411ce8810dad9bb6f01dc3c4c6fa49b45194aab81048854c2cb58d8b41cb1013faf82e16891170a0bf65079b28ad4cf1dda566958bcec04a0620547b8989ce02ce0cd5dfb22e5d7dc88565107ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7eec863766589581e01c7219b79396a3dd470ec47f3fe288e5595d3d4cd4f13f0bdf6858cf42e843fa1b72897980212d424fb537ba38013c553dd1808c47a780da4b57b0146ebf5da0e2fdd4b3345fd220f1ba7756fe9e41465ad9fc64223e02b919729d634996deee3b2fa245def9cc444fd52c6de7381262f2807c3208d4543dfa025ee43ab1e3d4c4f0c8a2bb35aec7ee038a62f6f21181c3bc6b7f59d251528316856b94f6399747c1a206fa602d5313f28f38a10f20eed96bd11343d589bf7270f37f48f39885080e1b8c101c9aaa7ed3d06e72fd77a09d04ba39f037c49cf45c3d328ceb3f5c3ebf8a11441ccb733bc0515a5e3a8b94e112e57c20ad5b1e72fe64a9f591cf08096f58836a88d224fb48d3c82d790abdbc42ebc24be2e8deb2183c3e5afa1f68805f90fa1c5baa50393548891637d3367a9f0bcd0343ff8151f6b3eac44ef07aae07816794617b026b1b00ebc17d40747de742e177da251f948d3acab79f0ef70a356aae539ecfdc954e72e9050c18d4d5f0b37ff9fa4c9ace562564178990a2a879f65605473e1d56d65d3bca64ffb3947884fcfa607a0089fca48fba48a4b39827276bc755c6730f816f7c2b03dcbcf54b064dbf6ab6434b474b5a00d2d6070fdb26561c7ff2ea18300d54c960127f6b0d1697aeb4718e19a566541a5060d320e687f690fbd48f09ea66277ec02ffdcb6c1a14566d9aeaf0e031a37b7cb08ec0fe9281fcb460343191ed0b156f9cfc982f8945779d1dbfc840aa540fcf3bc49fdb5d4f4d1a3a5d3b678f10c1287c6555e5e8fd1272993a47aba1619c107c9da3712018edb7141e254bf7b3439c41ce6fe74ddeda23fb07e6519934bc787e31117c9ca137f111b8e4c004f34fddae4e40c0451fa082008c8acbb3dbfd86c103baabf95e5a32c955e2c9937b572a5d60cbb69f8b378436a1bd0b5b7f6cdf8b11044b3e5076b63a27780a865a827138c630447187804f90ec9842b9d53dd8963dee4b3ffa501dc2eb21fc8ec16cf0db75e02b53273be1fba01377288bec9a8450346b5ef422e721569011c817548e5ad2ad59acccad3586b862d1b6eb4cd01be43669f2092454f57db0bb229e5e7fd94bde606b3c7303d8705392667acd3a2299c88277c2650c0337ddb6fcce8ee234fdd62a36201c48a286e4819d07ecdd312b218a9abbff6cc5edf5b80daf6d34d71195b0813aef335b5a822772ad230a1a4785059cb882b3f4d372d0e86e4bf88147deca6299580ba27eb68ab5db82c411f5fb33734a540c52339c46f8fefd304455fae9721dc9bec37d75bcdbe73bf0311f65ae417cecaa8e183361693501bd977bf89244b0673f5edd9989bfeaac0e8029c26176bed8f3a369fc768a34494a80eee6fd151a08c00454ae9dcf2d2e26f892fba13031bbf754cb16984d844688e4c124b8d9dc90712c7eb1d46c1f1af0643a52fdb178778ec67c5f50903c2aff61e5f60e8c65aeb8fc97cf6226b7db3e76b91647ef4aaaf2dbf0bcf49fc842047007b89f9c1ddbead8f628b2e69ef3971bed8924b0553991be6a209c84e62448eb730252b5aa21e3e24d9883d67771c1923285e8dc368a5c9f8924f483a16bf43b7b938664781c5bb14669b0e19c62fb74409f9e5ee88fffd1b55c4ecaab603346a8694ae7655ee02b57310ba205aea16b9f54996dfb51fa7ba5460c30203cd89d27a238bb8813773f0cf2a1046fe27d82cad2fefd9b9a201974975ae8eb34554fc9d720e0b7e981d2c8cd568242d476a14e69fc5801a7bf661c0739eb079d1af4ea15d4c410f92c3271d244c7e3da02adc724fc84c4d7c1ed6f0342af05eb164d17358f7356765424f3a013d980dabeeff592146bcd2e9041f327473cddecb7511966dccebbb940014f67611893976b67b77f5eb6bcb387f897d7e5825ce8ad9974374b121c0ebb5b2620f9a5d2e3814962ee62bc4144e0c67ea1ec2541c4403200f5483cd37be31eb2de02a98692bbd04984ed8428ae6416b7d2bd01050c2edc6284f320ed7c36e642af7da22c40304b6a72be854063ffcc553b53ee3924cb424b365830aa5c635c691882ed06b6fa4424f28df187ece4251bbb4f8481aa5c77e030d235e15afa665594a3b8f116f6bd62519946df4e233598926b3e809112dc20965d36dddb15b2101b049dc30cb27e0c65f0bc0d594910a65acf209d955c61ecbf6e9662c32b8a71bbbb0bb393c210a3122748014e2b7429e71e913adf1b974792113076afc6f35ef14358c7a28295b52fcd1f337107a7b3b15444bfa8f1c700087d5b05ee3f3d9cb88c071156e5fd6a6cb15ba332494a47baca8c501b048e73c823aeb00ec2505e8a39aeaa0b6cb4118fd9a0a7916e96271f503336f741eefdb79fccfcc576090796e52406defbd558849784a8483b00ee6faa453e3eaf767882ec010ec7115e5dc9a023ddda4ce0fbb528b79c60211cf94b54421c580b06656c22a47e8efb2ca3594b8eb28722b70a806cc4dcfb5ad3b5308a3924aa816e9e092a44b6ebe41bdcc7906842cd6b9ade2ff1d4d9ac6ed2ad092c3dec8300582cd60de294f7eb473bbd03f20bc35dc7f48523c0435b58a957bce5372481be68cb386485387f7a09d4b6709f27a840bc19ac8468f8778ebc8feb2fd7aa3393ceeb7f57484ea3457a39b144c46fcf8bfeb33a0efd2f4b7e36e8fcdc64e3438e666214d4992e168ae0238124b394d127fc985979409d71075a91223cbbbaac1dbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h85eb4a341ca38f3f6223d69370cb71d5f55870e38b620bb71eac96b9f72bd5cdce20d2c47a9e88fb90fdd609fa09f05315be9352debd767a72171459778ff5c9478ed0bb735360dccac84445997a2f5f52dc6d188727aa93aecfb0e16b0d232e74b215e649bdb335e040496926f5a1a12aaf165a4a622b9433bc0683623cfc29b33d0809a5653d4de71cd58f829edc92cc880f37300d4dee180f20b5a9ecb537bdde1eb50c3be42667ac1f36d7add9f300e8b4acf72d1c1639bccf2ca2a0312e2f9088c24e6e24b93fcd5cd86d75305261a355b8406a0ca56793214f178598276e9e564325e8979c1aeccde95a2373aec67f725d345a77a3c690974c49c3b1fa73725e4efa5437fce21d91658500a3132196888079c575c0cd8c2881063486a8aaaaf5e0fc2c51415148151a6cce08623496196f3ac540470f7bedab20101f5df9f6644d209087051e2e3ebd7d84f20fb9a7dd22107fd90e6f8b821e2f827bfb6deaf4630fd795a059dfc1384d42585728a8fe4c4630fd375f7d3f281af6df0dad4bb900159825b3bec3c85d9e6746e6cd6d8ecd6b892a9a7bc6e897e363f2d6beafac8454293ff39386bac8e22766dbbdf4caec0ea82cf892c1e53005f0d9781507e68e38b66472291580e3c7b479024a6891275e0c1537657f58ccb5b00eee51b5d52deb4fda3f19f97882e5bac45bad2a1e055e6277d4d203e19bb44b0d468f3c69859f3d836048f8c7e978d0d22444bf728b015021f2b6efcb43964c20d8f8354c225aee6b58b90bd0f169792af05d7e69bcc7bd1b89b2f0b7b34d9908e11f3bcca11edb6b5df42e1a029248b0bf6e03a02af899e1a5d7cac8b43ca201518bb3237577c89d70270bd7aeeb0707a6e23cd058ed5e074fbd2a3b92e9e56f3f823a18dee4ca31e5e7a5ee18170ed03efb20887ff844a6cae4532fcf012f8de25b20d7bee075b0819158663e9df080a1c469e5bfd8a11f8d9308ed479af3623429d8cc6f0b7b30b6dd28c83179e71bb25e0c7a30a02658b52a66a4349fd0f42bfa2e1db946e2cd8a0350ba6cce51535eca60d5e371f3b4889e963595054ce3549d500e6fca3e9d5c86840bb66f833c406e38508a2a297962e4483f4c0e8eb52adb932e5740a09209ead08b3e004c44c58527ed46dcd3e8f003db2693d699549cfb6e499ab8febe221e5b82f826a7bb2a6887e3c1ee368ac097ceda2f8a6a3b13546f556467daf105fb442a7ef7c2588bfa238544db780cdb2506a904cd78b10ce42b9ab187e25472b4935d8c9e86f61ac1732923cbd5a442daa4aea3dc89ceb6151327394c6f8026ba7a4dddc15cbe535da83035aa7ea509a4ea73e9624b1e545488eb3de305321e88f6d2cc011620d752b90efc47b20e3200d76fe191df08f70f97792dd75a591f1525af266025d4977b15a785c752d7e5428e91eaeec1a1aa383be7d0f65d971b4e437bee19704bc95ec17831a914ca46af8e129ea3afb18032960137ca36080f1faec158be34e61105332371c36f16948c622acc704a71d696ea079da6b6208994727aa6a4f8957ec290165a626d5323d373776e76ed1026e935ff38918977f4682996e6fefc8f53bde954190dbab7356d389ff6f2a36e72a3d07f0c3b1b358afcf8e1026b68120d5fba8fa92e8bda06bf40a42011a9b79b388a72e4bd11428250423029b59e7b8658ac76b6b942762f7489641668314d4a94ce2914538738d3d278a9c5aca92e34267716ad57a751af35f3b4893234decf859192dd84374d4bcb66054d70fc2f824500deba2de5b447312cd29771a9895bab18e57997290bb7716a256dbd1ef1a9c07e5e7b1024e70436e820f90899478544e4bf2e0e384b4f0076315c6bb2483182bfd1d53699c8f93a25039135712c856036364cc2e4d3b042c952d97f41a205667fe93d8e213c3f18a2a6a83ced693f0f454cea224f7fd0f476aa1983b4a04b94a540e2fd895778aea042bd6db81d614a39359faa32c11b3dd91c57b81137d8322039d8c46d87a9e537f4a9e26d9d99d8701060a6c019aa45b2fd8c8f12207dc93ea46d2df7b070f22731b3390e03c49488704f59ef1f3fb437493914ddd415a374f5c3f08ff1116d62a2b3dfa8a5ab54f39180b657719b06ee813be1e779a1c719f3d9bc13f7083f85c0195c67097e931cabe4db603b1ca3f0b8cab0d1b9a6dd3b28945a6dbba9297b4cafd895cd720883722eaff05322a5e5f7e53e40e302792a3798ca1dd9dd669994a2f5f0c5b083ba57c2e9ccb0e00bf8f285791ea7f4e53b43d0e896e8367aebb8f351d0ed9a5eeb9b9922281b9322be6573e8109b2e18583dffa06fb013f836362f85e279bb6096b7b008b3550bff5963dfd7f778c1d1fd7cc028a55878657eae7a5e090cafd88f7656c813e1e055a369443ad890a90c8f1452b4b26c2bad94a2c4fe7e265e6c9c387da16a60190625c3fc897ed2ec2c8de0518dde0a28cf5bd790f628d036ca1274cb39dfeab6b9ab11b6e5c91a5cc8c38b0c513a8fb0e64fb5c250dfa14efddfef8d0332a2eb6ccb7cf4c56aa5b9a899cbb28a75b229e03ba8565ce7c2bcc017ef8e97d83876a4bf3fb61c84616aacc4296f6f329012cf138201db8f8dfd1fc3578fe0c334266d89fbd8115809e67a06423853b210113dffca1816b3c6571c4cd4afba74d55159e5c6301b3fe84b3d7d3dc7fc79d500502f227adc564c69bda22454c5e6588f3d32b7dd90bd12e7e00727cd651ebbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc876e46390d30180829cb9ca07c07c115e1a23be2d3b250aaea321ae12d55f9a0bf72fbae5d1ffcae3a2537d51caf4ac547e36d14eeb9187fa49e9503fffca9bca57adaa17f6408b8772151febc5ab2a2060bb2c98d6a426e88fc0237f2360fbf4eb264a71c54538d3e2a1e80bff1051a9b41682ea3af7c7ca31484ebee5b061f519d474403493fa39f1c83d02ed9305b3db68cb1f972bcadb6608179684079e4d0f11f78ef30c2f1b5ce210122b90b54762eb9eec2a20849e6017e12b4a51af044317c2bb3002a7fb532b88da6b507bf18dc3cea673f7bd884774cc518bfd6e6fe8240dd8d030032d5bbb8190e387abd2bb41673e2478d3482d6ebf2f2885b9cf49a92d87ffc259ceb2d220fd501c3b24439634f8c75f1df47a89b8edb00d1d5559715d591ec6498027b1da198c65b8aebb25c4d92c11f3bd2c1fce138b27cdc1b5c0e6e43343f9dfbdf2ee95ab56d84b508ad19a41ed9374ec3963987f61b069f8ce11b3b7bd9a43bc5708d539f93da53d94ba78c80fce349876a1140e8215ee076e11d6d72697a805079331cb295b3ac05b77b9e41c41cf167ac8ebf7cbb08f03bcafc1be3de1c6008cc4139b3554fdb8da16ccc05ede71e30277c2253488c89ad1b875eaf622b2bd16d763ac0866d227b7c70efbebe2acfe9b6b84ef3bb07b80655901d6d9673931653603313b5596c97c35b26a52a6bc06c8b28c3ef4f16f8939e36b58e97859efdbcec6925b43671556994d6a94a65811d93f25e909d05bda75f45d6de83b32494af825952f74fa9fc4e472fecfad539722fd13843bb0d17717fc2423d53ec19349aa3fd3db5d60ea30802646c608b077b18e7dd5f87e6d5eb6fb56296aeb5afbeb07628438d7a0304b7790d2e1fb0ae4c3960ec73e2294b41e966077b6359f1fb873626a1d0f183667f6cd339c78beb30b25a595119cd7b6139333f104915f91471977d3b6028fc06caa1e4f68a31ef6ea2c4b682681e9aaa550bdf3e3e15d69904468d72c73c6b7140d26eb655193bcab027b4b4affff830003f7ffb9a02db46ddab710efbff5a32e2c43eb15f633985ad8bd63f19e77c289d988475abc0093e7de94f34c4b404ece5c64fdef73a51855c7570f932a6fda37522bfd64a361750e3df73e8a6fb68c14c6de904b0d789c683c5b26d32e04198b4078d46e3bec81e509ff4d7f958f2c8ecbc72ffbcfd215d793a0828eb2820a79341bc5e239deba619c2e29eb85025ee0faece589174f3464115f3cfcd2be0d5790b369fca36eb3cccc376728b667c33e2b05815a71ae6bdd7eea3884c153c7e2661982f6be16302936b24625442d7e2506f828f7ee6830eaf30e724f0f92a4d521c87f187e626c09053709f9f86d6a10289d86e198f3f2fd4c10e85d089c33c1f6114214ffe864ebc9c1e670c247e005b7e8872307dbbfe267012a88993fc1b93f5a9f4cda37b71191db822d507f8f2c10f612325626973e650212589c39ac1189abe86c78d74e46816273ec58aad45e7c39ef29ce0f71b8cdcfc4ba1aae74b61f76d12a38803c4de58e747e965fed6fb19129e8035a87370ffa9c32b8a5156de3a8f3b4b03d938378b4f14a0b2d1cfb4eadc87ffc31d9a658155e9ec6bb059ecdbba3fa676566a29e1760866bfb3adff95275f3d49a714a95275747d8e81cb4d5730d68d61ee50d48493f40fe85e6a4feff2fb6fa7e2b19c5e405ac6df9caeb408a85389a5a461f726f6a63db4e46b7e3ce3f8cab82ddbca799ab0df8f395837f5342c7c3543062b8a0b040d7b59b2cf42a5a9274ad1c7830794ebfe462490e527e7af190d7796a0dff6303d240cdd40129e620b8dbcbd5ab410deab7e9b63f209c2fb2d96cc4b94a02a5887625973ffdbc118d4e9a0c4b3ccc398cad39c763689a4d4febb0343621b25ac697d141276e54fd3594dd1515ecf54dad9ece04ab65234216c7c62eaed97fccaa446df1d273a5284eb3d8cb52ce9c0b5bf990a72a5cf62de233e3793f22eb29bce779a33a12eafaa7fe5dd5cf9e73e4e074d2c0d17e8a4825ee24e1a2b5b1871af2a6b458042c994438f923a0bb0ad05c0054ac61edc2d2b67171ad43164664709a730423623e0903ab124aad75634dc57b2f07a7f3fb7388e362d38069d31f6214f97b38ac5643b7515ac3a689d5c92c822fc8c630c7ec20022abd1763b76322858eaa3bec8dc79924b82847e13e592129f80d1b7d6c592e9601cc367927c5ae2713152d09fe8ff8f4c60aec1c25987f4cc0f4bb66fd23c19f03f51c7d6ada7ad189737ea33eb4d34f012b7418676df68dbceff3a003acbeb016a5b2a4739fefb9c11823e3546ebdec5c24954c4efe0d41c7f609e999ba0c3af64b2ff94357b3ccc83260ae3298d49f2ea8544273bc5aebaae9f8d56c7549b40a392a29baed5524afe3a3f5600a4df119e3fb76f04db073299aedbb41d96d6967e66a67681db8f869668da4cfbc057e171d264d951ea06995c9a076e15b1901e3d0891f3c70749b35386c9afb3afae55f59e11e1fc5563fb5b34f7e226533e33a0e5bffcd8834cb454fa0eab367495e004381a2cee7771a24df4cb7ed0ee10ef5f6c15eb3911011e7c28a64dcc45b23d49684f9d24c372b25f0ac31f6336a755eb185e4d0d37f59bee5cf38c274964efb81c39488f71856cdc3cc006279fa91e3e232b95070e35691bbdce6e5a114f9cce34a26518e8992ba1d9341a49ad91091d3503d38183200464b956966b7a22c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf5f0a48ea84eab2a20532392dbd4d83562271e889f12a55dd467901717e60dfb326c4c03344e5d9f0767081003896d26d242b963ed3d2ea9856bdde7ee0894826d85e4f3a439db0431a4511fbc3c95c3c7b28797ed99a499d6adfe96693f0cd06531ce7d67612f655c1a96b87305743a1cbf3f9a66fcc55a3d9e9d217a8f45d4e72fac180895348aee1f4324762fc9846892b6b6eda0f96f1c7c3797caccdb725a67885a90664a4aa9360697adca60e1efad68db682eb4e6b35c301722622810c05fbb83e78fe90a03d13e608957841fd232cec97893989cd506247e050c6f3da76f861792d1e66427460c04ad0aff057e2dc2b1236748994139ba962515ec15c307d94478535879af66b6002ef92e4a571dca946f83793424cd3aff7c7133af49d6547e3c743dedbd51b196e0d224bf3dbdcf451891ab2018b75f2de8c74850e1ef5c0d94978c1f6f13df67d474ffabffbf806bbe6a5f85fe8cacc456a3b1b6e8c9449f0cb7812d8a7b119a962c2396805790d7a91ce3bac7e9d1cc69cc7f673fd1cdcaf01dba30a3009921a455108f19ba5cfd63e5460b0e24aa6cfcb65d508b152f57105cce54c8e64189bd668237cc7c74b035f7aefa7dcd8306675180f3f7d1e84e69bb16728621f409b6c2f4059d3451e6e5815c99b5455027006ad2d182ab5c2308fb680dc2a3eca10748029c751992125f753297008604ef52776ed4ce39a53e4e8792a9ebbbc6c16720467d455c820b779314619c06e41ef2b15b00be138824a3e2357a9aaf049b504fdeb6618f9f1b871e0857a4d4e7fd22cd7726bf1d12bb58ede0434d8c3df5df317ed1360d434f56df5f8a6c110b8675a3c45a30e07dc46e6b13eb3c0cc3b50c2ac41e9b90a004bb0f592d86e99b004224bd3b4a82c485e984b309db198d478a7231c898efd731153f4866c9fa24b58819447611fc95bc282389196bebd6dc115236306d55aae6a9aa236d266c9da6559ef7c847c3edc8b6746bbd1522c323f5f77ed874f3221f3e8d91b14d13f41bbcd2b28c0ba8af98cba6861e10611a788037911974f41f170cd57ded3f36bfdaa1834b66157122990a642d92e246cbc50b2268521aa93165b65942bdd6a1de22d9ad2574eb2cfd28f100806a8b0adca49b860ca11bc659eae267794eb66fe70d563b1b982df9a21c0b9f95c202314bac33912a9e837f60e781b6da7ce8a46dc2a081311b9c31a709af454f8b2cf9244452fcb7f48dd2b862bbb9f711f19b569e9637e9e3822bb75fe704c08b7a433d239404903cffb0242966962cff2321591f638d10d4e4db97c66cb3afa7216a863ea75c74baf89232d299ce25abf814d1689482d0b419fe29d48f1453284971f527abaf51016c12f44dbef6f3ef88aa251101db58c94ce5fe09344a9494f5738bf46c2c7cd96c82fb422a09c3a736beb4bf9dedf13b6c753d6df632ea17171123c8a3676dc35f3d75995dbd5033e6194fefcd27baf7e8b5736eb58dbf1ef9ff6bc264c5219398a4d3aa24ce487d40c96f571dc897f11e58d40f5b72e2c3930abb232644bb6bef38d714057fd4b723f7971ed039bff0bf506e5f9c920d1dde20990ed3383358575c75242181f00d3e099031dc67f9b826b3cd6c7ab96d03489a549a27cdb1348b4564957815ab0f55a555a96fc3b1b5b50c09e46b7e9ecfcdaa0ab72ab55f94df732c75af9880618193d70d0c2ca3acca4c3e1f0c2da5a89cd9a02587cba8d5416be32f8cbd0cb8d835eac135016e423d378a6de102dd27f081501d1f367b817439f290f63baf088073e6509540f4a7ab63d851c4f3ee69849f1cc2858363e0c25d77a90419fc7a37d6a7d47da4771ae1a9b14de05731aa08ca1005c7d1b1a1d981475203cad107ef8549c92c55a8e9f4a9ff60ddf2960d4c6c48f352b63a2b33fa2fecbda60be0d17f5deecea9382be89214e2ef303fc8e8e0d09cc5f0b17bbfcbafaff55227bf81b83b861bb772f146a3ec4897bf771eb96c9a052a93a71be681ebca67362579b1e9d5f3434aee929e5edabfd7e9701c1817ea36b18bfa24df8ce8b18d15628370dd9bf1ae98de4d811a2c6965ad2d8946304cd8650d295c6cd9173a960bbbb7647777182ec088b2f37f2d6b81b539f9ec90b9c318882b8ab5eb77eb225785b2fc35a94fd4628f7d15123eb60b162bc2459596881315614aa27abb6d6aaae27dc3665e84bc6d436a5e2ad8956ca5e24d89217719f713a0d5f330d7e52b5d311a525addb84650f318c6cf7f9d523d2d42c1ac30186bb4a354867b51aa87ed38e658301d007d997b4f3e55d3c8a313782691bd8f2b3d8c91597d51519d5e52738743d2380df9120e6e60134288f52df5eae3efc44674a9f9bb693db15825199cca20ee60608550e1f2c066ac914da3c2e6527f6d70b95ac26ee0eba3c9eff9ccbe2965f1fb5d0933f3301dc1101d2d619c6f6c4c07b638bf227fbd1e469a63f7460d25e182f145d09f7420f6f1f11de164e737fcd7f7a45fbbf2000c2bb429f6df4db7cfaf0845ec1c06b8c08e37b125fd5eb6743ff639c0ea10a99e917283f3778ddb5591accf520acfe000fee11a2f1285b6e3bc2c287559c8d3448c9c4a17e58e32b0211b43c5ae6ebc3906c3cf9fd38169b1dfcaf4868daa997f827d3fadc6acf00b9eb4fc91920439eac291fe849ba385b0a0fb20035bfbd34d71bcbc7328e82ceabb26b76ff59728a0d37d39787f92863c6baa4fb33decb187e429f7cd15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb8fd2ec7f9953a10abc0fb8dbb066d8b148fbf7bc40e124724e70e810e678909b6ad7344645b2e9ec8df6ca870ba72956242b17281790ed93bcb22a1db27668bf6c60d2fa83af36874c8dec4a9bdf219f55a716d5b08abbb85b4049f5f6cff97dfc701d9f99c4e3a6926b390b3e05e9a48fbc3861cd65d24f9f00d37c05ea517042789367a70ea3baccd893f4f3ac024028cff757395d130babbd38623643cf08efa1c75a5eef7e955d6f7c2823e8552a3e628381d679a4d25300a3417615f1b1712e360f901314dd0e647ca7d55d795dfd041719ccb432a41731e7892ddec974f71e4a03b2fcbbd906a95cb3c4b4ac55fd9fcf908788bba1a691334d34e7aa4705a064c34e98a0c0d2ff8f7cbaeda39d03de01c70a21393d72c44e545a228cc1bc0d61f097823926c0fd0e6b3786e1cc70011a8d741c35d3ae8553304255b99ba521fbecf5edb320829743df4cefc230dc7ae3fae4a9d31523eab0385599a974c2c91243f8d4d979d8a9a809765b56112185cbf0a8c1cfe8482c2e1ffe749d22f23db40915b800a411ad8eb5bcc0903d58c421a5c30a4a7fde7cccb62bcbd2b99a5d69eed30bfe31fbf6366d76c56bdb70c61ba0a273cec88e15c5ad75d3128dcea70835941a7e7e9a36fc5c97bf5ccb50a28694bafd3384f0ba48dd56cb4b003698eab924e9b574aea6c412c12838dbdb4205b9f89925cfdbabb5cfcf17ab293b6519ffb4efd568a46c3de8063a08be394db1723f397ca22e8055d975c541e94193c59945adc3573aaf387caf640e3c99e205ff5c7d7c9e9cc7541056bc5d19fe072652e9f55177a4e1f5c6cced258301616c876e362feb30810e8140ace01ccc11306bff32c3df3bffe10a58dbbe9d4a75cde93b45786ad4cff7f8ed91413025e484cde93900ec6709e9b78a275ef369a0e10bfc6dcf56626d5880f3976529e1c30997a8049bf0742a8a937ab17ae580d311dc7ea88c9aa995bbf104bff0c250d3b17e4290b7e718549191c5acdbdc61c556e6ac44bd889c3918511d77ffc2f3c0c42917b56506acded2ef8ddf46823f7a652021d26f7f68d0c603f5a922d83292381e7256736b120cac49637a8e977e3cf4f05c98f2dcbae11fc531b817f3382e4743499b186588d0d39c6537e2fbf4b75d52b54f9e166ac24f20c1bc550880ee44136b15499c91202e68c69738c837d965dea0af2f63cf206f09a677ad1aaa72249d72a94c3b12b2e5ede03b44f3bf2f9928d141b906314fa9c0bcc5ac9f5e3f10a71093df34be4e21ee3f3569db109933fe91b7623c7b29eb40ee4265dfb376d41151080d1e1364857b2bb64b6368e085ef26e50cf692db53eb66f121fd70e4653e1246992a8970f375d9362047a06aad62c89830f5f1de93b1c1de5059af98cf9b0012d660628d39f14b8a41d1cebbe9a4337f1ddb4c3d6b112e3b84c67c38d356e72e63b524e2eab9b0e6394764a99b4dccb7aadad8d2df2a5fd97f9009ba8b039b0941a417a5ce067add43c035b201dba38428575eb857c1eda256ffad8bd620acb52ec95018816cf370a19cb1f7a7105d4e5b650eb41700975a804f11006792d8aadc4fac506929f7fc748fdd8580cba6b66a8733448d7e3e419d1c189b3da9973a6b7a35a5fa76c943a4e3a9c0a4de5ce71357c7827a586876bb600fb2fe7e6435d3cd1ef5a1d3c5e53c991997231209afb1aebf4f7827ebc46924f34bc08a2ca000e363bb743caec379a603f830eac13960e2fc8eb873ec1aaf5655ecb82a8551ce56b2e8bf433b4106805eaba6236d8b8044dcd615cac7cfacdd90b6632bd6731b38c7efcefa447c7a8fcca41eb8804b49e59f68b32703a508cbc6be95db6c6d0f57ee770bef8b091ceae838e399e6bcc6ea1598e45b1af67f6d9a272a451ffd009c74f94b312aef98ad8287fb7de829159e0966d9711bb69f46f8057e184655b97ec3d948d5ac0c2b00c8b93eb886bcee721e2b3b5c3779b408d4a60422729dbc5abbdc63e9ba687fa932ac678fc9becbe40ecf1304096c9d6a1da132edb102898276fe5da96b6c437b4068bed7f3232585b800143ba447e448df05b3014f5dd3ed320483c8ba7c238ec485cfec80d450f4fb869873253efa9b60097b027dd638d6cab3f39ad870c7ead96d832eec02258b62072a1a683273c41def91974218c0dd614330b01b95326841f15ec689529c5a56b51087989d84029de3839add0b1c8906e0814c69ed4b6e5d6b5fbb95a20667f2a7d94181da5e30344bea08d808d1f329306bb583eaecbd8deda7955cadb54becd1f77d44fc3b53f9f6304fedcab2d1bb59d16df821c20a03a15a324b6ec4bc023ae5e1a1b937fceb1632b4d4b8a8811ce9171568ebbbbf6e1aa58a598eb31abe252f6657f3ff142267e25647c8b1ce12c010c12a61d98eedcabefff0ea464b7f3548420edd27c2927eb79f4a5f8e822f2de2369b4faccc1286a7ddcfe8e867ee02eed412553a51849dbd306147dbdcf21d08e2874840dd1412061016798ab0912cfdd95c223abe030338343fa4e23afdb1cec5576efbba69cd3651b012cfe67cf8d315e264694bc6f6754d48d28183af8096f7f6963814a21e0a5c5aeef92b0ff0ca116e98741b8d4a03b2902e63eaff8c0320f0c958955c1ad6104967c84a9e521cdf345218ef5c6cf46ae6f0ec69908757b678ed2dd195972731eeb4f19b54b7f66db8d4f334f224e3a6c6037be7044ffd47c398984168488fd54452488;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1a3a015ecc9e222dc6681eb9d88f57537c35de5262da1362da18e9c9ad9a8543a2d41d5a5e1317ccc4c043989a98b35a87e96888b8e2b189621b5a1937bdd120e853cd8eef66ddc9609ebf378ee25ed00b4d104d3542aff08374f585a3319f3e401083346d75462aa3288893907cd2deb6b72aa499a4879108cf2ddd882d3ab5ae35597b87c008807f3eed172d41b7e9bcc5c7cf1910ef3dd66675a79da33810a7604200eb2887b84993bdc308779875e66aafc69e82a54e60b809978491b48720e37f1c5914c9ca7c74868f2837c3bf4704819c96714f1ca7ca318ef14fd4d417414ff58ad5c09b62ac6e5b6d23c5ed1a1dffe0c64fd9db4d058193b534f5f97dd5bbe7d6a4c2a3b83c17b6427db9324d41909a2fa3a975f49728bc9e7097d907513e4c137efa1564f132aa8eea212cfafc6d1c02f512af37b9d700b4783061da9c931c5314b1b4d1e39acfdaa622b84450ec4ec90e09ebfab0f0bfd3751020253daa6c9add40b24a4b2ec826b118a561f167d219bc32bcb888933e71ede0c63586013d8e793b510d781e90eef90088d4eb8aa2a094999b1ce21c8f855faa5db4f8c7be8e6fa258a6997dba380c1ac50b7bd498247190f91e62d485ac8111bdde12a1e80eb678e67a7fc3e83631e3f8645e71769f976c5ac86dd3a291e3582c577d9ef9583c65d4b3b57640c30b6844ad0fc0116e198c6c4a2baad5e3c76293ec69caf31e0617f7b5db11f23f3da5812e0c45d3985c4eed1d37adc1af5ecfe2b322a79f5efaa995e46218cb2e2a4420ea884b56914d26476d07ac3aaef70d9c7f7099c91875a9481a9f5e56272cf22bd07f1b68ade3c59d8126370178055967904c993e97e2d1473041ac8f65ef0ac75fe0eee49da38f6a2eb1cf57b95f3420b3b5d806a7185268556c4029626d13d2cb8c26733a0e0f4f06947248cfa21ed83890499eaa5f44a04e5018f17b45ab28e07c920232b5a5ed9646ed50a849d02e68743b979fb4ef1df3ab225aa46e0d691a2ea5c3944adcee18dd6b45ae81854954e41d56c7a3160b0b5f26cb5db48826fad1e7d93740b0de001683ec63fa25e90be57cd674752b47c5e37d3eba2c3464b044d29f29b171115c7b397bd35ac3951e705cba1c75783a164e34bc01543e8c4eaacfcbbffa0a88db83f652ce480d5431cd4fef9233429982c540bec4f60c83edc89feb934d6a041b9d56e37663cde4ca8211099650d360e93257f15511a11aa519525f8145ede9e9830ce54344e966ac8503b64d3a99d20f2186c5fe69c12597cef5e1cb16131083beb8799876e25e3b20090908a8b67c42688973a286a78989f2a16ce999cca0bf8a73227ede9faae04849808b42a393ca52eb1aace9947262a0fa5197947e4a32e34d5cff7e113336473b0d697c7958f0eb8c135cc1b4ad077b32b587fc62ac33414b7ba598977d936968e9eb7e5371da0b24bb07763d24f5528f22f2be33c24180e5b2b88e10d2fd843308c6b17817ff7998a976ebfa481d313e048f457acad680c25dc5548d3d07e0d3e2fc437f5a33c864d5815415f7a2ef9afa4990e03167a1d5fc1d3c4985d073d1a46de4cb244224ea33471a7fcf8cafa6f38da2d297b204b8df0da6cbdc2643c67e7f982c36293d5467af9bde3e17fa04a409ab279795a267d829b8d02eefab78a4e4df4642048047ce1cae4b123b2931da6217d68b5eb398f1f61295e652d8aad7bbec54ba32d9afedd17d2d94a9a66a95cdfb19c3086e862dc6cf3b97a534ce86e38966d457cd1193523a4d14dc758d80c07fb8bf6e5550a55d4aca02f4ba968f83604b21d5aea224142b14d9f2fc23fae53f180c5dad5918b501cd669d34b5d90a43b3dd0c4ca3924a447090d281c94e991ea4526655efe3c9125ea0f6064932f4e32c5bf9f7f5613a8aa964fcff9d4795d96102ec863c453f2e0633c1b8cf596d9e475e25924303d08ab16f52de507f871c6a7609ded8d37c5c6a9fb08b58c7c9c10d2707f57015f5fb3d5c332e994fbd16cd575a2bdaa6d2de2f0b9b0258ff76217a871b003290e65b862b6ad5cc7837127a75b90e880349e0ea57f8608be4963dbd9803ec12ffc9e784326cfe1bf0413829274fd9c8d4f758a8d5b7006bbcace012fd0968c8e1390bcbfaaa0cd3c08560c63f8b6a8c5aa0493eb2a597b4c458ebc25c28db908ad76e029ccb90d21cb940d5915d3ad2a1279256d657fe20ad209eb5fc85fb4d9011969034cf1ab1e63f591ddc2b23d5e170d11be9b4c9cf3e878fa4584710481afbd1b61d0ca26ca09856c8b39508db7ba67d935ba37ae77bb47ad0bb87f3937ce0fd84682a754fc2cb79d073560171d7960ad7c36307eb40298963a518053dd79f318b0049a50b916ccc547f752628d71c896f202b942c2b94abfc8654add7af45978c6c05e854af7ade7061b2a104a17e167f33013f6a0576b34e0eee7bd7151307411df1f513e64a89c5ec153187bb320d703e41e7b59029e756dbbc576fe79224b7e16e3af0f402655a4589a177365cd7e4bca21bbdbba7950f25374611160ee66282522a51712ca38d2c216937e1a1cb475fcb3860d19a1efd0026fe259fffc31517fe279257e8dfa0a4a0c143308ef7ea5bb58621210e5c5a238a5a3e55cef9c67d5bfa3e004a4ca89dea68a6d4fb11051ff659c78459f9104efe88b300375b167d0bc21d7cf5077ae6650d437a5794a43b381979eca622c68a492447c369d88babc11eecfeb378dc69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbdb5c8faebd3c0eb627235f9c9985475cffc2a201bedb5777d8ab2acedc728c05b6402cda973fa5a3062c14ad16b05963c892dea5f5525068b1d96c65df6e40623b1a11ca386055db6a0922a5274a2f3ae36f16a7ef767215cfce185816efdaa8a61d5049e31aa3099754574c7177563ec255780d75fab1ed518357867cc6034fb9039c9917b3d7be6f5b5a592bce555c88eebbd313fc6f20facb4c9b5e5095b382cc85444697d4c963c1c7bfad5e32ce1ea66b5c3d61ab188e563235cb143cb3ddff5ce63d05553918cf205110942d8530722694221ccc2ebc6e33bd9b1179dc311e44debdc31a840d5689d19ea5ed8c19f8c104d3d1453b5c85643363696a36324524cfd9427819d9357f10938552629c0154187ad3acb35806c0952576402747e0385f00c7f30ca03cf23a5f02e28f1f78302591fa455a27b37847ed441cd9e2e4e7964d091bf6171aee28c1ef0e37965fe42269c8794b75631230e98c29a92617e4f3ca58b6d164ee6e6bbb10b18c401419f8e26358b1543dc997587f2f2f332367e91d9523a73480cf18124d6375d26544705b6f905f5d8dc9742c7046951db1eb13d01cd490a3d88d7c2dd1be69862182b940336ca66a8c6adb0f151e0c524349b9e2c80bccad500d46a41fe572811d785a0b62a4e65760110ef18f245ac9cdd1aa0ed3bd87589c9eb7c42a12a46067332a7530f0114e203d0c69bc415e3178581d4b0d0c5078f498b937d6df2a2e4e4bf02ee45e9df491475ea5566aeb96373e7cc3b0a6a081f5de810f349ae5aaa7f4828151aa4ab813045d169c3bfe9a7c9a9f97558cc59694191349b1823b66606cb381491946a06700d654eeb42352fe087bbdcaa16d4c8c31f6e919e4db213a9a694f04fa3f8e6cb39d283db2d48e10906c550e1f45a404871edceea88be8b549bb42b98fcad3d908a4158fe7b661fd86ef0506e675e24dc5acc40bd7ae081c5f6efdbb4ccf7dd04bf7e258b72234a545389f6cafca4bd87c0c7833b28d811de068a0a5dc648ca8b8556611462fdf24e64be3c301c03986468bfd3d8c7806cd6ad0f94421545b0899aa2f91fdeb35be128bdcdc1d4a9912dcd0a188c6ec129e71d5ef25395e8953f28b0acc8df0c620b46df7de89b43733e49127cc5afb6ddf1e70c908f22c2a02a2acc7cbb7309336b5be5ea6758970739c56b56095848dd1538e4640de990eaeb55177b987c8e03e0924d4e2a9d245ef4cfbea1355502f36e202a8dfcbecf2c4ba4280c3010a498d84502be3995b11cad747866a175de90188ccda59d30890b32276676d836b53979c4579bb486a6674aad51b368d2709c9017025e6c96a23d7ec0674abfdcc1f9e118f4aa61d863cfaec8e7db245d4e6afd2c7f86d99b84d7687b750b72fbba569a926b466431f7d68a816b72619e700c08ea02b1cd867861acb14bbce33360dfe7b8636b05ce11dcd35da1889fbd24c11426feaaac4f2147dc400dc02a648e1027affc5bb1ef448138226dedcc8a202fd8d564ebcf189ecead7c57f01236f176b7f3d3096adfededdd9434e71c98a423722af3cca776bc9c2476c1a43a9c5e9fd9de9ef193ed812fff3ad85f83e492e16f42f067aa000357edce7e9252fa05558c7a679d9e7447d0e1e5d67466dff104c9e72d84c72aca4abeb98c524904ce02fe473178ad076cfc631f90915d1ec459346b9612694cb525884baadae5442da1752266430441e92ef5466c7ab5efdc4451cb8e70fbb9ca4c6576759c87132f5d8f2c3a614c6910d69cae54b5394d650f241dcb403ab96da3967574cea971ba6e59990a1aff6a3920285b2ddff4e54bf0eb3f767eda12dd8504017d5011e22d469e9a67e295a14d3a5dcb83cf8cc6f134068f82566e570316bc2e035ec893d901aa231de212474aa82f73100b47221a75b6019922db5d78e4c9bb1ce92b92f95b310c8717ba7cba9d4aeece2b0104779c19b9b969d91b943d57dc7623e85b1bd92209e084f7729dd7b304bdc3b1750acba0b6e6476fa030455874c2a4b0336b11bbb614cd4b6e7e9cd57e3f289985067c91639f6d701b2e5c5b3a221d6c5f0b4fd35cc76b3d2642a1e7addae7d5764e900cd00bb7a77fb0f8e138cbb55959ada9201a812e2f616a8443745b330a9384376b329373838a62c40fac59168f6450c6600e3df9fc3085cc09625e1f11798bedf4ab1cc08e4cefbf647220f23a2ffc2ba95ff2982ea406c0e90bf15904667b2f7983b73970bda4fb95d67f77a6ea3a1335a330835e3f4af529393c88470f574d2e0fe215c045cfaf57ce59c9e07c0e1de5d59be361b07ee7ed1768ec365af3f26b6e9521e26ef212153de7c511f95d631c60de26306a6016cf274460747700967405e3bb76dbadc1fe0774a1372136457c976d5ddd4bd79b62eb9e40a712e3faf35b7fca13f11582e5ac267e57d5817dd3687b77cb6a8f40f067c08a204fc846ad8ab62cfcc0703628445d4987e67c64dd421fcc240b642efa1a2a7e060325e7c961b286ce6c64ff12e7769468c6b3a910f736e630f10810713a75250e4d8d2a7ba89e9ba4e4b02326fd19cdb79ad32059605ffd7c846f2daea495b167f864e69f161e8b93e828ade451fbcf19c2c3ee554e4261fbf6790191539f19bf03125156828cf2efe70f5c4238b6bbd4024533f7e9a3acfa17a1c8eb274b93b56e5bbc7d549677c151ab9159e2537d8b33a165412f75f0c9f48c920dc43c997988b53e4d86777381ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hcf208722ca52494b7dec6d9c9908599c4774330ee86dead69d579594701f2ae22d91beff8cfcbdaf2d8e80a45075c6c102e0e896e585b51c93aa3d206f0bffdcda0b622fdf141aab1441551f9d4ad9708a1f23a0153e757702aa4923e8ed0c345943084ca9ed49a81581406e47f3cde615666ff8b8ca04e24f999f0ac85327ab6b739f2844d600ffb2d2e0b230404dfde744b0bbbe25491862123e2ae90268b8a7971902750340f3e3f13f64cfd805dbc1840fabe4fa47b404011425eee3a3136ef7ba3a3d4b77abeb557bf4b89d8b29e1ef4cca607882d4138b56b4c4ecf2691deadfcad50f0e5c5f8bdb90b8eea51d513bae8e8a30681bf197a764d407b083f04234b9fc7baa03e9cd42d447bff00959091235dce1e83737e498d73fdb14b05bf007aa0ce6e9faea17c1b43fbd54f9465bcb1260b2357674059187eb39c84dc35b373faecc5861653ceb6b0f3ab47a00d59690b538abaf9e0db09a0ecb97aede990bed986063344f1c70a9726c2ff672469b1323c9093dcf994cf561cce82025379ceccccb9bd03f00e4520212dd3acbbc050efc2f49e0b72ed57238a54bc78e5d3f11f02f49aa01b8c62d9e4cb05b92433980bec01560d1e3f27af41e18221a804517fd8728fec9bbaa70188325bc560ab7ed4435637140cbd0181fe1ecd9289e32820874b3648cfb839f028da8814763773b331009331c7b7bad3a1ea5426f4f538c0f35aa4b5f9b0e3ef6d011609956be369fff6c8015d18ae01e03530d863c450d17075823b9aaef8457ce4a78775ae5ea41ace50fd759e9be2360977beecaf519f73a352b3cc68b02aac15a8c5535b2e1835c7cd81e84170e3de6abb0815c7689bb7040cc7308d90f70fe54be418cb9e92345bde7221e5ab0b39e2606b137bc5c15939a70676f3ddf5d3e99a565dcbb8ea9fb8cbca7ed4a6d7bde5a2b387c82b1e0e49345487edd7972b065631e0e091c832f5dd09dcb14accadeddca1edc0390bedd9f0309c3b45351dbe8559a4264f68358e364d0968f8a7782905dc3433643d113f21294b25ccec1eaf1950d93ae91ec0bc5a86636e16985ebb479ae4cae9fd26d91b0ce277e5a15ba621d0cf3a2a77f7afb6deaa9a6200ae4b312d83098a4f74266636647753d54efd96a41184d63188b1b62cfad146f8effb4aa3450f85b2caf281004c2204077c874f11502b1620d8d5f2ac199411a74d5dd92c3adb453b1ac8c7ff7c42d77842eb95f3b22b6a38a9fb7abc6fd5be6ea17f4ccd79cc3952c654e04dfec708e216e5fae7553767068874bb858087edc0fcb6d50e9476a8c6323fb52902565170055e927d1e5c8a846ddb41c143ee9586b1db3c0f71e6f7b6f02164cd2088dd42317db8e7565bf4e710c1e1a950241d635f6864b813160fbaffe8dbf17a050288f7cfddcdb4d155065936b5a375f30b976ada6d6ec9d63c5179bd0e11e4b993234ec307b36b2099fcd091b24cc0a2d5af64b3f933f2ee247e8f6d0378c5ca75263880605ed6a12e91e7b1bf8b0a3af614a610c9a2ef3cedd41ab045468a77eff030d0881eea4dd10db6fb17409983031bc940d4f30091f79ea0c192e1d0fd2e8c417a78393bae162f86b39fce1f0cc2eb55ddcb562c958715f53ba5a35cb12c3a8bc33297bf6354287d3cb5917221dff4c59ed492155459085c6999e84c6674124a6c9347dc9d2205988b7181228c25350642cdad1b43f4f6a0c5d3bfdc9bee9f2a69e491707ce3dbe020201b0dadef5e19ce9c5c4c4bcd7eed0a95a5093b9f1442af8794e6ed3e3ca79a8e0fffc0a248d932e3b822dc2283b1a15eedab03ba3405cda3ac3ae10b93b31cc8de4247768cf4b9b628d1596a780e6972eee7ef9bfbe47576dc79c56bfeca30ab60f4b520f142e978919ff4312ba5b1db31aba0d5e5c522f60e219fd207b6a55370ae84c07b4249d52c9803b40cf64f7aee6a50a2fe12abee84a466862dcf261c12104ae4c2444a4f9f6cc28f64974a0a6c3f9cab1958892a13b967c5faa06321183a56ecc7d138f8111e579de9175ff6e588331c827c3946cac84fc8d219af676568a5ff06e0ed3e75849eff4e10195c0250a5b921a2b135dec76dd9000f717f65db534215abcbd37afd398b70e5e543c82e722164a123e44b9fac767dcc4aeb44a0bf66bead05524a8edc9e82956e3fe7e29246301727227381bb5fe5f0b07d691b78fd33ced523c6e58ab301417f4926fe291140669f7d87e6b6e4ecb42fb7043032237a24021e23babe3eab94bba7786a84ba4b9a121bbc546e994c06eceb54714b69fb59d7167c67d1b1040f8085fe29a2af38d338b97f295fd05fce9a45817548a3adb31b7181f3a0eab69f4232944ab7bbb6cb8514e85bd2361d1968afdf475747d661395fe1c2c2110c4773e6bc1f8f4f779c246294a6e2e77cba2c1a1ac720edd043fa164e9bd3ce5009f2ce2f226c081303b2a6ca23d5f61f11b4a1b73bb1863a6898a2fb519faef8cf3ffe9eb10544af3b3e2a23b88bd9fa69bcf58b7eb8ea51a79bbbe7e380ddad7d6ccdea38e572e42706ad7d193365ed723d6d8091cfa1c7e7001c65a199cffe780a561a476149aa6ae0538b0b6a180f5cb33e727609584e33543ef4245d63a6b39d19a26e07865705b425bf0c8abe235e218cd0251683026b12364f4cf6c0814750f45bdcf8095279f5e8faeecf095f3cf8c320011b5b12f100226d3dc5f779da025c1ba00a834e2a24b69ae97f723c57dd762;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h91d96b8033e64bb227ab954e41075b788368e1a7bdb72ac5e3f17e36d0c10ad1a00f9c14ee10b08f52b68a3e1c83814c7cd8e602edf6d78c7c5925631767dfc6e1d37af3d278ff94c62d7192130feca6700719044df6ee5c535b4c2fbb4a2888ba4d64645a62e57fcf93eee8376cb206e04199699dcebe8c89a4f91b49b34d4e2eef8b764ba4edd52031f1cac245bf577950729156d65b13e0c4d44b8e242c4990710551da160666b4d7c6eca838917cd71066779f061971f2bd902df564cd79e401ebf3d36bad4d18d3fd06141bf61ddacc5062d8fe45b96566c68fa5676016a1b7bb7a5819ce670c54add5c901c281e58669bf3c18c8339716d5ecec0a4ef65e32a5c07330cfb14a961217231cce4fc035abf1f7de42552b71f756c95a44eb538395a1d90ef0fcd598df98eee6361b8a5a88ef81df613fea9a954b9b4e7a0a87a1418dc30614c53598e1eacedbac519553410e0caa92d245c71beb9b6a3d55f60da51f2864f59538e2233d645b4ed0f8fdb2b05fa21fd6dd0a7b8a957dc86987c29369e6b3e7dfec665339f2e72af306227f8e221c874b58110bc7d3f65d85f50980de28471e8b986fac3503700588d54d008b829e938b73202a5883e5458308c932b883bc45d5b9f86e3dacf76c8083d1395bf9dabc04eed99499809f13d86902619d339a38524c2f7c5c61d93d7f170054507719000c19b0482b32429edc804087681d62f79ebd17ca87be677d155d32dbc896cad82b73b32eff419dcac3d37890d3f8f1241fe683ffa4780c660182b138080b0d904af4da2bdf30c7aa6eb5f87096900aff02028bffd010efc64d1f80acb60203b23a788d90975bcfa1e308150967185e1b899ae210ffe1f4c77311a22b2851538a57004dd4bc578e2d83b955d3986bc0ee094f1593857a2609789ca899da761b26f8f5d6a0575e9d4d6f51c421a36929382119b8875948ec15eb8894ca6a63489fa23388fe0b4c86b00cc70388974789c7baa52f985068cf3eb63c1db1b3e6c0bcb4802dcf4dc8c63fdcc65d92f455e947e36e7123e5172ad8bb29081c36009c36c112f9f7b2eb2bce92478dc184d6d2c42e05a4d1ae1bca4de29467eeb4898079db6911a9c6d5d9805f99215fa8cbdd0cb9af5f8dc05a7a851a21b8460b142b9847c3071eeeb55d6db2089469b019d52696731b53528909497aecc89290f601f739c6c8831692eb2b123a9ddf1ac579162f84b2a964f0d5b52c04a8534a69a2bffbd0d7ef3175f4f7ac43c463182c95aaed73b863e78a4338fd4a86ce2d8b8d62877372595d052645c4f11d21f9baca117f714aa4fc18b859616d9aa5c6437080f129d521e6cc8440f667ff631bd8794e241b87eef0f6f6d78fed2694a44c6b70fbbe6829b30127e4c97ffc3d3760ce31c9f97c6d0b5b33b5736a8f2426d658b7a8ff80ac08a055afbf23337a9ef4320f3604fd97dd51790f09e7a757e5039f9e38578af9073cb70032aeed9a2a24f9a0bd6d289b214835bf6fc21ab97b6dc1d56a80b0d4cf6c6e06c30f1378d05018133d75343fa915d9fa02427e8dff6dd0167c8bfe791d928b71fee288c9addcba4294d3b7913dbefb72765b6f36aa92aca9773bb5293dee2f89d98b586e943c2780c1f1423a430de1b542fef8b764f753b523c462c806eeda0d26eca1f574abc68532aa9972883aadd8af907ba21da8421c143472bd98d897b1df1ece1b6260a4fd604277dd42a10656a860015fa1f50f9b25fd78c8a2735875995bd28d0465cbc237ede4df3943619063f72f454d77309fb59fcc8d683e6dbd6661ab467e7eedfe526f2be0eec5657fc9e93e0281aadc681623fd37b29d71d43ab3867968d7b05497d55085a814f955d6e5f98821847fc1f2a1b71ff6082b8f56e5d230009c9ea2ea75195b3013bd920a6c09ecd3d729fd6673f508544e3948adf83e96d1a83f28cb983a97019941cdd353b1f00d68832a214f64560d3a9a43a1b7c02e971ee46b196e5bfe73796539f21180e0c727b928552d8649ca18a2dffb6fbb829f3ce886e4412346dfbc0dbed0ba278e8bb9d1bfad0a967d7f1c360602b469a169b9451de4e2a1aef40fbd38354888d9210e600639f747c085a5c63af4484eecc7f0b5e7667abbba527e7b81d424a8dfef17d6eabff8884dfe149a8caae6a2d09701da97a1466dcf728fb0ad8096f0be96936ad3158782acc82ca99b87a897616255972027c630d215fe0e643e697581aa39add843c9cc3b8d8d1f0a8cbdfd2e7df7cc69f90eb4b0e5df12c649c7f2b58dcf4dcb0d27736aa9f3327f135259edb776dc1e940000c5b4ed7e014f325248fa92f02047fba17987b6f47077f57ffb9b13533b0a78b93f8476cd148a38b26c49cf4c1dc74cd91f675f5531809077abbfa3098a137c86d193bc43e43ae024e96f4b020dad74df1b07d4ddfca96b15eac445a75e2e1a6e0c5f6c3711f1cf64f8982a3cf9d8c82ae4d9edfc9a08ef3ae2e8d979967aca1cda84fe902e3d18a8eaf5ad5cd71cc8cf20c4bee1de786f3a567289c83bfaeef3fa85dc85850db555e28ff6c240d8670915266ff7bc4de1dd2d505119503fa06e818e878ac6bcafa2683ee35acb018f5b12f28919b5ffeb59e0e3187260be6e2b9e5ba48dcedb15a2a01fe393257bde71cec1313e1ba444f50def60842e8fe4d5e0cc39d34befb652a3288320d73af33997b844b71377ff4821cea3f38b196e683b33a1fe846f5873240c09927c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2f4908409c286fd7de130d5f59726f34bdff3a2f7d558d07d476abbd303160480dfe51da501e9993d9447085e81d00b1605a9950c6bfef8de1202de75a3a19170a0e4118bef40c3762ac7f7dfc128a42e879ecfbbb0646adfac1a95a2e415d70bc3916c30a54e12c6f6b3ea4276faaf56f8e7f4a966f9ec8feb07600c830c2448735667189518a60449b19a2f960d210781f77a440bc4194bfe468164e859099207db037525488d6323213343d8bd45a868400145c9224f68bb81d9340f0cff6a3ace98f20f59729b3e6ab21d0a37c618519e6a8155ed793fe2dcdafbe91d967ebec0e654e9375e332d09912db70d39b0add2405911f967e96a6f257281709312f663e1172b9039b70ebe2a4617ccb78bdbf558b06fe4732409c0d467db1837368efcf24295308dd2b3a44c3ebebe7faa5e5732819ad9038d31f21adfe46f8fc55a21ffb1f5df7f39527bc7e9c8f6f48259494390692e491001447d89175bd61715aa09e112ff2e1397c87f3bb1ad3ff61576d02f8106088a742e40680f7958d50674a89e20c0273505c41d1ea295640eeb9bdb4445864a88935085a7e2866a86cee63717554c3b0abdf2f43c2448f865f54737d2d1b4d207ba1888fd881d347754269ae399324c12b9a82c1413b965955beb10f12d3e3af49d79fe7fab33dda66ac24a817eba06770988ce2322ad2ee0e71112b31639d210ee823194d872fb16dab5e8c3ce04f29f500a51e2ec68e6433434909a557863b7687f5f3cd322f439741d9bd41bc99dc26276aa9755788e56f5e2a3e9a80ea86fd36189d2c26d727099167c961a41a7e825021c5ca92e4b0027d7bdf3e4f0e3d1b5f9d34efa57cac83bca288da9bb6d1b53b557584fd0b0cdb56322b806dfc3ed3c458394bacbcaad95fe938eda3047a06a290a0d53ee54fa576dc9a4d4470ae59251d10f14f0376367e54e2481d09262c1994f7017eb1b67590691f70d195b60d8c3fa423deb3b8d53e700c6bc0956a70ff411ca979b6786fc8568f50e781508197ac892fe34b5e93f0456fda3591e08ecd438f38560bcf4c8aa4842b77e879659aa1d3f23af8e2a8a72d337a2cd288e2fbd47971e59c7b2920b5f9471f71a0dd0c5eadc8188c1ca5c9e2f231b04d7e302f37df3c88ab8d74c6339bfa762dba48f3bb3faffc7c3c79dd629ccb47c98a69a054103bd4d55cf02dce2eb4f17d7c87df623166379d92fef3580f976f87afbd33a4070ac817f6312f91d04cb6f9b3008fd403ab10e078c4bbad8832eafd72b9e5a2a3df27897b3feb99112ef0a606fe82bf2a7bc04d0f3c4db50a439677a1f2fe831fcfb1809d677d3b8a72cf7df8bd097680021670c42af4fc1287415907aea5df6c7ef625130f924653c9877a75090a99150a929412c61c027c0d26663b46576ed06b0e480b5c483013da031850bc79948118bc25f19184e81f4eda431827bd2971dcf0a3933cf3cf3c7066ea4234566c6b5abd5ada7f5d729db639273ed11697ee42ea816ea2bf901a2656218febe6cd748cfdf502a0321e6d8f18cf02f8da6f7840e3604467061cd22d76f266633bb25a8f9ec98cdee1e5ef1d774da10ef04d011af580736d013a23df0a67848fd4d84ac1372a5d82c3a0ad2ab686cd46612cfbdbbe6d7a031328ec087eab7ad03643c2abf5100ff54f818a0e4b3458cc4f2098bdc2d084b216d52837762574682494ac9c7ff0cd66a81e0a4c9d90cf80c586f9f1c2ea9d3e28555675c1f89dfe1b7feaf110b3a01686164977b20fae7b9e75be32287d98bda411e36c11d4433889c45ab15699182e826f155d0ff2a726f41c0733895200dfb653ecc04543de316c4b31f150b76fc44a6612e629eea79f785f24be92f90fbd2a9e3a6a621188970b7b8d633f6ad989c45eacebf5eaf14ab02a7e2842c36d9af3dd90ab117484aa28deacf5762e1497e6431270020b0f2c1b178ab585b32d7d682e8af5030f9cd543f6ce7feb1626717c4ba20090b4e7980f44a53aa68ab637737deeceeb02ede83a1038b3a356cba6e571a1ad9b80f88f7b275869e3016cf96077298af4b4cbe9e0dbc6e7ac385cf23849a2f47c1e9c86e327cb74f539646ca69e76866edf39957fae19fe07055338930966f5259266d7ff0f0bc5052d3c3cfa9912aebb6a7c3490c789149ea5e3da517b0c8d9e29b9ac69e02eea70fa2f83315dd0b3bd7dd090df29707905d784e91c9de2536bc208dacb8ce11ca446b321cda7c75a4a24070179085946b292621aec3952cf7a12033ba0f15bccf9d27718b48d32f05f3717f486091454828f623b2e96710710aa7a01ec7d1a5b5f25dd481955f9de2d1513505a64d292acfd615703f1e4489588b9ac7892c9e7d2235c68a34dc95ce2434c6852fee425b536983ce272cabd87884e2a0c86ca33ee819c6df7e3a74cbc4648c26243af71be0aa539234a7f64431e967641eb87df1e8f203813a02e2441294ffb617edef842ef24c4b34b967dfb1b913a0f951de50538463037d6b9d758a05f43033a0a4e633f29e07cc1f9f1113a8882ede95551624b5013da08a759f6b82812f5bb031d77f90e470ab1a278a82ebe509889e43fd5a884cfb9aba5d64d46495b6a4e88bdb319c97bf7c438e8d7b755a4a120a50b800b688e4bcdbdd6d191fd7d7df68c3af15579cd461cb1f2855e50416a1441e61c7014a3db6741b57686f9a02338dd2c04fb9c302f9f412aa0777772b14b502079b0d9ac758ff0f1d2c1ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7ae6737e940ed6c6343d5a05d30e9e72d37d8b7ffccdbd65d0781d495b1b6ec52fd06437d43f4d56552b888fb17614066a1731c778101f273bd40573a2de430e33c85abc59208df73ace36e76f946c6fc4539e584f3dafb84974f0c8cac77121cd9510b3949f6d1509bdeab7a06ed483a40a399a12b7042c78f553f154fd74c59d49609ea933a39d90aae345afc3b45c6e7e546d300e2fefede8e32502e481679ea54c214bf296127e9144a8d5da5622d05d08fe3cd85c59623801857c5310d1f8d19ca170cbde2944ad3af368ff02e67e0551b8537be17bdb8632906f16fe32d51254b4cfa4bf557289facbdcc349feac0c590ff057933617279cf3f4798c1288da68cdf01302154471d7f8886a2552e8ded24fc63662efb178feae9cb01060e2c28dc736d3e364c578e6875db4598bc4281ffac4ccec32ed1f9608ee199e3250a6d5b99bb53ea062a5ed15c16f9c8deffab6eb906f63009d87709a2d00f904013c7edbedfde024237bfe1edb2f37a24510ec5fac49aa8459e7f9cfbbba6607b94eae9ad4929eabc281006169fbacf885a7c436057047ff3bd10aa8f464ed9efff760f8cf6944f0c7483a1d2dc504cbea94741c93a8b0418aa121a84f7593e800c3372044ff9f8e2add08a31a2bcebad2a4720c6bdcbde6f959fd0a2a4affdeeb20c0a16b7ab9be1ea35e80edf654f92bf63a403c0eaa54da2a31c960eb16a1eca2a2236d286a8596b63ea463a2c2c0c5f2a799c56152a0a2536b0cb83f138b25a7b06d242151baedbfdca7c888eb0e9d8ee578e43f38c8acf4cf484c1d4eb7df58502e3c3c478b4b44d2e3e74c5478ebb4fbee2bcfbdd578e5f86a08f99be17121f94127f333a3da1b8a4709fca9eda3f67767049af245fc37294a4b3c7f67c51dc59b5c6440905a2de39153c76d6f412c6cac6bc163ef36dcb0b30e5500ebd28422d6af489a49c6b0e9b72c49e831c26b27fcacac9c4f7c5dc231cd7365902c80e59d713303f30bcb9bcf4d69ba831c24c71afc687d81f2ce2df1b90e0765958fe2ecd89becd2f1b369a384ecee77f5bb6017ffe463395716487657ccb5f274bae6d86f54e53161e3fa1e203c8bdbcebf0f0ef0c442301e8f9c7dcb86b62490b24ee2e183182d4b5b1981a0ecc530eae690638850f0c92c1d61e97b4ab538c1539f95f25ded3a47ba2ed427ebfed9fce2cdb9675d53146c1ca7148a1f782fc3536297436c772fd6d2a2f62297c03b3ccca847a705b8bbfd25d3790831bd52299c301462566bdbcda23b570ff27c043c01219518b6a8b78a392ee73ced256698691e9623c893046264d2440421955dd92fbf90ea1fd3aa848a7773cf3bf52c87cec9871cb1999b969249b6c1f0cb88440fa20eb89586acc92b2950a105b8f2f3b792818f2b1272ed2b1fbab4464df975175b37694cfa0f1f49934abff7c10f3effb6483b79b2fe6c565974d566f622eb2f56ca8537a0d3b36b668b7d6d831d93ab760e05d203c1186f7eeb7565f1f9a2d35a5edebb7fba96058146b7299f942c13ea9fb968c827bd43a946b5c22ea50177bdf9b3416f5f1e20693c580ebf20d9491ba54a5392b64fb28d2da3858e1ce0d0f249102f05c14bc679f7f9058a9cbc8edcba98c2f27da48c16eb53a30e9ade976dbd6ad134ba8f6f7f0423d00a104edc2086d664866148a18b0c4d5e0095880190f493291d66f54c5621dd801c8b6a33aae45119696a65688e686db4f0adfd303e72d4ce75eac29d129a3a3cdcdeb9f339a8ca7087773c8fb539b0bab5698500f2ff4a48c3f62e6af92a6bb2e10b69f874fccde9694043b0f97302c1ac7c80c8e91faffbf9a65688d395e70478f41ad780730c37db301c780ab08843dacbd9bee8ee5303f42d21d2e65089a803c81f63e730e1db031da6761a3a97a157c577b0fd64d1e22dc7999b227b429025c1956321210d2a58192cf64f57040a559d9ffe8548af9f12493858f74c0ba8071e04d1eb8e1a4bb9a793b2b10df45e4239a50af1d500f50221e842ddd2b2bdbe198d84501457a6b9bebe6cd4418fb16cd1e0a627f946945a0355fbbc25f34e4dc8e7f5fd2e40fe04005e3807cbfc45840295bf20dc9c03cd2c266f96d745fbed459c9ba9a30458d75a127bc100e7fd39b8029db18132e6834038031851166a135dca89397a76d561d5662f0093f83c00ffbeb193402675e0cb443ebf220f239ff07fd07affea5a1cc93fa693fe2f7fa3314f89cec446ca2acd73a658b593502bdc1bcacf699ec143a0cae85a84a1ec627b002a06140382d831aa29ff5ad98cc9b5b70bf93a4e2b2ebd131c06078e73db09ed02bf0f80b513bf924a7c2fb977b42dd3285564596fe594e58565748c90661b55f6bc0640ae27f9faa5dee8708e243af673021509c1074961c4203f816761b968df0635ff7d1c6122f529010f2c1d87385db6a3a77030a1fb61ecd6e6c7688cd71a5b65c104a03dc89dce6be462a771f2f60f5935783502e7c247ff3d47fee59564080c6da3c1b087ae5bf39336e26972ad60ba7c683ef848223887fbf8ac81484cd112c8ee99c74e8ca4d1972886ee3c3e2267438401d73c5668531e6c4c81cc092cbcf9c94b56e84f082aff1654388d7d48eaf4d6ff47e4ce5638b34717844d5033b4874538f0e86d7291734438833db3a6c5abe788bc464435091626bc60941b245158209a62efb5e2d572077434fa40ceda576aa36891f9aa673778aebbc80851cbec5a45d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2a0acba9ce0a67c247ef4196caea269a0a9abab361cb7420f91b869eb10f05474ba66478a8ae0b84e77f4ad1782e41b6d84bbde2a7f59c362d4a5b58983c9ec281a635062f716e0bd2e0842b41a278a137e4437fe69d1709107b2b3bd055dd28929320d1ebeaa5e5029fbcbd2e42645c988eed5fe12bfab24f619ef12ba82ef95d9beb9212b1d2750a150cbb693fe33a0fcfe9bcdb39abd11f7b41da42439a3ea93fd81b9ee959a02d3aaae19216724d5c1eb4b7d75eed64c8e24d28992641bcd06604ad17ed25610db94bf6ca111d68abd25ebaa57ec124de2e41c2db6f2f4458cfcfceb1316195f534f2a54ccc0f6114d582b839660b4c17d353c6e71e2a8ee75484387223a1ea9e157729ac6ed2a653f3f49b277acb58305307b8ce5e2e3ad621f62873e5e976d0d963b20c66f12b1bb86bcea14bc1e84c13338ca7287e1b721c1f79ec7861d2a182fd7f30ff0a6d4ba64ed8a4b369605104a6c4830bba1b5f0fa732bf71f28210dd5ce37b6b693f00c6212e7a83849cbfde7bbb67bc42982489b12c1c854ab7765c75735c704e87870fde18dcf3ba0869682be943884ea60e43604521d282a155fc2df671d34f927de4eff0213b6e2e78423f37c3c76f6baaf845884857d2321de6eff99055ac08ed1b447aa539a9d03bb6d0638a705dd2f93565c0009ec90733c1e1fb280a754083e25298f37d55a5c39da9b4b31978675dbd115c98cc774926aa450d6f3a527dc2a3f280596aa48ca8bcb9458f515bfcfdea9f9aab5c0974b84b09ed6ebf07465e891f8ecfd839447f3b021d96bc11dd90044874f912ecf3120bb32fa01a775c0c5b5efe9d7dac031c03ce64c41f702b65eeebafefb6e6c29575a40ff10349bc349405731b5a79f655b8aed43979574bd0f3662765a6c18349d09c1e9a8fc95704343e023b9ac67d363664905482ba11b2e98c90e98d1998b9adc6779bca0ef63bbaa36fb59f8493c69c6e9b6082e010690bf6267291f4427325a89b63f20e0cbd12593fd721479add4ff67e9fa933a057e2f1762d2f6fca09e21f579479676ae6272060dd63a27d5b0171b793f8aa7957f20ec53ff0cd3102e89bddb475db655387587984aae0b6f38d3da860a8a6b6f607baaad311382f6c4afde67b74992f63a6aa0776756fbff30758f9d41ec26f1b24209e10a0796fb938a8a331ae3b47b56cb67d48d021ecc108a26b1293ad898cd1c9ed65a9b730fb3330aa4ba087e8ad2b06c57863335eea423e52d6fcdf7b6aa4ec9606dfcef5b37ebed4e8edb3dbdb7ce246e9273c89a60acd7d6a2e321a2835b77cae44dc333327e71513263da4749339c9bd36e59376f23c14e66e67633764ff48d254a37676073c63fa816c4252c00cc1d4f89ec49395a82c696ecad9e8a7c0bf5b265646dce980d3488f0c71c97f138d51fd166800d963fc04fc38b90213ce7aac24b9a2ee5016f101131f0214c61aacbd2369bb577b75faeeacd69eee4ea43e4726f0debf5b3f1e09ff5f7caa0843ce22ffdd87d4ace34fbfff1dcf068929d536d2ffcc57fdfa507c788dad3627fd699e91941be75c209ded899dd07e393cdce9ccfb6a2bb16333075dd851ac07f5e379a3ec7a5f58ea2717bfc13b7599d27ae343d68ddb5c76bcabee93f1bdece636fcf84ab0a9e510c8dbc9623104d06ad5a336af9669b6fffcd70271c0824da1c3a555f885b5734c3f01c6c1184c9f4f3cf0636659a18dfae659758c423ae31a8e8e9c38d0e67bfe03d872b1de1955d2240d3f9e9b1de3c2c70b9793edd61c55b776d36cbf74abfc7abf7649816d06f2b0b2d8c68e16422bc05e11c785daa99e0e5c790fd4e8c24988acc9918d505f04f5cf3ec85d524a446ecf13392b8252bd933bfcd1b618b38079c9cdaf75dee4509400863d428009bb012a1f7ececce9d2888358b3671cde875e8a44e214ef350b34330e3c01ffd25e0a068ddb1542080fb28a6ad6e1ae5d49a828f7ee1d3da416152d39d63cd1c4bf73645e5a1f6017902c00a419bf75155fef862262551d3fc1da32f75c74d3a0806f003f14e2b0c541ecce900799a464b413083668ba5d962899b90c29ca12490cb1dbcf91bd3044c37e10c739f525d598114a8bc27d910d8a33913b9929ec98b5249135eb156c7e9d563609e33469832b6cf0d64826b679c43949f8126b66a078cf4e893461e888c734323cd23e11d892e328be0413083d3f426ace1a97b6b71ae08650418a45851045c1ea0a36c9121fa0a46fc985f9db76e7135032ff1c277718d94f24ddcc760c87181bbe9056543e065ccf455726ab9f03d6f6a1c8f13cd97f06e327be4f8dd6fffcf2c655ab955abef8ffff497bb5a3ad5cbfebca6fe00dec5740fc0a2e4c0800963004f5648207f5815dd6866ab232066cdf646ee29b2b22ee3e74d0efb90739680779af933ae6232be93d193c6b3c2780c8360dabd06b2708099a29edf31f525b0c7fd2f45625b68bc93006a4ecefb4ff5a85d257e516672c60ed55aface2224a620e4ede54d48206e690f4148b7923eaa33d0b6460c24e61f47ff12bfba657a59967495b3255f2d7919a95a8066092c29ea17c39457a8dba04b0105ee6c7c4aabd2d58afe57e944da0f99c1713e645586ea91536ea54d61035e5d763d620790af7a410922ec78a3ce7865b2405b9477997f88dd42d2a6375d5160f205eeea872efb697a4a714030634c72964b0ba10ef7d26437b5c300410bb9895ccdc8773f57c7bf1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h31cfd0987e9e9da2f661ae3d3e5fd754d925bc9b6d32c5eb38d1876e5ab2a4e6a7597e6c0e8421372194d9ae4999db983bb3a997bddb7cd333bdd2f822816f5e1b7a5453fea339c351ecc81fb77fe4ebaafae137b70a8e3b2bdf061ba659a15d3339cfc9d5b6369f23d3a5b8cb1463fe31b019e3049236b987d597a3e0f036c5dfbbb73ded63fedcc1024c6142b33a319cd82510cb9183035df5ff2d857375d486f89a0684f7345b838a362fd97623225495fd57e35add9b9d356c2aac7cdf280b23ae084f72133d45801714934fa4971c9906600c83b59d97942202c7ae830e54d49db9663028d67fe1d86831774d51ed0aeca36e6a3cb42354f1a45e49dd7e421c18e78ec2ca5a56648024def77eccbba1745b209a726f6b171f1956cfd163706d81c2c18bc38b0ef4775961a5efc1731afa67a7fa506cec730bb026972f2c9a49e22d9a10e1394971979e4a0644d2213a1c0a31ef21569f16364ec28befeb821ce8482c2dbbc3faf99475cb8bf8acc3073c2eab0b3fa6323d7a08cc7a2f03e2a1175828e0f1fa2204eb36cde6d5d5a659136721b60965e26f9cce95b39d4366a6fd616c13f6d374ecdad31346d364a416a2377c6e47accbc0c61ad6ef5f0f9c187121eb13b36b3b47def6b09ab4858f305eec2d78ef3ab9a191c63c5e16316cc94cc0948d4a2cab0247f2d6c809f09d277d017d35a949897e3f3dff39fc098a231df05ffc6e112d6c4a8b98b1c901e762b78d35c20912c01d85eae676b5dba8cdcde44cc67d89307189d4fbcaef37fffd96ce6da9aaaa243f3a60c970b7e78e153f9059d39e75c45f6415865b54d4a1b446a36b38e5abfe535dde72554f3d413ae1c22c57c7bf1abed5d543ce2d8016cd68b8957f4999a68a1efe857ba47ab1059b608a6c7b33c187db35f294676d8bdfff61c72d14fc56d756ddf61007f915dc71a605ebb9c4efcd9c172893c6ffd7667aa1c8198f9c608f80ba8003969e3f36669b81b79129a6696a4a673609df20b2f2dfea37d47ec56f0092b9a74fc422828c7b0ef2e26ce1f3b32fab48fa465fdfa6e4d9d2ecc6a8a6daa74ab9ff66297f8b8783691ab9959ebd8b677494ef155637d0b80fcd8024de086a020af86f64dbc7a9eaa3277a19872fbcf53be0ecf6b25870664cd9a5468882b572c7c1647de195f7b318fa479caa758eb09d308c93d6be9e9ec45b134f7736308383e3290a0d8873b0e60a8c5f0c3951c83272934b703991fa178f69ec767a840b89ebf8525b2e3d80f1a8b0f01be72fcba2867378cf106ef736b51e283591b308fdd0b2733f3ef8423d96b550a8a0d9ff5c631730d04a391310479999dd41edf9a39aae0a42c19bb89098c8741f936f3a001067b8932f189ea5baadd6c4ee3284602e731135d024795523e4a37dbc97da84786b6aa74daedd51c5ada4d4f2f418f16df4e71ebb9e2741ee48e70f0ce2e530b443afc9234bfa7c66f9d4dd0aa88010e1ebe7c121ed753b42c9d013c5dd9951a797faf4e628bf7cf7bb62333a8ba34712175c9e5fc39733e77daae84428791be141525da6760f3db7a5edf9d249ecbf3b94d28b21cdb0ce30e60919f620f72c01d29a46b2a4fb79187453e66780476f4476f32dcb620a5ddeca7402ada225707f2047bfb3f9f2c4e776ce19458ee03cd702286f148aca0089400a78e5fa40357e76fe98832c0f692d08d7fb90c09bc7c443e2ae2cd5755099e58165bb068e3f061c9235f5d481b4ee550df65fae73d30afef81dd40966cf3ad901614e3a93bc6fb6c1b83787f3b6ffe36d78b8a94632a62678bf6d6266e500815f54ce89148d882b4682f9339818455f21ee8b210bb9b32974ea4cddb6aef12ac1bd4e751a9f4a2e96ee0e148288da7218f99533ecf7553ecad396376197efe237902f91a084a6cd0671a9b44cac95f12484df624a738bd5d4d3759b8ead5d606cc4aa1d2107854c96df0b2d91aef3e2831517ed76e30d7e2b58036b90cd550a7640c58dde8f0e4d3d1db6ab3f79f66a0613f5a13eea31007a966912b57aea815e9adbb1ecd67519ae84f56ca2dc13683b2d4fde5ff1abf41dac22b4aed344fedf7f98f45145cd6d09198e8b0d6f623f0f292e82fb7587e2cb1d302be0e978c8ce98622df556bb1ea1cef3feff58f4592fd32a825987bbc5926a131bb85e88534e78f952805ffa86cf9488699ac8fb6e4d8d6aabc942ae27a88b93fdaaa6a1b05853349d6055e6094cc7e3a63a1241626fc1eaad2245153ba300e5219cb0cc7280e2a5c7fcb880007dbf15c1e7d20072405d888190a8e2c1ba9618134b8e87825e1e854d4e086aa899a0bea43d54872ee8f7f7a06f9057a5010bb35c2763ac8a90921973cea002818e3800a4211e85d52481cdecdd13ffcb724435bf1ca525571287734fa5a0ad218e3a582d7cf99ba2ce2bb105ea82c3257d730fbbd05fdf74dc6b5e84985f28a445f03a5552a60b72b79cf1976d4b17e81e1d3dd81614bcb726d7e525454f1f54e19379a143843b72a61addd4f8c1f9290a32da2b6a030785e725a47d9959faf779a5fb880382804a551c32ea179ae815e5fc53bbc965a7e2fa8601feae436b59ac9bee987641d0fb5ec51c1fbd0ea270475f6821c8811141133b5da77e75c2e753fe05603fa61349373b75ccd014465d4ee65466898c2066f1cf2dd1735a75ac89b43a965cfb1f4c8fa8ae01df038e857ece5b1b10aa44a871b6a8f2821b4d393d38348d6452139a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb98a0091cfebea51cd11ab20723c1f606e5b792d5a9f79811934a1f9fbe2eb317f9d22eae8c4aeeef1a193d4c8c95f88cae9f75b43dd8138eac168ace23e0918ee11b86d4ba10096e1e04af023cc981fdcd4146e45bcfabc913c9f47fc7d6e37dd2c3458cb75a58974c22c4d83aafadccafc36c6d72943b0f1ba671fd8c6cbbb21f1662e0453d1abda83402440a4298636b59dce837afbb836dc3b334cb97b84e7c1fc86eb0f480c87197eb20f25e209a58d2fd8c8c04829b1bb859fc89fb90acbc5a2feb84c05107278d36195a917ca89ae41768022e31e48cd6e24c51fd0242ead9211b114c6efa4bb7de3c1d9910ce44c95ad8006d998e07ff6d36de10a6f653d5a14c56cebb957f923d36c8121d7809570d4dedbc9b8426d0046b0447bed750106d6791966631cb649340f56e1b5b934e41af55bbe5343242e2b8216dd47398f70a63c1a993759b9a106e79574b7a73f9fe811c9c1512401e1ba513cd5363fdfce97b5ea3f4940191914d55bf6dd3c9cd67c688a9908f54ee9761138aa1fe69affb56e718677d90fd22c79f979f4bfef4e951e6cc8bd6cdf8a8a4a9ff525264a7e3ab62e9f2b83d0ff30c8d8ece0207f1f0583ed3ff7478ab07a719166a513c94d7be9eee9a8d8aa6643ec58624d7e39fb354dde3d122db5ce68b9cd70dad24a65a87bd1d99f82e84665754df67bc43bae404fff1083077c5fc2d006ace8dfe82eaaf26b8a890b6ebdd970e8ba2e48eca2959f6a310e4718580aac9f410f8a7beb72a68e7f1fb374fa46d600f444156a60a8beb2544944c18c553587847b5bea89faa0eddbe1f2d77d32705dbaeb5147819b4661286b5631bbd0cf252917e2bf7fea1dd1569467dea8fde727440c97b80e5dda52afd379f34caac673bbc293337dad97da9c21b7dddca98555d2e6fc8d42e11a1545fdb4117a27a9068c58b0e85f52d78f29fc467b698823a4359293ed89c15304b768355e0672e3b2bbb9383554965ceb8ae7d739dc53bad7e3544a578ddd24a7600590c61dd2662d877450e00df02a685c405d68908eeccd172903679fdcf736931b7647e52cf8b7b1cc9078ccb3552b59e14b7e1c2cb161f3d7278f52a574a9e79a66255ebaa1a9895a6f7f8db39e32a44ae1871ce19d3481770865bbe08373042fa01fc1337ab7ad79f451f50cc84d908f02e82d23b2cdc4c02533bbe2ff3a5596ab6b5b9e81749f8cb0927158079144b4628b8b1a76d623ea26657435abd61c3ea9772ecfdbf448ea02c9e505ef5ed2f31b8cfe1b222655184eb904103831248c4dd7fc7155041a6be2c42a3e9365b653c0813ebdf880a867ab088f140cc993c6d1a366ba9f50e4d2c562a6656aa73c596b3cea8c1d9a4800f4df34d5d04b73a70c6a24c6026f20cc6777a0a4e5fcccd9f0fe33cc9209410883fe2636d829729455ca92a0474b4ba9a17d74370ad67539a5d1f48042bc859cf0e6c8100c74df6be0ac2660b090c7fb5d2876616f8230212bf249d0f4124c10c87dc9726801909c3d7ae217cc9d816cc792750dc93b8652faf54c060140c6f2cdb91c8507e0aa27d2084b68d9b5e939819277e2e8c0caa9c2495715d68e18f5996dbc49f5ef1cc0c20d9be01bd9670377d9556eca85898314e8a452c18f99b70dc323fbd602174a75d6a1d326f6cbeb101742d9f9c3d7aff5b8d138cfbaecff648d0a06ead5a1b73eedbe0717b26f071ccc47aeb8a90e37ee4f77f5e29fbf1a575348b62a498e33807948c34803158826ccb82f5e194ef91619a1bb181852f38f1e01fbcabebe696d4e865563f3a680f7403b1a560361fa7bc08deeea479510090b50346517bb93a0e2849be28e5b8bd67e7b1edc5571e55c08c62a4683674d01e805e50ee2d601b62c30a71dbbddea940360c7debabb373364dc2439e440cd7f621e936bab45eec8787ca0c63cca3ecafd2caf05cdf9d63b0840c653eee5e41775557ae468785c27a6c58611f1132e7c9229eb467d958d7f5fbe09068064f79792a8bd82fb3310ee9fd8db2189d1c68aef415d404f3c55815033d6ec9fefb9ed8b80c605f11167176e5a5c05db70fdff44868127cdd884d13431caa7e190c6722df47ba42a8b3e04dd9d874fd9e16672ad9e8d5d46fcf164b4352cb531d99d694745967f900b764c159db73d8af05a9963833c47e7f82b8d46bfc9c1aae20301c09447e84f34b63409754c9b9b25e1e2480d4a5e960ad0b929558acd7a5789d7b4b2a30129157ad95fdd25d84cd28c3c7712e12b533b58f70ce05a65df6222a5d3a8d558db401a4a0f8e8e97abe116ed8d7248faa8de3b067b797da6a92dcdea14acc31ffdb985bb3e5118d1670e9c70a9225960c320e9892a24886a6b564d3079fbfc4e6973ad810b8c8081132715b2eb9f629f60c82d6587fad93c499eb60520388d40c5cd82d265ecd5957740b083e6a6aed3a25374dbabec933356b81330f6d44d723cf5c943fd5f4a1935d267d77d740382e1826874fc1b0d8319342427f39870a313277bea62e1b08ff0fba677f26fa40c48019bf2e0a43b507f87b3b6a927e82526b27ad7d646726c7fa7ce4a307023dbdbc97120d6d91bdc7f62bf20de7d98ac534f9577152a1c0f18a47f917088534aaa5395670abed24642eb9240bfaa26e908a2047bc92271d1a3110cddb454df11d93bd8943fba8a3c7538ad94ed47f63b5e900b40b09cae9f2f1dc491ddae4e12264fbf028afc6b7d681f547c33494cfec7a608;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4068b907580e3964ec130029740d56efdf5fe002622adcb99ef0678bb0d3fb405f08e0cea6cc1d061b058f361ded3b346e94046406cb1915615db1ca6c63817c00c18139845530cc748d4f06b019383c478c0483c22851e74a9f5c127d9063af06b772fb91616202f7e7261f37e5776414a36407aa6b60fea97c65f2644f1c64f978d71a12219393c791975c75c44e518e4818a6f2c26128302c2370dac88f60b6ee9915b599d61c40bb976976ece3f1ac87d3085e3a36e51a1ca771eec0caeb3b71f85c5e2ad12d5398f3cf8f3f7ca884434655489af06f55c787908988353b44988eb3e3a8c3544955036349766bc602a3d155c74f491e914f6283ef9ab49ab37277fb638a0b71418305cf3a74daa265059ead5771a8a4afb61fdf35fe93246ed5f8f0dd37764d33afdcc23547a50f62103e4f27822ed00017a39f42a2682131bd460d0679ceff9dfb63beb7d8383b4ea15b3a64c85ca66cfeaaadadd5d461ce1718629f30c30c85b1bae3c10476079dde7f33cf0712a81e68f6825925b687f9ea3073bad62275fd92d58890f172174f4fc49ae4b03e29ec7e15a7480ae01d09930ec7829cbc446008756525b1728ee9043aab201a7192cedbf543d3cdf43189825dcf52e00c41c62453a67448cbb7101933fe919efcd314a34a308abd35ccd9fa95fd209c28a17a7fca833d772f81a2bd4fc576b802453420e41cb633f06ecab7e00913bbe1ce0480b139f122ec0866bbe8c6fb505e76e27e1c317afd2ad1a0548f971fb19a91200610be1b8289c3c26a097f0bde7b7eaa4605da10f863df4ec9d3fde823d7782ee7951ff0d32e9a27e2cc2079055b9ea9e02ecac1a25c8a872961611a19496ad60a34f62eeed7b237c277bdc665d9b97e5ba8202404b3b9c8853435805719594f93f33d8a041c0f4add65adcec90867b465943522cacefd08f0a5a3f3a196e56da32e14ebe535278078f18b695fad854074d4ec877e8e5cecf95ec9d16dac3a2ee0884646b02723e8b930c3f8979021c9d9834ef7da655ba5e033f3ee015526e2d865a177c73244acec2b3c8745e2fcb24139918d4e05a01bcfdf7de4f2f2413f47b43567ce9cf38d6bd80331aa23c9cecce1669d0afabebee30192232861e7553f18713fd23bf5052b7682c52989255728db94069924f248de0148fb3bbbd8558833f1cdc45847ae4132459034220293a9d7949b4434bc4b7acc78e321e1722175416b58cffdc209dcf779784eb9690e933dd739fa29479a23e02292cf0b395779d75e4741f072f573c12c1f628631899bad21e306a16d265f7c5f7b3c3c43f761bfe8835fd85bc0fe89e76900a7fd23dedac66ce7be9d8295f83b36fdb3455286362ab080aa82f69dfc8ec515ae2c5fa639384da98a5aea65b3de6e83c9fe80468c7572acbb0d3943412170e37fb8b48437ecca8f9ded1f7db007bdab76df84e7864b7c8b429b3a3132586f7304ef0348318ffcd89e1f65485d5ea48fbfc3bb3b76bf511ddc2d75637d8cb9a7cde9d51575bf320e6b0ec96d3beff29dd960fa0ec82e83ac7fc6107add545131c58f241fc4ed49d40ebb21de88d5b5734ea335c650d194b7c7ae33588cb4a20c220c6395cf791328fc5db01585906d8647a1d16227bc20f354642ad5fc0c9267563ff882b582023107dc6cb3fda43f91570507afe61316cb06fb310cb90d1af5841850d0a1dad7cf36a6b21effd24bac8d9aa2165ba46dfcf7ea3bad372267bd2dba67f3f3975e2f5d860d5c982f3bb119b7f6f70d2bcfb9725b402cc9594d79c8adce36ca0ab5684608ce2da7a2d43072966e7a210c3076dfda7134f948356ab0f11857ff94100921696ac9e8cdf6d45baddd4c3006dc971d58dce4d1eb3e61ff572c30db94810e0991401d52402953aa4f432775e0731016de1f570c7fd4b50c3be8b3eb8521d9f9e342789aac129a7cd75f414407465604221b567c95e907a8eec7cae23ed26e01a57afd72efc92ce4bab2b3042867fc4647ef4f4e1a0c770edbf7be90251f31a71b194f86bf64f6ee3ea25c20554c2d8ebdb0816e53399f760c8d62e7aaaa4309092e69723ce1205076fa8236a252764bd83fc04bc54f25aa2501c484bd7932121d1781496b2c9ca2e440ec442ad67c203129ae05df53c9c87b3eb6724e465c2e16420b0c0e76fc089346150adfb0b4691e8e69bbf99eaf71905a7723db211d4ac60dc9b5a683062c33917e1aec28345dd5dc77fd17525f9e58ec2fba4b0603262486ec8930d07751c26c588218d18a6c5b82266997504ebdfa0689001721bb1e9d871bf8210f9dbddcd08caeb093380da056d4ddae14c28161ee6683acb4bc99931c8cf5ace9f271ecc0916f43e242c61e13f450f8267392ec0136277b16656c867bd0c282c846721bd65c24295c13ca0d6264e6f1e8079748cd98d8744742167d3ff88c5a9fec36333306cd447fa6879e67c669f56588ccba0ede75ce0a156f8ab2ce8ed6df999b6fd56f2d56a6dafdb76be4d083ba0fc2da57556c06e8a3fdcadec2709d8f61b1158e3d81642abd04762023a02171a9b7ab4d5ce873bc2d67a94cce3e17f6d7dcf1e28c8c43eddb461645bfa698ea92fb97aac843213bee7f5b31b0edcb5b31f3ecd1074cadbea23fa55c4b6171acce3ff82a04620b78cd2139103660e4e9f2ff74d1454bb4aeeafc068129a7347dec0c1a334e2f486bde325d846fcc89804c42309f0cbd87096ddb6fbc770552f95954c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he06c55ed903f099545051e22c590a4c44dfc0b7febfb81d80620bfde4329f75305782e45a0d98818cb213b0cbd0081a32ea76c57950b7a684e2a047fa216fba195f76f3878e5707744b72033d7d6e869a8cce276339306b14c8fe4f6e0c043b55aa5c3f8dd446816eb4486aebb0fb61572462ae5d36744f7a54f7efcc5b50a7fb130cf72da428e4e6bbe269111b688c6ff94a35104182d3f41ca4d56b5c27741b206c1dbdf4055a3154c012dd6556b7f473cf346762a617aeb2c90640894126eafb12473ea39b0d0fc34c6be74da319a89e2b596a018cd37d0d02b18e8487824aa5e85dc6c05aea2f851984d60698a2ef3831ede3d9497a936e31b7304253805bd573b73a0effb9d345722bca7cd514b56f1c7ee114af243587094866f77d28e7356a083e973e5b2646e3e4d0dedfb5bb4aadd8dd28d5376edcabd6b8a14cb0af5ec15fa502b1b6a2266e54956bdb317f939c15f78ffe9d83a2b4255a5f00df40f214c6886396043eb5550c21820bbfd6e050cf346e95228483ca84ac99ee6585d6ab472bd5017478db3f1becb2a5f63655d601d639460cd149247941b740c4b53acbf70a2877ea10c8c9c4adf404da4859a0ba0a70392cbcbbe3473a1eb388393843a9cf0f814ccd117c5e62cb720b3feeacd5a4e1ecdd5565080be29ff61e820f6f95ffa95503fc965c869701a4678f89f0dfbf201f6c1ac8a67de584387eb04493f47a1a12b0275dd6a5c4e0f3f7e6e383709823b39a87c0eeb6cff556cffd3ef958e64bcfac17fe88848582760b34d76cd2e85510d207007e2a400225d255ac4dbcfa04e9aaa591d55eaa31e8eb4fe46d4cccee39e6df732db0186427798ad45468ddf5b2d88a5cf28ff8fa686d55f38b6eedd0cf02c205c75a6389ab0c45bc0e8a74c9c94c99a20a35f1e43dab8acc79a2423214c5cf66d59bd28018fede2624ac83f4557ae9c61630d4b13d5a73a72719510dde7f907315ac6b8a1e13ca9bdddb5f23ef2ef8a1b3cbf02f62eb9f22c63182fc022c4d5b623de3b1d32289dfdd216e3c0079ac96e921889da2323258713c7c5d6dd95c431d7fa3620d0f05b73dca364fa03e80260075902401ec9b8c5bf1d1facd94d3a9faf3bbe904a98e1efeb75cfb9c07ee3cdba92cf33dc151fc04b595cdc78f17362882aa711a296d3d5f5755cbef8f166617046389cd63ec549470406daee15dd2e94e941565777ef92d90c99cf42d593e5bc4fd73d9d2517798706e7c98dea09b9f9986c0818edccc9d0c9a919c69a694c60511d1659f275d88312f87ee5aa2fa3b119cf6a6e6893a6e34b1c4e0b6905f2581c2d75f5a11be9d925221e32d9c4903f10c2da41a4c7f499f89aa61f85c52dec9e1313e614d9ca86ca81374ce9bb9c6876cf3122a6de9bc1e35b775753e9d430ac3de25c23eaeca85acf116b97217eae4ec3e32cc8d3248c4d0256c2acdb395f3b249a295eafa16770feeac47a35aca6e6b32a48bd536b978a0273f6c958bf5b1f4c90c40c535b579c2f6933db6e645ff415dcae813c5d70ac4873f966e1c20d2dbb2b2cd012521019d4805291279effd148cda41ec1935d83bbe0db1417949d23a8eddd7ec8444a05f9f6e99f5ab15351a90f54d8a63c3b1bf00f83aba627037b7cec94888d70ad2c0798301922bc4a57cb5bfe29b1ad3f8d110c213fc83e3cf62becc2d2b00374e5d6c6056ec358b0ed8aad0ba66451894f956b077c9ba7ff107d0da458c7fdbec2968b2169884c2d132b391b91c8ab1fb9babcc18982997bf23b675fe5de3b544f16e1aeefc5c814d61302f18a984fa87ca70225e64d8ee28afae557756068c506d8b8fcade9915fc2182b82e5d3848a1e40d917de829e91e317a967be023060383d2781a5afc7ef1db4635a432cb307d38c5cf3ea58865309245a77415a44c2cc4397ae74562fd10f3552f105cec73c2369a6462cd1c40c880d545ddb7b684493406db05bd47e58b434b89598ccf9cf6fda3b179c5f1fbee8cb6bfac012e121eb35c6ea22c5643458422cb966c9f76fd2a47794c6c8e31394abf1b71abaa36e654c76f6b9aafa1ad2e9b1d83ac799a5b30fca6322d12c83c8cffb9651319d87a889cbf24624955ed7c51d57e23619719dd86a8b503e16f54fb5df0468a7322df2a5c7580fd7492ac2aed1a8c149d645c9afc77b11178e6ca9de8ecff960f1feabc5e4ee1b6abe3663d0208e3ad7cd6c3cff547884fa734f9bbe5f946472ad772c4a7dd21365f2ad156c117de01a819f4d8cb5609b44355a5fd63dd3e97c2dfb4f789dbdd5431fd35952d3a647342a9507e6e1c74104ff5cf9024cc2e7942b88644f325f0f50aff814daa3ea85f1a9c69f768847d465ebfb3e2f72055cab1bd25551db655d6d9cad4005fbd7bbad52c91c971c1d5e4ee916efa437bfa940ec1766c649bc6e8a6a1987cd0647f4205e6b93e2ab0cccf377df4c258f817a4475febbcf23737486cd6bf8ce7068ea22902790074aba96ea3bfffad2f2747c34451e8f530739352f7235a36af9a78bb796bbd7c1bcedfc35d5cb318cff39b2f482cabd088f99890b5fff3b8f4bf506737b439e31dee87f4f704eab4166d7e14a1ef22b83eea853d4524043c404e184749f828fcc634e4af5d57e0f72d1c77d4035f849665fca0a9e5ca6107baac488bcc9ad92beaada4384356fe7ef2d62c82c97dc74990720fc6a63d2d3cc3d8056ae1d2140c11b883d94559825d3d5621b9b2bde0a9b605cb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7d7191f1f72e0349f0bb7ac6f8397165ff7b11334ae2f83e86e6057b6ee447ff542c0127a0a7657f7bcc8aad19bf33a309988d39d2086446aba9b676edf2de4f459163214a33e1544c63046c4b967bc826deae7f092ab6707111fcd20351ca9a1b6c5ab9d3018c4f5ba1340d863120fa6554caaa088be63234b4072113a52054404465502db764e05f9d6dec85c5c5bccb0b06eefa1f9d614a1a8b41dedd6c6e5a22e7efd575f68ffc01988736250d9519571415f82e293d48bc4413df32e2b9a8a7754bc90763deac80e891dfc98680c701974478c1175f0c23f2ef0719847e557a6567c3639aa3a5ef4c71f944e27b33a9f25cee8bc3d481396025593d4b62775766c5bc4c60143ffd0e278ac5ace115318b34486d1938493036531fc2d90e6ca907d0f582ac32b0cf8807f498455dc30f432cab1de7d8fcda89aee3fa0ae605ac402d7ba87b334b0678aeeac0607c429c8a3ba9e393bf85d0929784291c3657a44f219a3e87b7547bbbcfff344e03bbacbc4a9d688432cfe4ef31ad89638a7df284d7609b7bee47eb8985ba653d8f91ae67b1364e980a3f377b08f214695c1c741eb474149a870ca012ba0d64aa21349a6b779bba647bcc814e580832179364e5cd09c3da78f654338326fa50a7c04dc42ae909ffd4e1ecab52c8e0050609458f8f78ca30d0a254229a965b8a7d2c9bed54af57d5ee35e786063d0bb4f9a6ac063ba42c011090cf8e9f0842981c0038a1d2a36c012736388e5964386f0f9ed2b5dfde89a267276635657fe646174ccb5efc28e0be42ba120524b7d919f624bda62bf4e4b153d9380c461b90e1b01e596b2fcd28fce07e7963cb6628118d77b4160dc6c71a0943529b9954c2cdc40f8ea0bd3876e4c6dfdcce6ecec9a0917452e9b37b207ba08e94b6ff185116d6c21818803d0257693fa2b2d780266186246fffc88b4de6f20ec289092085956eec1ce71812eb648734c101712b78558a004c4f2d5b85d72b5d2d8f293a70f74025f184bd4361dabd3a80b8c491d4edafc0566f9c0950fe42ee6c670a944526a4641b77d8cd182941a9eec34eb5d0f7cb73222c3ba5df272df6e9131b4ee90f180cb6033f6d040e08709a5c004b0f00ddb204cd5d75f94bdd2e80c7b29c49d7d5dc076db94ad8381f06516280afcd3601b8de8cd81e2228d93631d736be5e2a037438bf13890699de6783f32b728b8b46917440775c8833208dcb3de466457677093735ed56dee13a1d8c9c04cb2de68ae9635d2211856cd313e7b5f19e0956a51aa58cb4fd66002dbe41c0f6cbcf28d466a3de5980f5eb7c994b193b8c6778322248a17ad4553ab050667a17bd53c6b6f21821ce2f2be824a46f679f14766657a582ede8cccf73da1c62635c7acc3bf592092195045aac7f4cdf825da4de74ce22bda567f47a196b9a0cff55bbf7d9ae9cc5efdd668437188f763dedc3ba22c4c274c5c5ec369d60d1ebf14cfdd02ca752eb9daa09c666206760349b78c4ebde70e44f1a6503a5620eaecf184652330ed467314df40350e8d4419e1c878a73ceafdb3d752fdf12d15f50bab958f4b0a926da11b653d84b45113e2bb3afb6f686757cc807a36dc6d77caed81ce94ce9e310e4a8ae0103c95e6c1e27f656cec413baa48fd580298bc26e600d28d37104f5783fcc6ec528199859bb570b7b0189e4d35347bcb6d617c0fef514d3bb5ba2b5d496ddfee401adb337bd03b23396f7e491952741455a7accdc9dd39e8cd3208a3e89c926d3321c5c254130fe60ecf362a585953ad462dd8f822504023f037e82d66dfc4c75ba6c4a6ee90e976c4ab048817838f736b9890561e51ecc4a3fbe626af7234a7b01d64af35795d5cdb9c4fb0331da7c5de54f8cfbb3ebc32b0845d43f9d92b73d01ecf4790eac2e064ea23e751bf47f833856a2aa7866d63a8ed2ca947cbdac725e46dd2c25b65d1bc1b69a85d4bf0a87a20d899c7d6defe7b5fa2d52c93486123a6d633657279daa294b13d0672eab4d34db6d7e2c9221e636785b98a7049c34cbad88c67ad3a0d55262e225c1a7b0c3f4091e8823ca3fbf19c3a19b3a687dfbfedb978829ee74c4b92a7d67dce710e98e073791dc1959cf6a8eab2eac1b2418e5c3bc1b1fdb9409e230b888cc3d2a9a7dd71fc9215171e134859a11dd13a599a71952c2b6b504c468d9571036c62ae2dc21c6f5875082dab774f5012acbb23fa7830a054bf391b69871b0af10500188e1ac194719cb48d5dd0ca36191241dccfd81c83aa3283115c315ca8262eea5dc4bed2c64d1dd97004a9ec065d73a512fc3d43a8f64bc57d95f57648a03d73870d247ffb80eaaf56e90294b2cc96dd908ccfa741e61c74d1d71d5e328d7aaeba4b7b69af95759ebeff72693a1f0e8b45539aba60af26f115b1a64fb31fdc570916bb619fb2a734f5be498cafd4cb506dd431dfa5eb2d1fe6504cd50118aa64322c39daaf150fa870e0d33a4afaf97e1530b1a30e88003cb7054c27665e2c0064bbae1fb2ca81e44aeac9c3458a789f374dca405c6ea9f5ac6f4dea4943f71669c00487521365457dfe25eab105b064e9ae107bed692abc2c4812abcece822ebf738f115c8ad4658d46494b55eec801cd139b942254da0357acd9342645a5ad99a038a04b3507dd0b530bb9e21689e2acf3badb0added8770a8403b4c9c66e3653fa3ad7a1031f62151cc100149c599fe332a4b5299c8f07a8eac145703b31d7f4750abfc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h26fa71ca35e24e9469f3327e28c5564d849978d0d290656df0a0ec2eba0a6dd7582cbe4856637efb845e55b858b5ff417c131655b30cd37c2a1f06312e73c34265e14ca15eb3c48b07665a2d373a2c839945c91ade992b49d30cf7d43ef55ff4b1c32b7cbf2e4cf1be32257ec99c29b17c474c4e933dfa7e0d52449d4e8ccdcc6d35f0f9117ae046f3cfa7a674c2c786d0e10bde67e4b869640951953a95494b2ea014297c56741722faaf42d9baa447d40584749f66545921a53e8fb0a07bf293ea78a6078504c75428a280c5955fa50d43aa2f30fd14c6e8b8eb0f9c7c4f51df54f22b7e9948f57c36690d0a7d53c1423f1bb2971d26ffe678e299f3c7a3a4973f7d4c9f9421ea41dc2eae64263bb55d6d06b31473934cb4fb286f44c7a4ad7fba9eb8fd0f6eb6974276651630906ca8d0464a5e92a7d66df72dd22a027bfd69edafc20f18de1907fc3cbe5413cf8b311e3bc75fd1b6294a12a4e3231c80d150feec3c17c12d04c0b714f6c1c54ab9f6ac1784bfa9de2e0aee9692ad974e263e517011140166578ccd58eb0764107d99864bb21025d2c6928343fed1bf763818e0ed95e68c017003e174e4b61d6b78a22561ce33c3db8b23ee44ff9d9c8fa6f1c20e6a7b91943cba93a741a19f23b70f4432814ba6b6c1997d291a6f6c7cc16d333adebe74fcc12f92e6f19770a707ca26c6e593d2ae2bd842850b88da4537263e82014ac23ca5bf119d04b3a1e49f3f40ff83b689503df4d50b01d75708d933ab4cb555350c2600068c6fed071181603dd268d9e226d7c24803add5e60547ad3c4094c7929328afde6fe39efbe2aebae601edb30cf79323fce6b18b885e0ffd9a05b109575ab377278677fb80f5b99caca88b48512ed754eed3a65a3bb3bfa20f28403878382688a88c2c759f5bef6547f6ce926fd6efd38b62ad3c359ce9d7e9f6f6ee7ab74c928325c68b4b109ec70013c0518d12452652e420800e10de203ef5e7a24323d9ceea32001ed64fd222c7f76ac2c44aac6abae99ad67aeba3cf6a6d766b260b66cff2ee455094c5dbc95818b42e910637e83a3c6a5e7444a5abedca9640fe1aabb955ed921d44dd89c2a984c2957b6927b2451c58284382c40a98553dfac1fd3269da578efc995712498e6e09d6ae71ac477a283d7f9ec6988dd45e852f31e9813cf2623c1649af4763e4a51895a7a6d61470a08f1c4c3c4034c4d121389595e4a8d1b18737291ffa75f03bf366477438d54111fe2143ee691930cc244d3a19909263a1f5ffc6cefc326dc959188facd85c414942bae90df316e7b933f0e771a4cefe885bd45a9a5b5f9301f433d18d1efe3bc0387f41cf8a5fc778670fcc7d132898a8c8ee026ef81a021dec95f5c4f0ce59c5858f03a7c38d900bb8c4d4839cb1086885042850ef981a603da2ce621ba4ce52660da0eaa3136bd3779a2f829d073ca03709e8883d166cecf82bf16de82da5e31215d7088fb75d8bf1c15675fe1382ac44190d96e6ad37cd5b0a36d554a05710308faf9a8fe6bd9cc06aac53d2d398b281269c20fb8ed1ccf3be2d84ceb120a417c04e7264d899c5cef15836b553f4d294e00badeb96ddd23ba1778e58c6bc155fc49faa2c7bcc65b26f63e6b115a63cccdd0ad0627e13607cffa1146ec8ca6e53d0ddfdd7acf23ca1ac18aca535f1bcda41747edc33818d824c43cd009e4f50c546749ab0ca5be80d726a1b3b079c2b2ad3d6a56adba16a376472c7490ba22b04a4d0ea39d7825baf82fa2966967b89409bb4a744abd8be6f2b03f6e2319f54c8973d24af07ece7a049c52c8cd99d9cbb8a7318622c93450bf19456d1e878960d3df1ebd1975de4178ef3be7ae5ac0afd879b0798673f23b3c64c43e048b97ccf17ab401f9b67a00b8837f4f8809b9be0da7b9e22cc2b01a8fe56471bb1fa16b12c364e1a8db778cb4ea396af117f273938fc29aa429d3fba00bd041c60042a3629530716805494b8a7b201b7746f92bff73e92ffc30c6ba9dca96c59b726429b8035c92cb42af826b88809e54c57627c132fe288d9af5b007873ac02df4f12835e14d15b7db7784ff765d0942cde718cde7989ee47776a50bf709c9a5e85221cc3ac17b7badb67e9c7cdb1d2181b5f379629e941604b1f72d8e900ab04bafab23aaea2d3b4b821a289439dec5b9fab0a282ba29b599609fbfff26aadbb4796412080df05b5178c05ec4e27a3f841b16acc7ebc330c81035ce3f48be2dc1e799411029546754266d730b2942d7ac94c941a65a42886b2ff7d4edeb952dc1197efecb4d027469fcd606be864b8c17d8f26a753c9341fbaec32568ef74d61cfcddb35edca4c590fee91d883fecbd587c4927a8809d6ae61f08644af3af850452db9558cb1de8d4cddfe1a2e95ead6878aab3372f262cdd85f3c2938cd6917f0fb2f632b059f03421f480734a1b61345e13eef203f9fd585bf32b5f477c6a108efe3720956b7524bf72bf2c34c7da9afcd67eabc5c199c9043738db0442e38e125002129834f4125088d52f215f300b119dffdbff2bd67d7e77dc427865d33f55ea77ef1e7e2a36ca62c7c3d2bbb6b5f67e2a9d3d70e1165905b03fe898405d13ba65654e46db55622b7e892b7ffb687e47d53926c3406d5c520302fef939b3332b634a40a86aba3663b25c60ef872651f02be94db5754dc8e554d48bb615517abb374ad3c796fcbf4e42490b73fb18a498eca8d38087f477375e1baddfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he187e3a974ea42943fc2484f724b06605daa4a9e80ed63e8cc38143716f1867a5f8dab207ea770c1491eb46613a6f1231e5dd9a336834b790ed381f1e5ecbbf30fd3a7ef75a3dc58a9c765bfc7ab433f4c1d82f39831e3a926a24da9ed704c31eaf1144665d506af4b32f87832778402e4831fc64fc0bc221da01c957903c8de4b31198e81984566b65d98acc168d9e875b25067d582fd11ba5cc59fcc52d796d0582b99137bbfae7044bc0e72979fe5ab7960b8161c44261564c1c20c787e8e54117329a811ea91409b2383a9c7d242a54006606644d06d63ef40ecd19c93a8fe5052ec095169bebd7b552e9cc7aa82029a8fcd74faf822fb8106f3ca18c097c6c53c3eeb9fa785d7fe19e49b2833916dbb8e8f8f5a77278c3f56b39a19c95490430f42d575c328c4e2c58aa737a6a95540a9177b536511474eeb263e532840fdb971dcfef5653a09b93a0abf13e5a0c28231c13d56994eee679d023c0b5a4b1e9a715f86a6b2b44b9840d55d28262ede274ab9c1ee96adb02817c6232d47fd4f6aa3b4c1ab2609184297ce53718df791e2e7146313fc51d71aec608fcef5314796bde00a4d5046b9ecd4195eecc352c76db3e8fa33626682309d9de5d9126a00452f3b487112571aaca14a4e2a533d1617ea6c55335abdc13cac06e6b411a0e18a0e76e36ca0005ac71c3a121e44435480911df418b871e16f3e49f32657437c5fe8ef1589b5a6e41006e5d2379e65eb5d313803ed832ac8ac5894bad70cfcd207242f5f5127fba43ffe3909b883d165d6933619cdfb246cb68016ab3d2054feeed2eca35d828a3fb8002e0564c5682f4e855593c0f2f230388416b32a8176c67756a24e18ca8ff588b99e20bebda6dd80b4c1617a5eb588cdbcc31ab874df3d6ee078a7e9a9c6b5514eb83fb56ad89a2583547cf6ae8a206e0dce58662fcf21aaf503e3c7644997e022413a7573f33a3064b6bf0ceba4d8255f8ef19faea870e54268fd3e74ed67a9be644ebae6bdbcbe31d68511e93659a950c494659a6ce81be4a0957efb1a987125b21c7cacc0ef5758e3c996d7711ed4b2059c971931e014add4eba86f886600d5521183cf7830e959b7675dbca9529589c067734de96fbfcff31be8117ddb01e23690c7babaad990e6cf1063d9ed1ab24d53a6ec147ac7ce51affd997cb07f225239bdd8ac0800296d80d917da53ed75425c32a8bca4d2e8c8085201784f06177b0f43a57e8383652df59de234197d6235dd9849dc5b81d9e5c60655f4e77ded991750915409e2ace50302c092e55105867ccb1226efec866e136d554b6b65215cfd55f82589642bbe3b6632aaee11092bc0f96c7c2df8561d61af152e52664584c584f2c2a887988fd087dbcb5a1f53aa5848c64f41a30aad991caf7eb3f058f8abf11c2d6cfc04ef173be94cd998409c87502b1d156ada4a95a280fc14a96e82917a37ade87a68de7503e07f0192ea07412f7ef19ab4a530f71911a0528eddfbd8d5d40b1ebba37f7a054b3afed9093a7d2a1fb8ab0e6accd25bd3b151172bc70e0942b6c834557c07cdf4e417b52d2c1c72714335732b701e8371c0d5617027689353be76692123f99d70fdbdcaddd9643eb8f90f3844653609e21d2d84e50863e374c9f29ff2528d1503fb8a022d780c605ea5b15f44a54338432af7c69fa8d0a7902e53acc6be67edbefa8e4a008d2d065dfb18c608176cb71b8f3077b9657bd68e4983bd3282d82a00c005c7e0abcb21ec724232a7183d42c783b34a7641b56643ba55ca6f831dde45022543074000e87facdb11a46c3709270a405f81228a8eb66ef900aba37845dfff5683eb203389513317ee879af761bed26cf6ccfaad24395fb82962607996d124b6c9ac5dfd87ecb9c93f68705649de0600be4c3ac2b201f90920d1cdfdfb660ad214211a517472fce0427cfefcd3817ad14337af2ce6c0b2cb1e9c1b458d7839a02cf43ef10a7223136547ff315e3dc8bb6aa44160480ec2b399e6027d39ff9a13f6694faf4b0e81be4218878435af5ad97479e41ddeb7ac9cd756efdf9f9f489bfe88792acd1b36544311a1e839fca05bd9d62be26874aee17dc84aa0b60f70f0bd2d97c407aa9d98f149aead7b95181d5210a90831a251d5a0b87c60a15c1fbc23675b8eeeb3ad31723cb6b2d7c50d1a046ca87e0a66f7b763fcde8995413c449642183708e038330e49d0112f25e5faeeca394bc3156b5e0af6fedf63e354f35c6fb729248e11e405493f84cd9483a25e72b7e1e8d76bccce07c9c7596b1cad974c2d46b2aea43ee8b96252a91fa782b56f598b315bb2097fdf6a6b486700cec96d64e1daa3739b8f9d2772eba2362601f25339e531bad07976454d0da3f7b14c4edd300f9697974546cd30ea23c49af3a1889136365c2e0b5e47c8dfefc3cd31f4a6abe79fad0776595e1ec3128ee8e914aabcbbefeef19904751d9a36792bf518e4f80099e9f21fd3e45716daace1940d2bf4abf7e1399cb930215b5eb228a51c088b5f8fa226aedb79f256c110e8acd2cce2476859790ffe53ce0558ccb119b3878d57aaec7cc8d4fc1677285d461b8248fb5b05107cf21208febeaab81484edc8740e23dc8d760e3439de2e3a113aaf374e4f616453f1cc91362013dea18e86635a7508c7abfef61d1148f8e3ed2dcecf4d117ee48693e5392cebbac5fa39f9a3e1a76adc66e8d8837843ff210786158a69f2ee8d4a2d8f67a1d0c3d9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h902546d622c96edca09dea2976b0ff07d2c1690d7b0d0b8cf0eea5be8a9dfbdca7c7f57aae7aee900e1906b86f2dfc1ec6d93aa6f16f5b0e66e9db2c5f56b4ff171e28a0a2d5cca3263909a0eb56d5e8e76b5ef4a68eb8263d6921e03b0befb61baaff730c3dd7ff2cd11608b1c0e1891b25dd63f0696c001447563b7ace41810db3dd0359a3980edf8878a0bf4a0be2079f274a7d200f9562e7e08760ddcc90d6acf46b34d0a70add8b2d5294b2d7c1a04bb18afc1ac83cfe21aaf8ca5944bdf992ad3d9706bae63d3e048afd265b672e0dbf8d7df58012523efc51f4dcf0bf2004b8e577e889185ac5c7ddf7e877dda4282a39f5f731643ebcb35e82212e0ece86e7cfc1a203957b693af02360d9016dcbf8fdf6660e53a584ac5480e32e4c6954168e2358a06571de3535196bded824fb4e36a0264ffab016c9dfde2a7c1f360f26c867d78fa9174fbe569c2b959a87582dbc3f312585c59804ef775e8b59b358e805909c6ae18fe0e3235193225f3f8c7faec0844940195833e9ccd70b419bc38aa25b8b24d6a6f4164babc97f3c785da64d85c7360b12283a5758e2c297fcebf8f44cd00269d8a026058ff22519b22a840c5179583218bed24ec212e8502ef45fb253427818da37a5aadff9e2c387ee3700777ed7c16ea399ffae71e3d1acfa3e8b78361ce56bac102db0a945099df20deb52634c37adb44e0e4047b9f46ab9eef2b211b8bafb945aeb88798dbd78b504b821724de8f59311591747c23d2da7a4ae3487d4717da8b1d50fd2e5d8957b092b9602a0e914fb1420c9ad7ea8182a009ea6739f36f1c93dcb29c8e722388c0444672ae6919d0ac17293df257c5b4e8a1bec558adbe3d65c3964b6e631dbe50e2822439390e4c71638d814fd9b7b05cdad6348996932b8317033cd77de5e330bb0aa932f15f19cd9b4d4f1af4bdb7a535e4e177d30a738c5c9c09a7e64085b339ec6d5e14ca5e639342f59b890dc7ff219f2c39023a7bf44bc5a4a32622df41d034af6d0f1cbb3b7f78d4789758c3829d781063a64efc1d90e0da5fc6159590a2f6cdfd8116009597fad384f30f54bdea0bdecaad8e867f96171d42a6e93e66b50dab5410e150b66baa85b4a9abb76f14d694c2760b07193905e4dc5620f7026fbbf18e4b04ce149eb31922e88616e3dde3d3edfb916b1ffa0a4e6f8ce311ccaf4e229c49f9569b76695414078b29bcf719952d77f882dad2640dab5405870f6b9ef7cc6f9ca901903221e2743ab662e266b61026f6a61d8e20df49512e1e74acb9bae0da8d9ffcb926f8ee0104e01dc1b170e09a85c830e0ffb11b6772fc7335b235f508339237b7316f625f2c4c69abbffa63ae5249477117dc0b5aea29c688fbcbb20ddde238790a289c5985c61cb737af9349f8b1e0c6e47e6625e773f194371ed597550cd82fd746376caf0d445a98d5b6715278fceec03110e2ec051803acad7aad4601a6ecaf0881dfe270ff8e6586c92f047b02cd91332f4cb7a2cd30cbf3dc6255b2e09775455279887d8bba3148aacaeaeaab539fbd9810a8086caa9c5c01f5c9b18df33fe792f42ac475171480a0121ff7808fb7dfc3620ff8747149d66060dd356595802375fe7b8ac77bbc98b165bcf594bda1127c9267a57c5dbba525921e0a35b38a8f610631c341cc78fcecdfcd144c2ff6ff1f9aa27754bf7e077abab707727f1f698b5a0abadb3cefb6299a83b732fc27e0cd324a18eb1ded0265b0375cf7ad6b693e17c595ae5a44a675060a21616e883bae8013538f55530594f8a41210ee3a4cffcc003c9cbdd6e7537f9cd2caa93d5b90223f825f8ae78ad1bdf2dc01d29c779bfe80e8a590f22dd83b358535cd06a73a70a945d1d39c3a7ac26d1a84af3f1d8cae2f1503d3253432c58895767f70987410f771661666656fe4a24172462e5d3dff3394aa948d6345e7a2fce03b0789f91c6a42318e2330c7ae278f41f3fcf0ffdefd37533440245fd5090e5333d9be8a0138dace3279d496bebb289b2dda97438c72a6bbe4e2f2a5349e9672e9d05449836a1fb2be9b298d9a965c46d29cf437589ebeb106003650d9a456020c03dd995225eb6b114d39c442432e260f794e37804d40ca1306c51474b68d41233a40875fabc60b61f4517fa1cfcca3a0fcc67ca3eb7194a4d3d183467c30c5e66f70ec397a3f00860db68248037c1370bb6642c84e42696fa17d2cb246f0c3a83165d4119bddaa4fe485c566e5cadaa0fc5d6bc66b7bf7c9d3d411a1b577565120a792a1da889eecec9bed1f4d52f009e88eb75562d6182982985b8d3afc4c92a465f8f80eb7477d7b291580c120e009fe7926ea77327b65fa7a6d85922c3f3902807161a4e460dd4443ec99c53d73cce12468538e5ef740ed6d812189d7eabf0523a7c14050a5979b7e8f7e55fb3c2b1f7fd8201a8406b8a4a4f1b4eab14dd0d90f07c0c0b6689e17fa0fad9ffba72b1e1e4acc3bbe28c1e045a027b30681a7d8ab60e80b42c36f7f92b95f0bfa2b20cd42750938618aebb5c191f22b29492c5f667d38c981d82454a86d1138b3ae79cac1301626014ee6b8adba66ab25da427165257ed3f1ca733d6908f160cb37af48626380aebc5b50cc2762165136524e8effe284ed0b1ac377224f174c42bc9d552a11c17f16dcccac58e2637b2bbe61653c963eb2de7d21a4a1dc5eee1c1b345eb41873c2fbacd9f4f78a43f3b8f802137617a5598525f18e6710fe7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h38b7f36f8c0c4079f79025024bfacd44e4722b4472775b61d30233d4a9c3550ba7f7210e84c5632385e16231f85fd3fd71fdeacc87c38e8d8083ffd372a0709eabbe7ba71f5c7727db15560848756977e69a0d6b7cac7f959df4abf6cdf4a320845c91bbba4deed71e602158dbdcb921223de346ad9ddaca47c10e3befcb70f0b033ee627ce7272bf49f3c2fa0e56b5d7479f32ef39eefca9a9dc27bd5ee9c577468a2140a405885d4d5ace5b7e8e7fbf8997feb9132ba9ac48563dc506a1111afcaa00b795f8d05895cff3faec35bf42edf2ec8f68337f84b551afc6b23d30fbfdf92814a2bef09e77522b761172318b2530f12e6d32e381d1d96f1379f08ead8dca02a99e5e6baad76d27da6fe57b56d047c90f0f1a42992be726e36afedcb962138e23c8936ab7a70d33ca0f3236a721b7abd9bc13729454744231a52da3aa7691f98143622908e7213899396642695f16ccb0e9880c1a46e271bd8142900a14e66ba3e5e10fa7d5c02c5263ba19f68428d547b84d29f26687e295ff1b7b2a0c363c0ef3fa66c6d7e6d9bd604a97b47b2def656f3f4b031ff9673e61455105ff77199c5be9881cb00b82fe6df6569ab30ff64b5deba615d54aa5286c4ceee74308d90baf1584bc285c23ed945198c12dffc9cafd7e8bf4ebdb7f2a23870ce83ee4f86db525df9e8c914f572d23dd83fd5360814af4458734cf8d2a99a4d27e6ab4f2f1005f8844914431a4112287e366203183b8309624241dfde31ec532fa026c817c1262fe18f3eb064e6c2a2afa9de98372c636196c3ea12c42b2f75c34501ef7e8fe045dc7c85a3836f39c55476e3e3a1359c40ee5e70f4437f3ff77fc0506dc501dbbd5b48425bafce82c1fa56bd41bd4814898c5f96a647b753caa53ce9a260fdfb5996448e37fb8ae31b88a1c48034abb7c5dc88ebbd75cd1ab614340c76ca10417d30029e9e928f677369ab7c53d7d725c6d6a576a2436a37713def038d85b4f6de30a82bb1e0b9f8ea396ad7fecc5867016677c604958d563cf69725250227dcc7e89fd73706795ab3341428009254cd18dd21e053fd8482517747cae497a45c64befa0df8468483b69ea51bbaf4a66e0f4bab43b12c272ac894c0ebef09ff24825bbdef14581a6419e2b4bcdfa9987d6c94dea0ffd5bcb2671c6de7bb24e464f82e49f586ed9d459f71b6b61a4a322e036304065a0e000416b702bbcf60c0ac7062770da1ac694c7b1c0b4170dbfcbc75d26f8ff872381141002262a2e641c07379fb355ff3a83bffe159b683353c5a1e7d6286be44aa7a131a1bc78efe08a2c6c15b05ca6f5f54c79ff28db933be8cf1444ff85a043b73a0f0f35ccab224fb8b0fb402c4b3ef90db15b27905b3d6b6dd0e1752dbc80de882df9b14566f3fdafc8d850918efbcf375df83c5f12c343831616ff7d0857975a0cccc31b2cbdf851d794f1e91ecd192800dfb23179549c3995b12348c646ca482138499637822405bdbdb68d599a5042d8a2ee85776b51425fbeac9ede16ba8c1a136ec5395ceada88ba5ab73d34c708548f5b0c70040d73c9cffaf80247f1ca06d60bf9b620d62d49cf5473b13c36ef03be4abdf180ac9e89aff7e81743aabb818bdae615cc8702a4e218bfc3575f760ed53690c077a54607591881f20353aeab4e9a26a4558280b480cec71c79174bc8c5d1a7c7e4a4907979e25770ffc03c3af71d080794b09b67a3a8fb8caded52c1bd39c612e969f0b202483289886e0f4582b5c7544aaa3ac1767d9967b40faddd05a775b084c8638c2e7439605b96c5897fd689be6e0416e6c6bbe9ad9a87f4180c0951785119e326705c801f7f650b8181031d0d557751030c0f15b6558caef29c6ad8e1961659f0f224f9bd317dc84a374a075e442b0893a4ca769c220dfc9adf8695c4eccf09941bcf8ff50200a5738b5b7047761c8e18b0ab66d7b4ac1afc67ed66fd102624b1fc55fa29973402dcd9900dfba6d69ff38d66b10ce69c28c7e560d561319b6880e870e16cd4ffe0c6cc6dbeef5ce5f3c93f2a8de2278e2c73a803b984d79117d1f5cd46a7e82ffefce7f1d914530b7e583ad4201929a934a2826c997d502256c770becb5fdd54ebbda153bb05f70e16fb300db3cdddd156458936568dbc9e32d90b6f0f090b69cef25d4608a28d4158a5c03235af3dc24132307d8ae2e050ce55b96efeb145438992ca2973e83dbec78dbbf38ec842c55f0a90c0d4cc50d6f5b26752494070ef4c2a6d1549dbeac0c468f3dd7ca993602c0ad59629e864bb83d9791cd05b1dbe7dae21d6edf946da6d5a65f21d4c5eda1ea610bbc4c8b1451785e8362fcc7e19b733dfd0e1abfade4371faaacafbda1d78dc8406a66e1e00b9b31de88b347f7c00c80b685e41a12aca9ccac79e823471d1cd9201308339ee17e112db16a7b7ab265d37849f1e05d5e39a1ed436ffea5d32b8dcbe3a197d08b5986404451981563ce1cfca3fdd44925a9cfa9a8e1d60294d16fe3fc6ed466a67302d0031739b91478fa35a89ec921333c541d7a0ae393aa11df21ec6323ac3cf20acd74250751961c7cb0804ba63daa738276142136dbc9fb85db5457780b3f2fcaa48fbf4859d7df227ec004592d29b533f6c04dfa7c5f60db38795ee73f9dbaa6963fb5eac7abc49978b234ab322d90d3e812ac53a4e9ccadc09a266986de6934237c2ac88a4a97d8e47f763d743e27e13e33ba62529a83e6e8a7f0fdaf58cd78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h717616353eb076b8061c8dc9bc21b81e84e9a00282985f4b1d8848fe701b227d39ba600e7d975944dff508ca9d947fddf1537fc1702cd93501e0fd92621ed8794f1d319b7060f541f488c967e2dd20c83097dc1f1b96c0f48cd576a48c31e01ef9a805d0969786afc248e3daa93ce5a4147dfb7198b0298af9e09c45e616892ef3798ccfe4c67a7521c140f8bc06120cc775583eb902b3c92eda2e443aa1ac3e60c270a026b760b12d32a8a79ec65933dd7848492d3f6fe03ac871421ff09b72c632f29270355ced143b705ed94deb0b1200f54ccfe17d454ef67e5e99e9f0b2f9fa43787a31a7b3eadd948906904e4ef15ba4324949924d72a25fcf0674735d21e49bf107fd968285492ed479207d7062e5d151b1cc6d12987dcbc22c9e807165990ffe66066b5938d5761a98acc2a438b0381a45b727beb92ce39a24099f44cd16c356c631a6276985a665daa657eb04ed79417b7c31ac6246655fa554f71e1551ae2b9d4c68a33dcec0f9ce67dfaff447ddc502d23ad892dac49c7f0c8fb207d95125fe220fb77352cc359f9c141374c91218ab8e3c4dfb2dc922d3a9a389d5f70feeb3a97ab229f5c64515b8f6ab1ebf79eb5784e026a22fe9cee2f06963f91e2f737cec6d8d07000c2614129177c981a1a10e10f69c12236a536dbc5616ae4a1e67bfd65f964eb8ef62e4fd536ae78688a9bfb470c25bc56ef6feef825eec873bdfa06c5c809964839d970aa77f363e842cc37de4c10b380e682139499864c61b1951bed0ec3f91f5a4fba07a1e7849478553e4ef1b140030a3d94f065ea2c40f68c2a18cc12f39e1535990a50cb130d9598605e6c124a7696196977a78abc0b725376c73246fb1c7cc74222bc42a7eab3acdf6db39e1ae588a6127cf55470546d7f409dc524d7a0f11fb739cc4fab8b60426ce41311d1c595120fb3dbcc47f2cd198a207becc95d7fe27aa961724540a2c354d52d4a5f98a47cbd5cfeb46c3a8d15a2c5e942cde36c071a4fd5a0ce1190439aef76f967c37203ba0e87f242e4121a0dd4debfba91ad8ab6050d3c0dd49c732a8944b8b3ee995879cc48c68b4ff9c43850076653a6e24435d03546ba8a227d3e7265a4bd76434814bca3e500a228115e66a3ef74a0caa5814c1588b34511f5d2c8c9f7482c8de4177af0a040418f8091682efba2fd02a99c6d2db2502d0630bf8816c9df489e5fe4bc62b3bf0b22b9b97128e3e3ac4518a48b381435f6dcff57a40df3829527c6ba4506ed0756000b3150a44a29f2318833b7f701ed8d6958495423339ccf66c252d1f4737f5c8641b69f763fe263d8234a71ee1ffa52b140a2d11851bfdd27bad38c360256075ed1c2d4ad4819b2ccf2382342b625edca377933f0c2a7075a15a4ea0c47dd22d4ad635bb618a0e5d2d86977902bbe3d0bc04b7c64bde7ae0838ce6420c262f7dc7a3f9b039e7d7ac00d36d8150b458cfab5d184cf961a412e6c632fccc00330945a6a890e81bd057de47c8950761fe97515301acbb92e324dcc4896aa04b80cf45011cea533500604f7a83276c51bc657384b89b52359f4f146458e46d6b613c4d4713347d3a52430bd38a383f623498c4c1a80b04f99253c23c07a1c54613115ec97b49402c9f8113cf6947cbb23937379107f102a34efbc06e8335d08df3d33e76bf7a0d2aa863214a50646e5d1558f188458996b8181a3d7b1c6434c2136ab0dfe470a5af3b8f9c53de6a43f0e5d67f5e92afcee478624b1fb4fb2d3e2e0af98b7dddbd62941e406f015b23d2acc7e3176a968a938e5edc7dab33bf36f2e29b5ef5f5a13fbe393122f76a5ce6ecffd172c01d394d079d33851590df549c180beb8495aaf5d608396c2d44c12a67ca48f0ec6a13b006d2f97bbc302e1407e606ed1fd1bd9433da402e03e8d893ce3cf17f4927ed27355ecc00aece2207a0927256c3424e5c2505567b854275e57b16b68d0dcea275341aebc8ee2beaba674619ffa3dee2b7caa02cd1d502fd289aaf6931150a39d690d3464b06f80813093dabbe3c6ff4b22481e8883e75e430f2ca36387ff928ef387e6cdadacbb1cc6747985f9bb8e93d189ec17da23645fb3d8d2905db9b62f95c40fa892de272f224efaa945b87270617f88b8c16f0de7b7f3acf62e4e853796c027cddce23e12c632c9f10a0a4cc4346228068e7152fcac6406efbdcf1fd09de71caac0d0d1c7ed0441504b8b93f317c0e4cdaefe6c18d6d438e0deb3739bd21a82ffb4170ffec016d8970d04dfa1fb7c55ec8b4d5b264420e25501710a089c5a3e8c634f15c069665881b20c879f78867f4144dbe7fd920f2216d90d8ac7c6ead4f61d0992c77c87ed34385043c75a06d17a606ec42eebd3b85e505f2fdff4bd53fe0b49b2ff31cd03d17a5c3256bb2453353192dfdf771a58c92de5ea766ea7dd83111bf295e7848c45624a2d14ad2abf46640aff311b4b30fc4f7ab4a2b80a01121964b8eacdab3b0b906e955b7161645110e29aa15ccefb3ab46706a82b6e189bfd8d583de0b2d262cc59a10cfd08b3c9c4d34f93959d2aee73cf52540058ce2e66229e9536f97ff7196b6021ea6a3ee2057bdf281814e82056451c8ac606b261af1756c6b273e8aa38a152bd38e19b3fe3cc13bf274fab4beb20f538fe4c541ad71c6115c21469cf91661ba7f229facf86ee81ff7ec69176b61b9d0d6aec1de515d2ae96a37833324eb378c4bab7ae7b66ca75c4d636ae9604d0c57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6c4988a658f97526541b3172a706281b220b73e2566c4e02edc05cda35d68c05814aeb15da81eff4f0aeb03fcf83c424637af09225d41109af9d8f60149f8f9fce1c53e48f96b6cac22a92c6c6d26763868b3ee1ede87791f71592a082c77449e7e1b94b1b6a79209005b65f74430ca9ece8533366cec8aa9650a6c914cafffb52a065e3ce12ba11523cec0c4a025ae8da95ec299bd07a14521d1b1a1d5222e80cd348b7b860e13dee1559bddc74470c19781f24db5915d3f30b2d55ba38cc5ef9fe9177d11c484052652bcc7c590572e6048521cc9bffa743d071de11689f13b286f6df5a99fda0887730a21e7103e7b26c0a7b0d961197c856678571b818e81276e7a1e285771b824bd23d1c01b71b45cd048c8af5fbd140544b74af06e543ea8d947d235ce70ae5d8417f1138d1fb28072a68fba533e7ddc744b7fd128575a3ac0c927295a95f1270cdcb8f8f1364e78822cf9dd99e18293f8d262da83600c13ada94642b7aa3a88dfed92e6a73aa648cd339acda9da4d802d59b9e6888b5f799b25528c178148ac3fefe8f61c529c9d9430367248dfcf6d6e30b65af7305797aa463b6ed7610e12489e29e5298399616fd678ba02295483c1613753530475edfb6d14331938215739522dc3c1d0a6eef6e5caab0317825c9e4ebc70627ce5744b92f45394a1be4dddd719d5a54055b38463367e83691cd86b74c695663e57d79a247abb3a64915a86c6cad48a3e893a839475df474f88f512e6dc005a8c7fabf686c00cae1faa7f3d8b49b7ec739a321d37989217341e073c8ccf4ac89b3bdf7b89b96f28ebd7346ae4773a85362a242382e97e5e61294f3ff43c469e3d09bf10aac68d26afa70d02f71a24f42110c373e26ac393cd0a015fdb3504226181b7763befbbe5c0ebb51733dd621bc8b0fea6a2707bc78135a426199e093a83b6f1c91c4888953cdb389fb06ec7ca58ac3bae4f6b473c1728cd7c4b2c4cd860486a9996009e63a19eb7a61ee3d024fa87d7961bc7f0dac406e3b472a99da36e81a0b94e0c0937a81c4f094aa56faf4840d66e88078c9bd48fa4ae4389160a8a6e217b8972f2dffd3ec1cf38ded874ed4f47dd8797d638ecdc316a303caef5a5b408e4ab13b28acbafba70223a9577e280740e385c2075e87556c0c36c77b6047e560c33f52e282061a2e4a26ffc813b78bea5af78a9760d0bcbbb6d0453e38689f7ac4cdc404f9cffdb2e66ac4f3670c0f19a64d1977e9aaa37a293284ea3974838859a439da42ddeb89dd2ad928d59a8c2c6d7ba7fbf2441225b6477c798ec89cfdc97b7928694d619833428755dc0892e901ef12525c495201186299017ba51daf74acab608433b44496cdd5e2344209cdc3a58fe844cee64bbeea5bcba5a09fa5a64dc811751dadb0c82f358773826f27b143a15fb1acf802ad4d8ee12af08c48b9ad96351d7e1f020c1f8d4bbd79e07c3224663d8f6e5fe0088452478ff0a8d303a7dc60eb4c9e522110425b9efd00803f24ed0857eb4d6b6726ca4fbb4cff5d1ef1e77264dec5ed2e91a249cbbc350048e472e810c23dd372d1c532a877b7bd20fa659f2ff6f1da32e4119aff7430be560cd8f380be049dbc1d7cfbcade621feebd26fed5e17aea640ea3dc6bb0c3d241b3d4fb270d269d9d01938946a5e43f09b2c69cc834942c4b4c7a4f2136966d92e2e095b3d2d1df32408b48aad808c6258c3babe48bbc876ea894c7aecba79539fe27c2664749b03c260030f6d26dfb7da5018a9d8f3e792183260bf31b5dff77dac4f8441ff38b9db7bd5696712170a38fe542ae5f28781794b3e109832607001bbcb953969a40e43ed7f9446d549c510d47f1b91e97b4ec4dc9f411a91d53854876bdb20525822c3d54fa2ee306af9639168dd6dc98099bc2fd1f983cbb72b0d84e6c88fe7d488e5d2de609dbee8c48d65f9bf2f9be92bd9a58a6a9cde68f988a18a095ee5307c40f59d60ba728d01899defc6298df19917f707a80a63aa225424a8b65de6325f6def728d3fb2e9aa75120dbf13f6ddb0c6acded44048841a45bb4552a3a5126a71416f1c28d45eea84c32da6436b84e6be8568494435c223421a70f5689c8fbd3756ae573e74fcc03aea2611b4c70da837ff4e6913f77ae48d10293ffafedd726a2d5d0365337b018edc0179b6e665fb42e0ceacdb3672d97dabc861d98950ece88c1f69c844db0340b609cab8bd4571ff031806e71c1e3f4e7779ae14443bcf13ce0746ff1eb37f91c93df6b9869b59ff066ac4635ef776c208549e12a5908ec10107c4a3ae3845fbd7aae0d6a836865b7ff81bfd7777060440159ae870ad51e198d2b5af0ae276e5c46e9c85f8bfb76255636df56f10fadfef5888261dcaa0737aedfe3774cc6e714ff8ab3d914d75f2d7d2f86b53609f564b0f8999f92378e9b2dc8d885fb28ef4534c8ef01dcf1341bda89b8d7b0e57f5793a8a21d482b200821f26220284ab91f0f5eeda4fd5455234160bae1eccf454a21528a6b45b1c27a726df747e874d8cd14b06112c32a6c6ad3eebe84db54d51d66576a5b5b8459ec7a7b76c6ef8f3d19a7bd7532aeeb4c9300fa203af66ccf9176d341915ca64764a22784c967faea286e7c389463d6a21b3663687c88637d11343a2930510f851997af9dc1ff6d5b371f3988d5fdb1277414d8dc84a2c3fca22c18d918db888a4f0f7e9e9e3f6767b8a5f1c7aaa0119c496a5a6a5c210b17804f0baf57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6c05fb38592e741d06c6990182c31ce60bc84781002cc86d5157bd6ae924ab1d3e7079f1c734e2a0d2bd9b0ae6ce444d97fbaa7b469b2f57e0c084e1127213e09140ea021b8d86340bdd9bfda5f78243ccb8ad60e56752f583d600081f8eca5d1625b03c8d99421ea75e2b3a33e60774a2c2aebbbe13fba93c8e967142dc08fb7c4278bd90ed29270f6f376b3651d7a0143001174ef97f3bb8bf9b90c30fe790d36b0803717e137d778bba21e70565589dfa25a5dd7711dc4dc253775503f9d43aa3085026f332d7e8b4e38d78cb8b77ae0220b02a817725822632cb46cbc77a312b4fb878c11e153b718120a4e818ae0d6a904165956e44987f9c8041fccc014aea1da8b6984539f55b4c5faa5d05b5b911ceee5ffc0f6eda9da3a5a5300e917a070a139c988d423717caf1b662343070f679151c2d78d9e6f26d5734250d6d3b98515ec907132b7f00756492a7172de72c95119a15cbd7398f3158b8fca53a44a8e0290f5ccbccd1405cd87a9f5ed27acedbfdad5c90cc26008ccdeb8082ae63143073e64b12506adf67d238b9ab1788cefe12026dd733e6aa782bbcbfe202aded3a91bc409c587dd20eaf2e7c0c564464bb13c6beb193b1698279c49d7e11e6cba424f299f70d88f6cf7d57ef1288c6b17289d83ea19b79bdb383a35bf1f6984ffd8d0c1fb2a51110c46ef5fbf55d97bce0b01981f09c027b5fcd1534cf387740e1917f96e367770633784cf3ef4e815e2dd979c1b7d353808dc27990b5aa3522dd5dff82f58ba29e76f10823b62f26415aac5fa8ec42927a149171ed556c18873fa73e421fd4f71fc16ef42e733e1d76ad5cddec63a633c72e37c0bcdf77844dc22ed45d69bd85eac72c35d4ad2ab79c8cd90ccda90349b148580980b9d1ded8dc628819b888eddd46a4b362a5dcfb13bd8c16a847588595cb544d1ad842b357d156a03475495de2a2399eec91414b20f0e8323e99fe54eca744902dedbd90e2306fbcfa8a2c708440ba85f0344dd5f7d2ebedbc34c5b5ee75a98d76e10ed0000e767dbc61bc3644e65ea4cf28b57f896d8a7893364cfa243c2d130179871c5016b5a75a31c2ec4293523c0e5cac9b73025fbddf717d5eff21b4ae8a6df9cbfd9cb7815fd46cdb76bd2efc9e599f91db60b65356a82331781f42615c67bf61503751942a6c9c0eb0df49e795b8655c67312507396def7f5edfeeb72ee172cd3247e8505d7df0a824a04a227a3aa07c0b034e9078a7fecdfc21543d57bcfcd8b6c27740afea5d187785d2a88eaaead58acc9826d0c18a067f3b16e5bf32c8247e05fb5f34457a3beda20aa63f1a5dedf2e2202330760e193ee1668f4de164dfc01c0de5dee437ed62f43fee20779b6b18f2a36764ee3c897f66112002491318f658426c18040a282d0d1b43c63d06e778385b0167e7edf699bd3b9383731b386f374b4dfa7ebf29a86f3c772de8b2c44aa2b816e7b09ea20d948e9136776a8d27ff6ef6743c7ea4cb3f62a5670faf5550b23bfe1b025575948b77f2530d513e74d718248a06a20d80bb1a070ac56ae6e2059fc146273960b1c92c52b467d190f99d7b2e1563fd2a507ca053edc74bc11e368f72c04f68e1bc142d80046e4597b4769f1e009f8669f207f742773e54cee2feaee3c3ce21f340bd355d2904f49eed0dccffe0575cf2a76ea3fe64f6e939ab29610b3e7651d3e6f8f44add96bb7ef3c880fd71935108b8b0ecbc564fbd0dba1cf3a76c6e1c9cbdb38e498b25b3cdf2529efb68401115ec7cbd87f295b5b1399f88b943970b915aa3a28c4628c30c0339114748c46401de783abba9de08d78766079bc87fb1ab15e87903d47107d15e8d99e44cd5e0f5845155f8c30b26c232baaf795017e350c184e225d06278a179b3ed9cc51a549935756eb7c5c765562878be0f49e9d7380b403170a9e1ed8416ee4dedc48c6d85e7de2fb08046f3395e61f211f74a55397be0e50f534ed26b3bff9fa2f820f2eba853e0a7dfb641cf045a62b64120a4d53c83f124bb1904e6da308c6eadca300eecb28edb2a9cd9965a9c53d23a10101a97a97371b2b110d1fb6148ff5c4f005e3959d75d73a4527269184862fffc0c1880143684c90b16a9bd887ef58b8a05b5ad1afaab9a88a57fbd062b20c03626008492c4772c751ee4ec512b1178d4e94235f73bcef765a4c9780b93b15080123e8baea9cff3d40c0fc50ca47b80371e7574a07a76bad181ef9b6f6d75eaf63ec2a88aa1268e9ccbdfab8a06f345b5e12779bdd77f663c12ca44df609fd867b7167409c1e5789532d250bffb789040904f53021f3a767f96b83aeb0965d1debd6603f8b064559d50234f266172dceadee95079a1c39b135848de2e08ca8ebb9ba76c752dd73dea43d074eb6c7b1a581dc6dec84aa66e6aa47dcee906e72100c07600c7185878b56eab92e8aaef0f9e95e47baebb146ef86d2a0e35ad65eefd146e19f49b62222787518b26501f5d6570e32ee4f30f0a8f9e38d8a5a56aafc527d5ea732f20024b3d65051eb637ba71c094e468db4933ceeb5f25aa8367a2c25ec68027681814edc05cba272b110f159f43c37b33cf91218e7df5553f11c3fa2bddaaa0f94004eb5351b89f82070ac33b1f1b5d6162d0afafa839d18d486dd9a7fef1e9518bc6d633760059773920b59b4565b47014a0695e9d3eb76ff6dd96e270e54eaa1e53b0cbf452c8a7baee078e58781dc3573c66856c84ffbd823ef508;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hcd0058eec48826432c064d1d9680cbc666761dbd284e297f0f26fccc7fee49bf3e427cfee7c2f77979a3dd45cb696a8d3d9a889337bd9d127b107e0a21eba7b9ae455c08c73b33a3369289962aa96b0e3c7f4aa25d0ab026b3cfcfd52dd53eb644f5f472d5fb36f70b6171c235150a918e4168b1329b9a8da49cc939cc1853b81750a0667f902bbb24166d7e8a274564be49f65ba6706cab8fe4448a922d6fb2390926027c30f29fbd0abbe06d5722ac429314541ccc4d7270b3d0a7565796f141a39baed8e4aed58e910ea74ec1347caf2774c0244282b1b6a95d49891d1ef3d652505c448de2181345913b808688615205f835ccf556f48a2835fa1a4038d2bdf6d22dd8ee7be8b56d6c9373015557c6f112d68a8c9f97587d30f8449853a3fa0ae49dceb1c511fc5462c02d00cf136be6cc71e4c4dcc6b713b961620545e50aa7b34642c1faf7a0c0a38532490d4887c6c6cb6c97a8a2f348bce20cea5d27cffab9733c3de96f8ba384bf5d6ca41638039ce707ee9f83974778788cdfbc5e77f913cb6c073d243793093d31efd672d110be71cc00c9ab639e8c13117313324d07a588bcfe3cc8c7e3675e5997c1d083d7f846f296b3714922f9985be9914497af8e7b0f786485d303c0bedf485c7b1b86bb73f6371ee89028a7ec4e3d8f80e78982aa8d92b7be67d34bdd02945ba7c52fbe3fa8bb8913110d55375295933b8a79a4bcc05bbfda4b4b25d03ca5e82e48b155150c670d8c00be810dd1523151b87e6fa433e92a8361ace2ec04e56e3738f9aa7b34662835fd571deac10bafa0cdab06f2e4923d2666b5c0570c71b6110a4cce1f62bd7add92977ecafba710bf6ca1c997888582531f26b4b2dd44a1d2a965a895d4f50216725b0879c0fc5e74e8cf37a997a6121e132ee21eb9cdb9b657deed076fd4f05313e097cf27bd27197de70d61ff12d60403d7365f42aecb0bf815738508664bc98f61f8897b2ce3b4ecdbbfcf61261038edf4fada55d38a9d7579e8d0469eb35d32499e164765e76ac5e67a54d6762e1b76b0bfece7478ba5d2bb5ae50eed9590bc3d083f89110edce61b57d2b986382fb035d6a952c2037c6b3b600d3f13ce6b3c1e52357fa648608e3cf05d278e6a8a0a0ca21058d9a7c3014b257ec6b0dcc100e05518f227111cf8e0bc19e5732e1382417b1630ba18d15a011725d825f835e495850d7b2929234a99cab3ea1deae1c31c0a2d19cb68c1e477fa8d637d2a143fca0db1bda918b9e997b94c22e5d18e9d4e8471227461309d6a5d978e9d4f1405fc38a17373e75baa713d1b979bed3864974417dc5d556609171065d2c6eb9e39f97d681d0fb8982a2523b1a08e52a09367bb0c11d324357368fddc7368651c5ec9521cb2591429e1e4a6c5b0dedfd27dfeaf0086940c1c2c65a4ae169e8eb9081ec617fc21ef32b648ebbea290b8a1b4dd356bd2432bcc090faa4a1c3ea0ae8c87bae3486d78fac4c8e946a0d0ca735febcc745f0738e0923473b493f920cdbb21836816665382f4b77fdf3d64800321c785f8fd6eea4a28b31b52ec7f2c7274fb8ce0e6b7234d3753a4b7dbf54baa0ed0649b7b472b949fedaa5cda9aea33239fdb3d4fac964c466e7fe005323858c5e63172790104977fef805f7191732f929077804f0718251c521295dd9473e476c7e563528c960b685c72682b532fb0248a2031e2348ada589bbfcffb7d1c9f47fa0a6eb63e124497b2841b3148a19a5e88bb47960e7eb58b10a5c3e2ada56974957767fa2b6749ef511b6b660e5aee715e9108df26beee0c4e01911635775d160e24df74f450dfdb45bde61e7e436611c7077fbe59cd326d78a9fcb31137f149cc25f9f58b9bafa3f279197e8b575b429d5f0607c209fffb1806fb7e569f7a8568694043aac620df593093d419b0191e9635546881fb5124de2839f86ea7a38766dcf8c9c03814f50b661aded955e38fa737272d63361b1c956f6bc3fc8e8e19ddb4e9a92fd19961ecc055cf936ecd421bf94220f7e1a56f4397e32dda8e190e0d7a1a09f83c2bbf71aaa50a6b9aeae98405d3effd81d563bc95caf4f5e78657083f8d3de799ea31752072783409791b374307318fc039c41f8e42043992eb45c8b21a80a0520b8f1626827271be3303436e4fd4651aabe2f298a0f4aea1bb5f64daf98f5ac73e9561005dd56995efe8afad31c5e402ac7cb46adbbf868e50deb4a8a79da2b4c2ffbf268d775a1559f06113b7ce749ada6df04d279d085701588be267a559bcc6853c5129e82d10f90bf214d4b5102bf641ca4ffb6b6f801ed2533d70943cb6a2d0328caa2a7b6fe21c1042db15b263a211ac92a247d84c335df2f64ef1782d2799f513cdf04a0a5357e049dc5afa145d4d8d46e8f63c911f86b9db5ba2822cf397ed7a2e624ea6a75a11f8a950b1ad87f546eba9b5aaf0021c246a26f25955af362208f7cc77928ed2e57640426dfcff210a09a3bf5a08aa5578d38e64923b2578eefa12ae1bddb8d7dbd24ba960fb846ea488b4cef67c2332ff8cc71cbc32265279981a1020f829bc7ede3f5c630e7359a1ea72b4ff06fe02375b5f0ed640b38b08d6a39595a63603880cbb7dfa98c1a4afdc0c5dffade666ce050304eb6a854cb61b3054765aac086026afab4e0517d0e3909c6956a37805c58e99740f2397fee8da073e9ba010005074d9dd494f302c8cc0a0766c7cb170116200a96920c9bfb69974a39203ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hfb9d913f9250dcab7c13138129be11251876c2ce04d37a5e5786ced01528f2f18217b7bb487528aec821226764915b2da1b64c57c81c3ec5e33a1b61404e2d179545f5d07eef54469fad35304d3c935526724baf026013ccccc25c3628c20c064396720f9d7d6b5185ba850b712f141c3d5c53d885a82e505e267b258b60c25dadcfefaca665634ebe4c93d3ffcc050bb940f7d55a9e74a4a2bb1e403419915484fbb36c46d877c6400fdbb819ade974fc39b70e76d4e594e16f7d61391e9a31b97bc050daaad8efa26de99fb8868a125a72203aafb2acf14dcf39708ca4468ac213bf44c1fee12db9aadd045e5e5c3380752aa5351e481288217028382fbeacb5aea8914b1eb4f22ecaa1cbad07e4248a81abc30ec336f67fac9a52b6d37f4923d539033622c1fb9fd768dc10a51d9a26dc51084eb425d15c70d90e2544f8584fd5adeedc00f69257c1945e8df93379fdc12a15f5bddaea9daf351f5254a5002c2a1db1e5a96f4d90523fcf2b18346507074d51bb16791df96eaecd94825999b138a487455c6fe710dc9968e5b436c15c0c385b70e166c26c75058194828b88109e553140190e6ad400be2fccd095e85df6f2c9a66090e712f5ea64ae6f6a78fa63972c10040f02a4fd3a568f76052850e6b55c630297c306745d39be9616d236e9fe9c9122b4e9151b2ff822111eb92e195a9ff7210ed83dcebc5129bab3fd7fddee12d39ff3389abfefb5778b6025ec05cc8d269712c87a1df6871ae747c2fcf2b3256eea1f2d2417574820657f142665859e87b2e7ac07b5664ae9c3a351ddcf3c6602d5529496587eb4d533d2980cdab655af0d0c4a0a50c2e0f5de1fd8dc5c6cb3fb2677260a7d0d6cc295f6b64251cf9f3b43fec0bf026c79aed5ab887330d0a15b2c277cdb3649cbd03ee27e7a6a9b992c6d4178b4f0a46fb227c078aec26b6c16da4f0ec7bad91158561dcfcb8a22f82ea6dec7dec163f76b2675035837f7c86dbfc5968bfa5b2300a2d6901f9129db2fdacdae56b2477674bdfe26124a8636c170453429a3dbffd80424aa206a50dca9dcde45902e52809c4210e9e13bd5cc0d6cb046c89d2adfa2bd71ea24523484c3f1518c73b91c5b6fbb646e8fc549aa727bc3f87c96eb15b74ff3d0bb5225f661247dd4938119d98300f2d9b160e4e57595e6e01f60e38f2de71217702108fa14acd218161a0fbc3d08fe06f192d6f3a10a09d1fa7ba83fb1d6d96f2c4f39aec19e802bdb9245b6f405452fa9d8cd67e882352a96dd31dff69eb053c7ca21e19d8337e3e8a97978c250e313e1cd55669dd7e81390a98c72a7d628361775d910b58b45db11402bc0fdedfbf992da0fcf725bff56cbba790069ccd92ea560f7790edea9e28317547f0d0e6fe17a97a10b284ecc98cc6764a1198def04de3e34192cdedade505ae077391472dd9dcc1a4a3173c7b324c2c1c51f5f4e3cdd628751c0d963884d0b5c3e57968311b6ad83cf5ed75dffebf332a2de07644fd3599bf617c6f5927a09c4ee45da5617b0367bc764e5510405f5472f993788a8b610e60a66a42d04cea31b70630d5ecc0eb1021c1aa2e7b0b1eaecdf0366efe3864dadde811fbed6c43d020de08a1d49aee0319af4c5d7b74d53c3dad046aaf401f89c1ae61eea40f68996d6ee4b580c8b8a874e12b810eda57d803a170af6d33a60f2d9f46d9358eacf4235db86c73095ce9efdb7222705da35cb0a1edcb1c9ae6d9aba44ef9d55178d8e22e6fd38d778eebcfb42ec74cd6af27644f9cde484f1b6dac5d0e999393083901594f80230861c8194924b432b151be98de303ea4291c324b2551a41270343ce378313b51628c449e950e57d5ef21d94131a42406ac3756868cea9cfc7c36ba48a91d9159a0b908b725120aa625692fe8ebb82ba2c7c7ecb4b524921b4eece1a3f721d8cf9a2a5fa8050cc3b4d358c06bf5a1f3c63b78838b36969c873140f9f94babf7f5d803f23ec2b0d806d499ab5d37f93b2a7d1923dd9aaf78ff97134e98595fa6edc32de78629620ce79b3a72d3136a59c813d4a6d237f92d8d3863fa12103661d7b594ae8dfa4ebd2530eacc10fe3226d98c1e36af3ebb9f977074c2b588bae5b8356003e3d4b01f8b08bf5798d191d1138199050336b7806db97f9e7e2db90d72a1ad9218dfdab8885a22cb7ae1c8c81546aa39db370f82363f24c35fdc2b13c5d2c8303eab84e4ceb5545574cdd989cd3c726fe2a23e2a07f38c41a54e478254d77eec36c375b4ffbc2da4aed778d0ee1cdf86a144af067635c70e4787c8b9f75db668fbd77d4dbf61e63fd2f0568be4602cbc8e785f8e6ec0a1495aaf7993d1d0ed53dbe1b4375c00f956d3c935c72a4aa1df2cf52564c5f266a2912d588d453a9d06cd68d98dcd982c94d87d8b83e185ec5c72ae796b6d94a68768ea160c2e66b03071ae1c64b25d6b49888d615ff481cc0e71831fb341d627c0b3bb16f92297582ea81556b71bcf4558cfd644f4de8574fac390668840a976185b6741a73518ce0e7e30feab18c63306ee470e35ffcf4e6c50261719bd0fc27988914af9dc224b2e7eb5f85bbcf4f4a0517fbded42f592dea0dcc6b9750646ffeb92eb9e3c5057689d9664656e99216e3f68ed315de8f78f82a6fdbc7bb32664b0b57f25de91219977fe175337f96e84fcd4617cd6aaa02d14fe71c7d082980a2672a9782e2d891f491166723c933f3c6e10e0e4a4d88fc13bebfd12e69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h50044d689739dc1f9820c629fb76fbf22b136990265cde68971dc3caaea887d87f8b83b3a44d5f99dca16e7f81b814adf27f4eed2675c66f9c58c2fa2efc64f53d1927cf3023561f759929aaffba6edf57b0bbffdf44bb07de1f651f5843820672c0a235494eb4760b41c0db1bb1257f814474ffdfad719480b41dd0dd841f0daeb9a6392f1f927211ff153500229bdb5842ee771af49bd23fde67281ecb4742822cbf934b6fd7a591adcd1001fd77fe6f21c3bc5c68d4f72ebc8c088d35b4f4b169638298274556bc5bcea9bc2bcb5a5addc2baa7d8a2999d2d275be5b3b2fa377f8a518db654242c533ecab06265db5a5878d1c0af5e847e557ae394a598d6a0df40c4fea874826f69f8c2c8207683e3c7c28e6a904ec296a10c9409e993432038dc2d117a529afebd6f8c3d3071124d075c57a3c551517bd4b1f355e8d91660d34a74a3f8e3c5b8a8f0fe8ea31516f759da591dafdb0f9b205d0e388177e930b4aea4670581d9ffa60900456ebf46042d671b35493c812328b268b0544c1408af202a97cc24d072b1b810a5a99d2afa90c21258da420bcd7fdb249c6aaa521b81be54ec5c4eb27ec5859aadcb37fc6b414579bf9b57c67db4a794e4b1345df19359c4baf0df05756828b372d765ab703c48e947fc0d7dfd10c8d02dc2164fb3df6f9099810125680525db765fd8893d8fe2b8f0aad5c5914e8fd24becd9fb0a3c89478f7c431e19699315f67cc328e8993fd322705cbfa9cce8e3b75fb323f74aa6e406b4d49582494d7c1a98e788cafb5526c338ad61c321b961b04fef9a41c1237888445bf25149e2a24bc709d5924e7db268cb4e99902a14b7c008df75c0f518a89453fb3e61edb74901c8989d523811000f43053830cfde8989138a4db1dee374d68d7dd8b8252456fe64ae239202e7d244be3d50b3b6af56bddb4ef5cf1eb23b14912439e6eb0069bb06df68b60994f3dabb68be532217758e85f405b70114b6d084bf29e6acb7d9c6fa4abaee5d8939824eeb291b8e30ad6a3ba60a90d50ff84ad3cb1c2c44b44b2f270acfdab8a84379e57b90e5a91faf04713c232bc787de35fbbc017cda3382a0409b1177f7d5212e86519c182549a76022dd19e904d95ee5f37a7e7260cfc927edd6c0021a0aa51ffe7ca6aefc1e1dabacf1bc3de306932db0106e1db7ee595536c3349a7245575f02784ab3effa71239f149f5acbffeefcc0af1325785d4b5f93dd9ff1c468ace38c5fc4f55d9359bc6f0be67ff90fcc4a3b140369a372ed825ccefb5e3e3c9c15a07b2f85453eb816c5546fbd358b927bbe02f1916cf9b0df6c9e096027efd370df2071f3335bacc6e261bb0fd31f822bd2476ba66d8b0f5f8baef05cd4e55c5ac9f947770b5e73ae65df8670c6b9a6a022170c1f147e8dd57bd4ad1dbdf451a29641e4909d85850a89744d3f4601161f2ddf16be9e38ba26759164cc4376b04a6abf263d6030af7a4bea78755eb30f9affd583cab23539cba60c53ceb1d0a726ef896ef8bfdbbbe8be588438ae6fa3f29673a677dccec338d529bfe310ec66c85f7ea38449c4d7ad9c37c084d5098addc20ce536a114cb28201bc7353546ca112381ea993fb26edf58f610bbdc79a915a4ed054ad2708b9ae41aeeec6ec6000e9e96a7e9fa647dc9ac850534372ee5b17ff7bf27da00caa89797183f3c30c073600b101208afeb15f429dbe668922a888851f0bf5dca19ed52ccd60f999cd4f98af6ef442bccf05344b2093dc99a30c23d2660614f0144cc74865c891928121057758100b695ca3114469cad60920a2f28444159b28b27aed10f3677d4a2e5805491cc213539652e31081c723625e5d47e7be531dc43fe9ae522b8e7f9cdbbb7fbeba2710814224244dd21d2d4f9b64c44e87ceedc2817b103ffb7429057d161f7ea488e72d7f15449f0f65194ed1a93959101bc6e2868bab8ca5cfbe3a58a23fb4e1e4402282b8c8eb6bc61ab35dab3c3a8868125487a6fde8b44a9c5ff15b6572975c901c1d9bc1fb56268730ece746cfef4f932fb483f2e1ad14b5e9bf8b17823507a17e4d0b1b04fb32c4385a9b2c60574e917ae420c3a0997baa163c7e7b27347a78a09dbf4cc463d84556bffdf74de612b025a8b42c73db588edfd9b148563d4a568e7874de741c5959d1bacd63bbac743d36cb277153c592916ad96e43f4beb35d2544f368755da566d0b4ce4a5f218f184714a52b57c5f2934ea3fdb356554de9255fb1a0f0f22652f98ec5879554abf6cf5824ce64b2fc83843f4f9ec6f3c2243832f26993515ebdf92458478f40ae59902ace038b24306d5f2c8da84ba17a6f934301aa928a6f7779f0dbfd3f78247b347f30189d8a1415db91219c3db8e3085a0dd447278dadbf1abb71da343a78ff7071adf9bf5b2bf9eee3999441d5cdf2a46de4907b201720c6180372a49ae9acf285b020e1d7576914c99ba4eb749ac82512b113dcc25289ea4f951b0df24a9bb3726a73419a0bc1553f1fb30744385a84d70133dccc53dc13ebc955054f7fde7839c8bbcc8be1aa2fcd4b05b65363d2e61b3c21f16ece01b9d53ac1c08704d13f182090bd89b71f650de29a44a991669d2e0962c7fd4a417b0cf3ff77d180e30e272a263b93921f379924d81404c85cfbb57b2c6157a44f904c083555223587b362f02f65a772d36b67eac3974946ed751f431878d5b5662c37e94f8d9ab88601b86b5fd975d91aef1ca563986dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h99b6c765ac8015bb3547ed495e92405f32e32661adf90e595638c4766ad251183e9d8a5dc819713f331e2abdd0e70ff5284ada403bbb9254a5915d403932c8f1d2fe3b98776eac1fe6f42d50c269f2623a07bc8775a5e19de7b248c2dec2f038e60bf6ef0f7dd3f8e2babf5106527410792c0139b2f20b95b8775205f8910e445a39fb060f7a0f718d759ba621f1f74fae6213a7ed354889346f3aec835741352e56cb016b862d92ba2ab8e5a06555afba67068b477f0cf5ca3d4f5a48a1fb305b69e1099f98f44e9c1287597a044159f73f758e7719eaf01071787af12ae2a7a2df3295c2f5c474d07b4788a8bcb9606df405666536c08e83886238e09626e58de1c625dcbfc686b7a37c572b52a07ddd073f4bebb6ed071508ed7f1196079e3cde1ab28b9951b9db7bfdc3160805435e85cbfe72f60ec1de473b0d2b7f530e1dccec9d59a5701ad6469057cda7e029471e24f2dec2b2c0201343449689bc546908f27e2fc6ef2ef731f2954e0b4e8d9592cc5ebea11af53ba298c86afc6faec660f4d9d2006391f8852d544089b3db4692b90be703068cccb7cd2d902b6fc532fa4a20dc756e61ae88e6faf74672199edc2979948d14afd15e691e237762fed0906b6d8022959bd71453ee6813965c6e5a2fc4ca571e7a126db9e09219090855b24dac53d36a7fd879948b02f7765aac36418521bf599f56bb53b3e14bb59e1a4b5e21e449271679e5698f9a8613c19408019d8024f2385125697698a1ee2453bf9fec4febfc4951ca6ddbb646cc3aae370d038894654e8865f9047b9e5e43388968073c04fd9e3a192917dc33626380ddf72f962285af60b9418d3f14d06f1cc35b981080aec8f1cd03f051e4f81a03e5edaab8f429528a2a70debf82e653d8700c0e657a1dc3dc705ce8e4e13a344a4b6a2c086c4bdab1dc4bd00dd04dc32db2a63805b50b4a61378def701c42f05209bf53944e9a2b0c06adaeb703574090405284f05df6c5b4a063b17837c03b82eb30ddb94c68f3e10fb9cde3a76a5ea65acf1bd6b7bc6ae23bbf974bcc194d7c303c7e8db1560101482ed19045cce12afe65072e4517d397184ba47f063f8cfd1ade055512489f72372b2d7e4f95422a19e3f54f7f7b07a5c3b41a34232d55336880a2deeab7ecd0fbaddfd8d7ae6238a0ab8d6fff58c8c642342b95532eb5317a1f17f325697e709125e57b04519806a32b20d204e36625e8997fb6d4451aac40ade3fc1aa3b9d4d93c80af9b276088e98736d22daed15fc5836a35b8634a588d093243c873d3741ae88ba9dd3b089c16eae90c9442eea9808a524f51e23c0eb95ffa59598c400d532616bb4bd9bd2c826de68fc1204d477d39ec3fb4b9a5a62dfbe9669c7b6590faedd6dde2ac00e90cc40629763410eb7c461f874afb29210b56907d01fac6cb6bfaefd6463fa20536a91d951b1b5fc68c38e8261ac9d1030db9e2356863e44e426c60c13c21858ac981a520cf334161927b277c69595ead2b6c6c7aa1b77a6ae1944e5110014551237f6793e576725b66a9a096a2ba57a24dbecff063c92a85b055cdaa3d6227af17bb4f413de94da7b6d92457c18c50df16cceb967d6b31a41f53b53632d1cf69bcafca577aec09cb888156e67d8501bfdd4820276298c53b6927e563899f27fd029e7fed6e70777b69b9ae0e22ecd92f3b77f6ecbaa59f796390591509c7cd437ff9c8baa661d4bddbcf2bb658f43b1e9385d3b715e7971027332f55a377156b4e1aac2f30eb6d865a0b59f1d6e75979b8f183c3c4a09cac0921bb85175e75df6a0d55272040e8d6f1bf9a20efc51871f262e87eb4bfc398135c8244061a017521045b7ab4bd715cd22010f71482173f92df8f4c4a04197518ac288937b0de9292ded1a047db25020aaa80ef0baf4348e17f7a9bb89c60553864362e91fe2be9b7486fd38e62aac11e4e8c6ff76f91ff6eb2de05d406219b7d6e78e0773c7dbefe1468c543ae4e7fb91490729155bdb91a9b05616987f104882afe32b28288fc77a29831a51cbb45f8d172a9a6a3520b0a1ba919137be9eca41e14ea74a2a16025e3cd4d177fb919f5872f368cb2fb83b540cdca8f817457d6b6ace94b83dd3d317ba261a0283174f102435b0e60636059e95b280f308ac8e1a1f8aede793504a092da026001e51ee3ea7b1d1267c57cb37ddf3f59889ac89ce82eb3f35245573509e8cb19d7f76318440f7e37be1db5b7f6ca8e6be09d70fa47c30c7e335641f8b70738f99f6caa2a5fc40c33e6e4e9494a5b3ae53e78c246e3119d44320a61d112314ad371a26f7cfa5e884da6a53808fc02aa4c75ad9217563f6a18d70cd46da53af23a0bbbd5666a9b9f256ffc5b7aff52434e13fda7edd3c6f58b838bb6abbfd87777cc250658fbf34ca09e2f051463f0e7abade665600b651b2c4bb65de68a94279fc238e348205d79d53c6ee76fa5921abe18f4f6e4213d2d33fc49a87bdefc792770f6fbe2fe508310da8f9a12a4afdcdf5a9cd35a65c90873aa75262e098902fe5dd05a69b6f3355b22442cc789eaaa6128f1441c26c0c8db0a04cca62a51ecadb17bb5d8a863993488a3b695dfe88494e22db6cff40f04cb9b874024a54218872df7042e4c35524af3a4cecaed13089834eaec94ed7809b5071f515ace5d3c7e9a360d1f97c39efbab43466c2df182d39eaeeea93290a094d41e3e7b1c673bf157175e96537dbe9d4c7c5c5b00f48e544238;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h18987fa86d7a5fbc69ba5866ea45bc354a1fb56cf3b040c6e948e94cba4ecc42d45d2c31837a462f677aadaef304ab1843d0a0df32dffa70d85c92736405f0985f77b8741dfb138beca414c64d52bebfd1d7e115d38ed728e81e3dfa0fc2ef1775ad190044a97dd5e664ba5fb29213929656aa59e778701ffc62853a1ae4abd488593524c799bcf3e37af5bf7c1a177fa7d0e2fd2e2b3862f3f78529ea53b2af06356fe9e29ca3778d418c9d2ae3284b0774120f8b19663dde02fcecd3a808661e11dbec0fad5c2ff3f7b0229296078fced67ccb470ca4986cf5650e93d45dea9b2f31f49800a9ca545e0124a0f1018cf6736730194c57ca4082eab0b4ee0e3abd1c4f623b17a5091bc0ac9d826354b44914f51aa51b90b66ae40b81f86e569b5086fb6ae6c1d2ef77b580c425f79ebb13b24fe7d76394135ae82f34542ff27c24df5dfecb13060ddfef877900877c2c5caa0d05b3e2ec8a4e2e29d6153cdb684f6cea5b9d06621bfe9404583b8bf25dc04c687dbbf1a033ad657d3c901d77f50fe8f02d07b5848dc3132cac88d499b794230e352f26aa446fea7eed19935883d9e331da1396a954c7e8d95a15474d7d443044111b07e7e8cf58d755c76b12700d5a314ddb5c0303c4ecd15f29fdc47922387bf8e5346ac9c6797d194b17a99b44ed9d9869db52772455097ae7df7b3c8a156fabcea0020d4dd08e970798ce0ab9413d8cb3a90fbb5ca48aa39750b39547a4f264f18ffad933b09eb3870403fa4f4cef98fe7d92d91eb521af25bd7012c44c51c566d9cc1f30bd17f36aa48674b72c67169026c9baf73e42c804bd9a1a43e6224c2ad4ac1b06118528574a871089be32cdd5dc36097b96d99415f5563056f01681e405e7f0bdf7cb55cdf27b2859232ae5e5419d9a3e559a0e533de2eea1d5e8f18431095859bfd9dbda0f84b72c8d5175ff23a93f3b0e22ee2e7f2c9ea0041870ce6a9c8e1e1f2c96aa47e5506d37a7256b81bf545e51507ad734e32e59243dc5591e280a5322755c1252c33b5089b5df4129e6f6646c0e05384e20b4e2c4619c1133c1cebb143af6e20f504cd3d4c95733e8885ae8ff4e31920e350f81bf2102864df79666db19e6113a1a845afb9554adb43813147c6408e367c71d2a209da58b1958e456e3e01446efaaec396e5cc49b53e61c6ec3d724c0f7888c1278c0dec8fbbc12628944430ff2f8049089827831de54a4f80469f38244a0b8af6db6d485e708e38b1ae94753ad429e5012a744828a10509a9358e1c4805d8c679bca3df7d2ce9b63eb80373b016729e0882bf2b11ce68cd6b0837a250534e06c658172ca18f93d47d4428e6a2a398e749811f74209facf789adef2c929809398f89e6fdc9621724ea8e274d01faeeac5a2ba79a9b9f555478650076332f8d47884726d51195743fbc29a21feb0de6d1c2af838b9e2a04fe242737486719937e5d34f23670c9b225e64c10bf011efeb206745ee61a5c8e72a5facc1303b9fb3d84617646e4acbb2d1186ba0c22f542f2b8bd691c49e4b057078844d652eb29baa212f7226c59c65d3b02d575cd4493458534e262e427a17f7718a4cadddaf2e00f3843e0820a0a92a75ee6ed4a435c236cbc620ab8ae4e82836a6a205b2d1695551ec7df7828551ca1d1ce825df16785be4e5fd4e76a2a6d807379a1c3fa6ae4b589d5ce9328a9003b13fe55228b0a271e73895d6bfd2159ff64854a9a778c5c7f89d31c6a98a9d41c11378ff3dd3252d9498a7ddf92e4e72e3f7ac3aa4e8a0cfd237b5bc22754777237f6415e3c063844ea81f96e6bb05fe10289dc0dc7f05c29e3211948d359ee0c176b7ef975b02d8eb7aff7887b50766640ef613bb244fe813ab42fdf0c545f705d64eda8acece8a1822b594a81c4ba0ae6e976b740d200c948776406e073986b61e337da5713f08f1b0e0330d7fc0a1d78a9ed9ac6950a9680d5215ebf13c4517c13ade38feb19e02784f3bfe7a35facbc85732a0c6ddb66c04f56296c956ca144c710b57342ee167c892b3d10083d68564cc0d2cfc66533a4ae5b6d7390f8ed17eb68ff96ecce31d27fee51800ce884ff55864ef0b936fb990c8129431357fc8e03942041048139fcf7167bfbf218ee698dc133b4dd12230551da1f32632b382d8207398a8fe07c43e29d90b4c8e861a387eabb7ed74e16cef93fb4fbbfb32f43e6b0a0c3055ca2c8416175b50872f1e06977249077eaf0b6bbf874ebb8be7afce3a99e2a09c771bcd81c6448caa209e8de1efbe10f98b0bfb57d3f7f4da3364e6336b74585e6ab3667f300ed92eee33fd71eac1935dc7516d0c23e57dc10864fc647e673ea83d09d93381d0c1bb86893b62f63fbe22e9aa198e0a95c1cfda081b33ad38be3805e4ae53eeb4c99a7c4fe9cc4fe1c80608b9331bec704640265a69490f14544bd49d86238c86b5c0ee314724df39123b2b769893b58d6c7ccacad341897342172d31c962f2b7d1eff1e8b08acc5d226df8e73a3e0bff0a5834550a39865aae92716986a1a06b6718005b15a845674bd8dc580413cf044bde57c9071251c78723ce481fc78c8c7c897d90bff62e7107888932c01280261c782d3e7e89d2c7b3cc485e6ad5844ca0d28a85f18aaa34ce495b93a2203517ac356280a7e56952e6373a9ed7061a8d5787c38505efc0267414fd0d03b75d40a037b3746058d18128071ec10426ddc1672d4e340c6fb70009e71ac51f1c8c35fb15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hab21f1450940ae9e82ed290876fb4a7beb7c273ca1cf62351b239f03e47c97943f1c5e8206115b7f5924b4e691a24b6cb305210db7ca88bdd2bbaad19a22b63f967ede5b010bcfc83a477709915e14bd36e618d715654c5e9a08d8339274875588f732cae07369be70fb6f6bb04dacfd156ec1ba69855b9cc2c67f4ac2f5363905ebc7e7166ef73534cb1b50f4d52c3eeff3a7c1ad62bcfbead724b449eacb99bc9c35c625f46fdde929dfe3ee4723524e271da25efdf78b2f4310c4e50edff12834b0b1b1b8484cd9af9ca8b9c3be4dabcee8c383aac54d157e41ddb9117fec0f8cf8a359c69be69f536dd7dbd63f6278d334284a149c0ab4aebf7f47b2d74554cc5b248b22606723dd889387446f5412cd18d107153a6f919ecc940ac39a90dfdf80a294e408068163f551841ac6923d7aed4a7431abcb1071452c4e0082e048db03d26908838bfad0139f7e879151923b7d593eb6af3cb8710c4d7a1a471c4c6cedaa8845201801f0e3e145e833768e0782b3aef9c447f05127cc32eaf9f1b6f398c6ae45f1befad48b33d0d6c32c5fc4b3f672f26b3f7430237fc1af052e7966de3990f30cc26ae137d8f3cd2ad275773b0c2ee3c1748af932ed90cd75aa6b51fc35a1b5ba6ce04cf3ec3d00a68343de15cd34867c8ab605af96271c1ce26c1b1f3b421b0d8b83895bf6f4036d8d16d9cc2c4c4631ff665f96cba636789f7787169468259b10a5b146b9a0294fa6d529ea2262a6f52f1aea7e224bf39343a67169b97b12df5e8eed186944ef13492a96c71c08ec3fccd1809e88cb54d42f2990a3ca2390baf707029902970f23e80297a7fe088c130cd9423010074d491f44074deba2c9e5a675d03dd55010e65d7b05ef4e00052c77de287d0719b1e6290ca8985847005da8a0b2a1e3e943adb5c1d2fef34894d3272a9a95e1b87116fa266bd421eff2853b8f16c314acb1412775f8d2cf07ea6f8de80b2310f26798e1ede5a96248823ea559e8c9975849aa75aab4e22b2a78d0cfdb542a4b4c35023e4b58a3df1b8c0132a32d2333d5be178bcbdc0446c1e1c85136d92832cd7158122cadea178783ef1bf4de545148e97b09b8b5503ddd70b1ebfdd3245fcf42bfac61ff1a4aa795c4b21d992e812490386d94f528d091333e539cf183bc8f4fd27f622e10f370100c3a55b32a93f02927ca90826d8530cd5012c6b06bf788a08b12afdc41057cda9c683878734fbc409e6ecfa84d7ce69d840789574360a4a60ec5b601c8d60fddf8a773f9c4e5971497aa03ceb6df8c9147ffa39d930004abe993d9bfd03ea3fb2dcd6f0f3881dcef724d82567560aa40f1d992e41391c35094d9957d61bc4ee99ac29fcc6bd4bd4cd3fd1a6603a5742d104c41a7e21cc0150acaef1272699c2458c236a6fec717aa7cc3bcc572b6f8441476fba6a3117f166bf92874d2d4cc9d80dd4ae451773ca620edeca3e4e6850d2127e395016d4a6cea6d2fc427d610a474a6d5bea380da0f2ac95ea9ca9ddefdee45039bb610bbaaa87ff7027ecbdf7523a586b31f32845d48682f1fd23407ec81478d89c8871f79d826c97f69b79414ad5c77d5c2832721f271441e87ff3f412e780b1782f7fa8fd6acd3fef25b19a35c8c1d94941839451124d3bf6c28f64d57bfe8f4918f1d6ec73b136afa8534db4e6c2b6060bdf3e40a6190d0f0457b12e5d189a158e7b376740a9b7dbca47b2acf2dec5f6e136bd55a576cc13535bbc078e8ca8b1d5e0d507c31012010ed4bf10f04b1b59c4da49a5ceed6c5f3e3073d55675387d14c83743b66f07960f251f0ca0d36726a58b2a2159ead2f62ff00e563fc62e2477a5b50fea798119bd0a8a9d33b49d86b8f8ea3b0cfd9bced1ad17e088a102f96a6b9b8677a5115ae4be1898bebdb69c16a40aa24652fe1eb91cd5f6719bed655991c8dc67ca3edbe4f936a2817cc736c6bd010dab758efd1706308cff08050038506b0d08edf21edfa3147fb22fff789248fb46c089a98d955534c0f5f4d635fb9fd0ca91e89e7fa083adb2623f61cc4273b5e8278dfd64cbc5a966546ba593a66a973bb3cedb1e1c42668c13c8263b9383a28898ad242377590d08b252999f028393c301faedcc55df78897029e42dcb7e5311815770834dc5b430e4616cba1db0f45ba0e41ab45ec09f35b12c8d6e360015e607e8e4536c57170aa877e2e24323cf52cfdfc28fc0e502001a5d24bc5910ea46bcbc80f8c8ab12beaeba63208de075efdc000aa505b122ce384fa5bff113cf401b1f6d007769e768fc871a2b7cf906674a67cb2b2348919e3c62c82da621aebd40a914f8a98bcbbd59379f30edb841b8be784b4de69a0314532efd37916bdcd4758213b6c1aff11be080c96e18340b0d6e3b83f95d14b6fe88bf09b0fb720bae20d9cd6c26fd0251cbdd2394c2d661f35b1a7d1c8e2e4c4dfca622884ae285a6c869194b84aa27f4c71e9e9ff6972a4d2dcbd60fa42a189606e09285910c577b9a9078cb943254d5d975164f082ab512930d5b56e5d3fa7c76eaa9d200493aeec724da4e11941933652937258ca1cd9ba0a7f4a96bee7a3360668707edc428b972cbc2bcebe83140d6bd3d3c70c594bc9604ef9c9df842a807b8cdfcd22288314b0601248f3eee2ef81972636b6fc048f122c3fc8022cdd4d46fd15a7e3d44453d11371efc8b38da8d6ea0bbfb7e303a71dada31c70e3b5266e60b6706797cf11b2641a4fdf5e133b85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hcc34e0a0a4ecb3a645258aa4d02d1ca0c89779fbc61fc4b29c840a0cab5dbecaddc1a4367bcf50753295aabfd06a8fad6feebf67da7947c3b5e01330a75be40029c036935a763e194a05ff5ab40a4985b6cf397c04940080c1c4206a05a451847ab12b79f1771c4574e521980d9b8ed1b7d0e330132d4d565acb1d5fe088a89ae6208bf618019963155a26a0bd2af7154cc6e1ee33970f858573b1543d48f9a66324a8803ae4651f77e5c5976169411560e2c22939e848527d9b1126c1d3a73a1b4f6bf8a9f141b503fe13de3d39df376a13f0462e55e40d72e8882971ea9f1d972472033977977442c1488e764bee4de397a4edeec4cced3e2897437f29d6872c20fc07364ebb01e7736a52e3fdf2e812db84d920bf5c9f33abd3fd1f511a58816523874a606a31468beb8338979025da57ccf72b8fac959dabaefc3db775490aa2149908ff0db5fb9a5e078a0cebd26ae968be00c940038b1b2a7174b0bec9e2b27b6a9bb2113cb4c723b96e51dfa20c441e477ee18ebf9a2c070966eaa4db6c5db89179e2f6a5219cf4be028d2f490a164dea4591c59296c6617719589ae0226554097871044e550ba4bb61c0eed18edaf775b31e6c3f20ba30a2f75ec0da9aa70c763dab1468e2cebb5e26a00ac4a10f0657fd80408125d4c1d0c671d53feb45b50fdd5886ff37cde9dd557c8ff25bd0d64ef4c9b658d23c557322d9ef15693e51ae72bf33e4ba3db54c4a85c0a53175ec3fd73d3d772cab3b8d3abcae3aa2ccce7065a7ae3ce10f5f752243fc59aa41372d509400d2f87b412f81aa09e15790b90877e518b27dcd1f8e6c0e40e3fd7070328b940cb8198170d56c1c068732b3762f009ea0bda36bcef2ea1f0bc33b6ae1eef63096ac7684285e9d02a6ed2b072ebed55129454dae45cb414cb49769d1858ac723e54bb4cfc2295a56bfb1838272ffd3407c6ca6ee9f83fe34c92a6c9b6790773c8d4ddb99c627c6be0b1924881989652d0756b0b457f8b72ac7b395289bd61541b71c66d849b76ad5b604b23581ee7a4125bc903b3589775ad10e525d6800dfa4415fa072860b3fd11a11b394c27603ce7541965b4f9d7704bed3eee862f4cb2a369263fb87ee413bfd33870977ce54ff54d805eb93dea5d4683442131feb3c9c13c4adfa1fa5f30f2a13b3ba06a0a6c7a4d93839870214c9e8a10282778da143e4de05eadf88876589cc4a82923ed468472426bb46375a00473c4e0b9155221aecd71356ea9e3ec641122826d1d2180a54807c7376fe9d057dbe003e4b961ebaa06393094499c6dd85bca6069f8fe25e78ce9eb3fc4c7752b3c51cece13d6ecec148a1aaed4132ceda0b82f1e5ff3b5ef6f605418ca90229aa9cea25b187c052109633b9f04ce51c948ffa4661c65274f5c967c25d36ef14ca607272d7f9a6e0d5776f24d18502e2a8ff421f791b26753c13c354d0d745cb01116c33cacc514d538df7307056c12ce90c8d32ff9eec27b6412a48e71305a25cec3d91a689610af69ae4a152dd31f393ae1965cc506fd1eb323e0aa9dc83d3751b9d131b25a956c088bcc80270fc461782b810c081c7b556bcb3014b803b47e48548f7a5e01c75321083e6de36dd4cc51a7ea673270e8cab760027927a4f42488593e31101e64b726668326db6738a433b68f1e643b1c30127a67fa5c50163cef3b52d507d242ae45d39b16d8c4b3250750f74f6b262bd88d4ab1e9db735b5c7ecf5e8f396ba3fd1cfddd62e52c652595b0995f484e635ece06ac506eb4bcff61e7a6a80e2b1ca3f7e9f355645ed9da16effdd085d0736713510be941bebb18b4b9ecb213675d3208c79b01bf4ce17de1904041d5a1923c453e1c9d7824b3c21a7e123baa66039736d9ab2529349fb5c6aa7539e4fad5b02e9faa89a49f50aaf422a5cabf9496cb18157f742458d1ee250e96ebc00e791c3bde36feb66a065dbe375d5dce86ed6affcbb94d2aa834a7e0f7f460d8958cc8b0be93f495e5a18b7fdb0943ae94e23dafc54df8cdfeb4659e8bf9a626ac72c32de33e4ea661212764baa8ede83faa9e35379b5f6922b87722c117f7df6a5332f864c877c1f321aa0d772d16993ec5889d06b1f25f23d7ce2043f04d9485de6ad55ceb8fbe94ecd236201ec3493f90b39dd32351a7a20d98fe8800d37359037fde2e09214f09ac29d69987f1a6ae182b7fb308297a8eb95f363070dcd8a80fba6eadb1aa649e9d54cde440c688c8fc7ab0258b6685bbd7730e0d55f5f90c86328271f82aeedb0393db7947c1cb7e14e93963e507a400fa19f94ae68cecb6d82e0f78c09ceae2eb5e4f16700a4ddfbab6d8f7f53575e626dadd6d4707641907e002029808235ca8b77db28bce755c6893b15663bdfa67e115630613a173c7965415f166f5c259a7f795d1d33df2f54531068facf815cd6c3f2ab287d78123f0a0f0fbfb3791a6351d4c0e1d9a2380b588ce80b004183401df44fa4b3c2bbd1796a6d304d84174cf3a772ef2fce8c23535d280d7ef918dc864386941878d86e5d4becf4e2d8bc58ecc8d18cc8e0baa977576f81613530f2c8ef861609c37ec211e6a7d053c5e690d4576f5abece6c4487bb584c6ebe8a65fb7283230f34b99b8ada2752c91c6b3a4a516d9188b1331d144ba6a932b1ff07790e96d29368a4a96c3c8d87f90519c4e570647e560bf66e0442ad273be03f76cadc34e1835e4b930a6a5b39a847cd8e3a6a907b4468c9869159e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2a4b3f5fa665cce4ad256aae39b2f8f69b7fd36f5d530fb8a20b7d8d5baa3742eb553faa9a57c8a2e8e735c34eeb36e64fdc4330eef02b2789151a5f52075ca7147aba47a6548aa7d4d125177c4c1f29897cfbd611f3f891610becf9cf46e117f849bcd09e67fe27cbd7904c91dfdf6fa3f23e5610eeacb1691111e4bda049644adb4e4a1fabe5966ea026e5bec53bc3d0b4004861596f9a708969950521b80cbcbe94eadee5bf59b3f2e3ad7e7b7bda71087b2a0c31d08b43d6c6d4e969a5af19dd581d71bac2c326baae9e36c9040bdee31d0456b36d7e2399b6fe5aa474af009fce7dd01a4dce62ca1bde9f334c503f85bce3f5cbf162474110e9f90d3370b168d3eab81f7cefd2ed6f1eed16cafd52ee7988257f1b4772b0d8b77ca34a639d5938995d017ae22b707f62029bc89f01795c38c2f35b004d54873493417151557433a969502a5a412f12b96f894e440fe7f395aba921f0714d373740175213b63b1867a9b7cff4cd575a878aac027ef2d2964934d70f8cae7f5efc42b86c06a4aeb72dfb0d1403b59370f3ea93e656fc73821d933d291b5d19268327b4b794fbb126bccf380d1c36810dcbd0744452a9f91d4256d56b86a46296114a5fb32161c130fc9736641d47f45f56435ea2ba3dcf57ff01324d2fbb033ee7d9c2b89128e6d0cb268c52e0386fe19e23ea29d5169e7a35b6a4ae355b8bd14b453030aab62a4427ae37df68bdd10e9c1a625e81010e72caded64d4e4e5c6ac4ea3935b2a32dce914ab69c175f40c4dd59b2a8fb5583d2b44e591028ce01cbac1682e79ff15d8b613121668fad71ca03a9f1ce5049664928229553658fa61515838ea79508fa594109ccc696bfad27ed6cd608d8c9309f4950a6a98bf25bfe9356e7694545ed0a9bd136c4e77ce553e1fdaf195f5599c32211df5f4664646eb35c18de86257762515474e1085bae02fe3b431625927a51170a2448c5a98168d4ef1f6d92fa45375f6b584099e98c6b7667697e3e237b3b1f7cd2da014cc3d80d2ff82f3206b111c1fa3acddfed2623368055da4ade20d0b318881583b0c8cde14fe8d0eadf2c466d4405e6bf0be63d3dfe28acbac7d4cc02da0a5e1861164b7d8b175bcbecf82289b6ada62949ceeeaa8b58c9c64dca9eec3fa84deda010c23007a010c58d999ee0fad0d3753655413189caa1bf03a4ef944de26834cd88db8e392fc57dd6169fa8beca1125fd82c82d5074aaef5aed5805d8880f108ede6c6a33ca83f0064c0edaafe0af828b28b7083224a4e3f13f52719bc165df243046d134ede0b649282e3b560ec56beb8c23336814ff66b18b1e26abd5c3ff42d73c3899bd939d9ff5282e5f21fd4d9b510a20a05ec949c402c1f3ca2b0bf21c9f66739fb8d3e1b1356bcff7a40f111da5464834f1acffc8197ab5a21e9009a6224b634224e0bd22f9bd1122fd5115e9740d15d4d3421364dd9090c6b20912a84bdc1edb9d6d56e11db029da736d203ad6cd5c361762fc6545a911f046d4136c2d8f003cde3d05003d8694cf7bdd1a79008501631d6d00e55267c5f52fae2e3543a33e7478b4e02b34dadd5a7ac220d0836fb661809c8292c60167e1b2c5e1ce6825cd91dd60bd92d8c7e324c8076a328d9750462ab2a253afae123dbe696de6f68a88f1145423e0bdbae5fba9945098b60732c18ea6391c0128cc676821b53202068b5b98829ac9b28e0ed009621c53a49b91a7b9b7753f105862a28f65d597e8b4b72841c2fd039ba2c83f35a28d833d351a25868131c040f925079653b12e49e1cd55b4e824e1d7efc31a3cd82af3844b9e48b786624521628ff65ac864f177646b42f7160024983d3913890aed4bb665562ab214f5f49c60da32a31807f36b426e89fae6f33553b05c47bbe89c25add999a45109d49d52a74f6b2c9c54c383cfda994e396c04ea1b52933303191a9aea85e43d12600646ae620a56861019030192f88724825bc2e837c4d3e552c88fcb9fd4770307545f7c2aafc81eaf34f3286c99548c3889bcf486019271cf082623d5606067315da22754bc62495a4e545c5a782d3309b4d0d5d58a09e40cf62e4044882c9d6dabd8438c6c7fe3f1519a89e6e2e0db90730d5c2fc80cf72cacce627a9a42a5fc6773eb7655169b37c23a9f6296f3ef7720314f2d8abb3742847d63a333a3a60444227901bcc966b7d4b1e46730af5598154777f57f75829dbcda968a59e303546d9d9e67e008cc7f62a4f9c556a2cca80b326e1299ce740b3d0d052a2aebc7ab174c9b6ee12f8bffaeba4d2e0f9dcfe8fe56567136c2b9ac873f850597db468d74b9bad4e7e556973102738230d108f5fcb2fafa3c635a81249753216776c7769ee4b3aada431740f60c80e399b69265d122347323b225e52ea0bf741896628e2b84c86d40a75e46cb7d2be3bbde0109a83c17ab008a75d74d99b78b870ff340eadcc40523c58563cecfa626163cabbac7047b5501e1a3df698f53e9db1cb7165265c3018b34bfbd62c652a293c4889d191b23ec728553d20527fae29751fb90d3681b99a29ffaea2bc6433325708559adbf95567a3466a85a5e2c1f6090395f5f8f9cf59b775a38c07cc14cb3c8969c2eb0c8cfb911738d2b97ae11972eb933d3ede73b0740e10dd34bd1a8ed4bea9180510c6f0dc15812332f54b1c20cd33edf8c521bbfbbb31a76ef6ceb7ef3559347398628857968cc448ed56958cfc7cc088c8b9f3a2a6e41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h43828fb5018816a696cc5b28a576e1ce0c02063a37fa773649e54a0cc54560dcba614e2f6c046bfd5c2b6b658b5e2c7a5f903c4f825f34da905855532462d292e0a67dd649125a29141ee4d5734982d32ace4fc6572a3cbc12545ab493e877885e63324b2afac24721d46512d5951657a14a8a22784038647010f44e4063e54eb3f908ef1b1cb747c350ad74bd1a2a876efa587ad37e75ace334982a8d424b1119c534ef625ec85f2673013302b1e0c21fdcd43d4d343141c39d1bd24cab2ce16601263ea99c32848eb901a09978b1ac8a6068794813088046420a4bf91b86bf99436f048c9493013d016a38621aaa4d7e7b9cf925930f46f2136053fc033ee0240b6a6dd94f8aa6039bd170622addf3ba48a1968853f5445e56268fed40d198246bb8911a69ce015cf2f79201c409e452672b0d9e3df75182612b6757da1b985e70d1946a9c81775d7237ff0a39bf5f058b154466fc8fc6041ddfc56b361ddaf07ae0fce34d41998ace5c3d0d7e41ac0f20ed5664aad87930a261081ec0b88f64ba6bb6f79c4a224c5dbb12ea50cc4777d9c9f38aa7da34bd19cb5277f543f64ac113718feea6f25bdcd1dd1513cec94dc22bee92df9e668ef302c3b99c4e5ee172092fee1c875a2c10c6cf97348885cabf6c8da7e9a2a2724fa6bcedfca4d2bd2daaa7c9466b889319f18281b1f0453cdc75cf094905813c98ab3db2427e91afe7f835a95ff1522ab9f392c2660362b84b02692a63c3bc6dc84d38249515f559ba8ea2507fc1ab4b6ec769cf180bcecc3ca8f087973ad6fa3402134d7cb38cfa59a81c5e82f15c15065119d9c1cb5e37d291e248187cd3d820692596afbe065920f610409cfe7be4e8958b8d1635d79d8bb36e95abf3e9961a4c07e73f08e03a3a982c3c337ed6bf5cc109a54a05e0d7762874a9557eb15a854c0775cea6b66fc6463a4b9b422607875746c1c1adb45264da93a345c6b10c4dd9a720fcb3f5d0bc6fb4bb54ba1e2e97b9b87f1d6e59635754e46871fdc16d6639fd3f3ec88cb3a8090ce75a712df647a594f74eff0c1f520aadcba3b31548cf9be732a91d462929714377adc42971f9dca4ec8b2a3771299baed00c46055ce43cbe6c3b80a7532a193b206100432fabe2c11d0f566501529144457d87cf44f54c7f066fd8dbd5a05b1f84d106a00d268fd485d0895e39118d196e4820f36816e88e0e9df179bff303a8eca84e6e8d823bd9ef0b93fbfbe595f081e968b83bca44dc211e75a296f7edf53bebb78ef3070feb2feb067d7c6555d27bb414134b504a78a7847037c2b770b25cad66bf3fa2eae6796051b4267091942a608ed40c27309255d355b7a3c070ec490a87206331cd06ad20c417dc113c414c6630cd04c2e5d4ab654c976bb64fe65fe0ab22440d2016a9501790f7a362fdaefaa1c5b6bf88f3da745ab39b41487a9055d391695ef2b005f6b009b33d8f2e97725548e299d522ac5337eb5e6773daca356ee4f1031ed021b9c6d7735bd399a014e622ffed78e87dccbba4300ed815363bd8f4ed4c609636450e4feec6d202cb88fc2421465b32b5d7e5d6a7c67e1fbfd24b02e121ea5df1d9dfafe3428f3bf6c371f27103d5176c2f612da91e627730e4d2e6637d1a3ed78c7133ea3be6f6225f4e1198d12a8eff638c89dc76c176890b21e8fa8ccc1021816deb3d2670c34c942f16f5080d9f1b326d946ec40ec28ef2aca6b7dceecfdb9895c2b52154b1c14e968b5e21213003fdceb234f716416df66418d419cbcfbde0d914c15ff9c4cd3c5cb8163f7ae0e7d5b5c17795290d9fbfd16ec0e72916b4bc143fe9c51edb1d2a09632d9d45239d3c5d0b0550df38054aa465b47976481fa52d6bb60aeaa8a283465a18a8231f32a4bcc99d3eade06fffad0aabcfda1ebc2c599ff14cab4b7e3c9f943f9ed379476e97c1a7bf6e1bd446cdb9593e806ec14e891c058c9013e34ea568ecdab9f31ba803bd88ef1b84f7a64cd3f9e0ca594815da6f2b81fca0819411a4c01510aa25b57ee6018e32dc1acb3d88adfd976b0f64622b83bd0d3526e0e318c46cea3717e705f0827d2927eea4ad5f0066a2eaee04681e435d88f68c2998e3103d820115809afaf32a19347791ff20d554bb76e3dc37f9d7a2f05a5a53f66f8cbe4af8d901cf3c53dba9b954db43576fb92e6363076278f0a2d849d2f88560a3d3e82d41ede6388aaba4f7910505e75eaca6e1bac8886804885e85efec28273b10f6a744d05e6de79ddb600b3658e811859d2cf09f5825cc473ecf5d035b7fea36594833f26274f5a2ac4f5476b2d2726da79ad110f14420c97ce8915105cb2963660d077430144777cb04322a8af1300773e336f9c6f206af99d3bff718334f9ca9e02d98b31c1e9d1f4a8ac93ed001333d0d6c01a6d152cad2efd8ffe29ec176e57d51682baaaa4980b8f41d4c450da4057cc89fc27ba2ed04a2f461cd25d441940a74ec68f4c8cff385e97aba59843b702894fdcc0e58e4562d482a625ac03d374a9aca25db52d9f7d310eea93f3f078a62e9b30f2e4acfded1a8dba70a62a170321b17241d08ab1a419d74a7d6cc9836d16b529e019c1f15e95e4835845d3f94b5979ef67d851209cefacb8bc3448ca4b44562e1b26a82ec50b2a4a7111b76f9d74339cd7cc0496ff84228674112307683ae05db7770c76cfdb292ea62f38d772f233b3cd0c1b98c8a7aa40e446005a5cb4cb9608562c7e610afd9edf6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc1fdc33618ff0d121fc784e7aacbcc5d68ac57816a789046585f640110e6d121133a316291030503a863ae63e22d2dbd7e4afca244b445cc47c3dd7263b20628a8a70632d1a5cfab0034dba0029e8c8c0791b6b242db7276600e8ea4869a784ddb56cf2900e86dd4847057b71c5241ba2528b1c5e06ffb19d739c70c0f4de0b9b3fb392b4bd873d01a79ce27af427b11bfc70642630d024a8e5c481e21af15d457654a91605fd16af32beeee67f50d36bb28bd7b4695bdf38f30d8bdb52bf2aeebe87dca0ef5f012074f71f320521e0321e4a420c8b713cacd3bd42ff247817e8e39199e3d91b3a37248eae1e426102ec3b2e991bae7f435a47fcdd969134c331556201327c81e29b15336d845929a0e809d4a960216719c1000537377e9f2bec42fbe9fc76f928afcc0ace1d1222136bf03106736dfe39f91a31e224cc5c0b1da1ac7f635b4a93271e5fde70612fc7d97daab7d62249b3263f9396fa2aa0b9be9cbbc8edc84017e7b15f46ab6211f3ee0f24f7790592b7b5eea544b919f7ee070b1cf29f986203376995396d54b074f34ac5c5252bd2901bf7583780fdb480f4fc690c26354295e566abbf1da44eb5582055faf3330558e4ab9e22705dbb0e98486a0f1e583c9aab20f187ac6937f4a5e37ff19c5506eb47c7d1ffe612c577bcb478e4f2ea0ba98287228acd4cb055499523f541723a15132e51a707be7cca69d1a80d07270a55ea9739e5150bd8518c8299f003e837b425b71b48edb91f69715527f916161475e030e2f102213b1cc9f62b5ef4172486ba0a73e5b613a085c2a7b962ce5ef3a3529d8f4ccecbb4d0bdb7a75695ea200dd8bb53ea02c5ed9e892b4ba4cd4232da9ae21aa6bb897979696a00e9229a0a79062f5561eb344f41e3a266ab25ace3efb13f71a24a12c26dee4598a2242c18dfcd2c347a076d34b92803f291f6474ddc6afaf15ef24b9e666b4fbdc387146ca6d0c96f8fe5e63305b36549fd20cf587d14f3f113318d737ca7083a9e36c5c8abd48d364a870638643982cf701a4549174c9a0c5438130c8d190fee639bc270e88963247be47af136c2609b0badf81ad0e1f6b39f91b298813f41b79ab9cc761df38702b1f44c01ed8d0fd711d376072eb62d988552ae9384cb69df1e34119365795b92a31441f2ebe51ccccc6af4f58643df6a46d98cca4ab3908a129a40dfd6cb8ca85eaec175a5f7b6263e4fa2c5e7d47043d782d55b97599d2ac3d02b88350d059a6651344da3370653bf5a9bc9e3592e8b882b5b3a343c14dbca48fb4a6a2bfd200564d629b840b6d695ab83267d5898366982f46d5b84150aa20ba7494cae6be9b8e704cb4a8db1895441fd08da021f1476793036cf75a4b5a37b946afe4af7e5d7488f55e6d0cd68a74fa2609e7a14355a5ae0c64e7018a74a8b00ecd0ebf9e86d9af39d5d5edec6b0bba1058951521ea807be2750898220a0758437c3a5e2e2de1938f6ad5709de99ee2ea4620ea14df16a2dacbba892264d99642deb38c813fedf092f084fb2fe17af232ffafafc3323cf8d2c73e27a6c2fb54405d3b79bfa99e284409fd50e3a8617b549d172ebd92ffe6afde7fee051b2713f026624e61023c3da8b9ac0fb0e1e3666ea95e5313126e39faa4c9d33946b1de64b1403cc465488a0f91f3a3bcb6bedc209e5a1c6c54fffbb0bb83eb326f57934b2144cda07a83f22162884c7e4d8e6b785911b751e7f2926456c377f1d2011b1d320c7f291a6fe98dd465c32df2d8bec722b7aa09bb48af0a591a70d6abd02a56312fc237c538c3baf200b4fc1aadd5fea691ae3228607db89ced8662374910b1791b2d47b2f3f1be2112603ba3cf018a71ca43553ec45a39bcb3693139f6f225ddcefebbe00501168b8932b631059a599d6d2aafccdab902309c30b24342c18b2c180b9ff6a2506936443644fec5078f86acc34d4074661aef84198b2d9048065d021b02e65575c48dc1c03f89dcecaaba21a329692a73e1398f4e603c2ef5d9e97a38e0a15a25f0e7583ce2350905c3646b1aad543a9ea032e68788c8d9c9936115574c58f494df8f19abfd242b19cc4170e90bc6c10171ce99aae3260d33f2eb455bdc1037f58ca8a8a8198bd2c8d3bf12fe0d8ca6ea32593c910e464da820e79220ea72a885942d2a6b6e35e01074352abc495a3550f533f35124001da3ed43bb1c9cfbb7d528d93baedd84223b6a70e4b34bce11cc014c6991ebe3ace8eafceb6154ef8f32cac841517da50f822db9456a293e6653a85613241a1e515fb62f7cfd89b9e2a0fa3df4922a0a523407bdea97ae74aa4d41b567661b5ae7269fce920ff766a12a64724ab228225f2478084763b5e3016892d52a67d1bc41aa08ec8a8c8118385ee678010d60ce4be0a6b7b99cb268f47536c1b1fb8552a11f30a3508145d9a4c680372144ec86aec9b176fc0dd3ae09d321e7cea279da34ec462618330f767556eaae693464db6b7ab1301fb701eeb856f2b99ffb2b2a21b3d4521ce8baa1f2da2257e17552d60a6e3a106aefee1e1c28473962dc1f52409a3161be476dd38df1ed52e1bd5922007ad7158112092c1a57fa43eaeaaad0c1b6e3f1b03c39bd680c53887974fdf795a8c94a94cadab1402be7134dde8ea8dc67b6ec6e55a61b592fc19c457b2ca68a7341de19acdd2390ef5fc8b8decb93ac6bbebc9c2ea62098d1e4df8aba2fe2e94f7c9b840ea736535b9365b3b37c76d49a1fc16a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h64470abb86b75cc32e70fb24d3804fa5223de40f6af64a626b2d4239f4558818ad53b3100afbda4580cc0e517149ad54a2cf5776acd0b545e35541b9adc1bd3424eeae5517a68810bf13627f38a6e83405bd0419c9f803f9b95a8bc0a51f44c12bee06f1db55071d20f8a570ab2240eae43d30a3c30a9cb86ce78b199c5a3e92d490c141233cce096f4af9d5c5d8cfe05bf637a8c92095540b3fc91473a306a9f255ac525d1e72bf1f5c82e22a39a88ad521d03af397dcec77bb17f4d15b59d92101c05aa532b8d76cf77d70ebdd77fa72cb0dfada8696143e362438c0e1a2eafd0ad03289b765b52824667bbfac53e08fa440c4eae3cfc042c2823bc50b3ad1c9e8bd36aaddca1b6071dec5fdcdf28be1c841d8522c84fa5de5ac9e63ab0b0186bff509cddc9cb87f2c7cb32e392c3dd7b0077b26013e7fda5820b5a95b88b6ec113ce6cd713e6b86163a4bb89862b1ae900023f12449093641a57ccac5c9124fb3a18c3bda6c61598f07a13a3637cbd1c08068f16dd0233d8fb76de3fcc852016058ec3cd1c2624df1a19649b84a6c3418afe9eee4e4360a6b4649e8d809a353792b019250c955574d9a87b44ce948e6c6d00e851eaa531f282b53c7ca2c03d9c5842f4bdfa376da16cbd05faa2457e10c332f30996dda68c4f078653bd026044cda71703b887f5f880cef143885173e95303ee46b1cef1203e09c7b0842686608bb84d07df1b3f3b2508458d6810568bc67e8a24869c44c9fe311c0b2dccf0778b4aaa716cd88ccbc63e99e9d6dc5dd5861ed2afab17a6f37141762a3aadefd69ee1a66b9356d15d36a46017dc775673d28db5759b1b10a6f26938be140aafd9c6da851d4eff3bca351680113000d5365c34148f264d048f59908726bdd4bedd3c2a12c8025afe1bc98ecf8f9b524044742e4ccde21125d6c47529dcd16df58b6e4334b9bdd4b366346d79cdfea6c2c8bfa8b72b7c5c7c2da3394906526d8f55d00f53261fb6bfceb0875d5f20696e8f86a4a945b93a7bfb061bffdf3e72a1a981363c69b14a1487dc9e3dc9b9a7d14ce6bdf499f293c70d188d68393d60c22438e34f9d6b532369dcaaaece14d92173d6e028fd724665469a3dd0d160539692115399699a52d7d47098418bf1cf2e833c877ad3fa4558571249383fdd5235eef4a088ebfa1ba46f12e6b0c13c97b7e8c449df4be23880d532c7a12f9fe8a95f2b0888330c5ea3a2310894f8deca5b28ea329cb4ba43955bf1bd41012a2c4831a0d1279775d6f135ac43a7d5520dd915cb73a65867fb91abc2407fb79b685b717a98834bac265460ca807832f8f1fbc5af283b2f1844a270affdf8710e753578b28206994dc6f5da420db8b2907dd128ad802124bd11820bcab62183c8f2d6d3e00349a5a2c91e7ee29da14a6c2b7e1b00d80e0a50e4b5504a820d4ab7d55184935ced38d8c02597d7801ce96d20175c57853ce819aecdb29bab1d7e578e689a136231635323246e51d90f20ed4a7517d8ad158e1fa3aba209cfa9fa848b9e3e9f8a6ce77a7c98f0b62e95d67f7461db527cf4bd8b2a79bc5cfbbc3da94747d3d6f7a69f30c5070d70e64bcb78588fe2c8ca442d41e5f10a17e463410c53f3e696015a2aac860b3c68ddffa518e8024bc6f9321cacb53ecc452329c2274c9042bf37a7f6e5653c695249b3a4ebb2f9d19a9dbdf71452c224b4a6d2b461733d4f1047dd834d48b2d8c4daefb374ab14d95c6e0062dd51009854aafc45cbabd75b2811a46114c9165ba607515b05dfae960166240d543ebe61cee16fb295169a459234037031fd6714d48d9fae4938d74e97589be0bd65d6d2ec174c39fd2325d367560ce13db4e9bb84de67a3ac559c69f8c4c1b649f89280a47829a58603b42af436c68f8d07b47a6a6309d837497160df6357d0801ad0e209bce5abec26fe8a89f5926732f8328c91897c1390a5dcfa06d98f512a1ada2f03414fa5f36cb029898c6c44905f29e8704d9f25a280cc5713a74e9ec601a1c9575da2a91506b3a148fcbea6380c1bb718c6f60eedb9e16783dcbcb714ab54c06656606e2a343f80f5c5b266481fbd8b0fcac7b31f0a9b64b3030563c375ced30afc5b1d171fa51d484dd0d66c6833bfbd30619b2d12d1dfd6092bc4d2fcf56294d58d52bb364d75bc15fa9067d4156c851dbb63baf33db61cd3714a3f559d4c75015d02a19f2a186dd0fef51c2a10d5048b12837d31bfbc154336eb0bc70eb260f76eb6471ce6b594919496fdaeb0447201afb3813ec5dc12780ee2861e97b44f51e8f85a46e501906a3b53ed486ab707f34ef925168c6bd24df1e4271d3940f895965c4bdfc7a80f6a07037e9f752d391a2194bd81fec2435d3f3be9de3cfc2bd04e04e7bca3d335cf57371d84770062e9b8dc05ad53ffb0e4809231eacdc891791b426740c3fabc7046b880106801b843cde6f93cb1d16e27ec6b96aa3a7e6980785b7932aa47770fbca4f68b76f0f85afbdbce7fbac0a3b2879000df8862831b7c656110d0a09aa26bea52e2309d9daa4b86ae7df1452906bdd385aaad94452fe68fe910f4554773c2fc6b343ecfd6ff39041c77e9b1caacdc5c4a33dda846f57a8847caeec0b792101d4c508419eccd549055f20ba1e679eb7047fe82c0ba68440d4fc12a015ffc211b86ba353a5aa2c59c0a31f6d3d6413d783f69258ad33d2c0271acf1349d710d144d37869111843e728989c86efabc5ac977193;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3608b96e2e94ad79865d4c2467b515917be8925eb335b42cf03e87574b95e6a6b5a87a24192072907b73365e7e53f35c745381256282fa94a19124e09b999da390cfa82b6585e2f287c73e93655eb2150291673b351d8b5707a74e5b4b5a9aabaa839f23b243440baa161ccd1ad9ce0c213c73b4490471bd7ef5b89f8a39a4617b5f6789cd2ad7cacf866d05e1a7fe1e6cd96a447fbd8e89d2a0639886424140d517ef07e2de10652c81fe1522f48f40ff577c2ddff0094c11145af8c619c2d302b3bee940e355554430ed0ac9e05a355b3fa1673d2dc68a5d35e7af261fbb45e1e80ce2bc376084cea0ce50a3893d10ed896a5f94a6ea3e25665ae36b70ffd515651a41467d4372b0cd07599437a9893ff0b19d6cdbdbfde9c922c9d461f2da8d11aa7f7a4501b96fed0b625bdebbf682dff3cfe3a17ba617bd8a1efd5dcb8a3ac5b812d4c921d0f56ff5cec7b78199c974f3fc5b81345fec71314bfde1a272dd99a72d95d5e9f1cae2408ff462b1527ea81e36e8e1bde2fd1c08f889ca885eb1378fc7c21a7f9768b5ff33a6ccad476e86981d6826a04751cdc0f53bbf3f0330280155e8621c72a98ec9030708d4c39364ff3edffab2a08bf3d68c9e7b7d8cdf47332a44cd0da61459c4ba2f7f6198cb4cc8e833c3d5afb31a1c9ccee9b6ff3a1d1dee742b6f0536bb5af17ea8c8710aa020e89334cdb0b670f5ae67b291609f26159398763adf292975d8e4779172db10a9723a46ff7a25410f4ce3624f22a50e39bbc57defde6feb97c30140c315f6e6ece5a5d45dc6bdb7c473978da2ed7ead2bb7f55cf45f094d08173a8ec6659a928f95c0e50add02dd6e8a0e90b87fe835c3b914b51ffb3978bad9e5fa5fa1f19301db625340788a6fa66e193b9d6c3ebca715f8f85b20da26e972aa6b23a8f4b626c6d113b0bc92ef8f48e69aea909aa630f2c2848d662123c554bb86fed16e72dace97537a613fe6895973b8c790f0ec99cd45f2ba67ecddbe88504b7acb962f88739bcf770454773a5015a25bba47ed26805f2deaf797ed142d9b729b94c742c5dc9ba2b4be6886022fd3bb0b1c396d7ccc797be43ee4b0cb4ff232a2601bdc8b05fdd083fc58fe2b23fb5c9014760a53587ada195507e37f0a6ef4cfe367a299660dfd86d340a6683bd0f72e517c2d0222e04c6db555b4cc050fecb1299e611ecc0d14fc58cc978e56ff39566c6ad15d5026241317aff234643a60db0db912c40f61984ec72e070c31b75b45abd6dfcd82c39701e42a5c7a8f87b6759feef8e0a942df536a763cd267b9c0d66f1b4c9516616f6e8baaed5e1d26cf0cce542978472c3b921bc5c3c3fc0ebcc3d2f312a534043e06a15954783b06ce0b24a4d60ee426b622594141dcc751151ad41d1408bd88c965d6732820adc0865f60274dd6978930d4446b20a3eadb93d060c3557cb5b9d8eda587164be5ca12af695b67cc0c15f8e0478854fe775d2e05ad106f2236ebcb71918dcb194662c7bc45e5552460d0a00805ccad98e7ff2104f6e4a2c7272856b28cd26d87ea5b858335eb1788f1e8dc9c2b4b3a855fe4c110727581558817d951c69e0e7b1467600ea8f657dc024c2e390699d3c5288ecaa7a88122a8b566cc7dfde8daf64031fcc4932a3c2b509b0c93f0848552b5127c8a8f98159e3134da5c3bfb81b3e31b06ebe9dbf0a4b104fda8588ff0f64c0ec1be4466d499df5d762843ccdd09b552b1234004f451cc0959c01024d959a7931188d5c2ace95d06ee9439abf3e2a6addb06e2c3bc6032c9b6a5a6c8528617cc3bb6d2a19331a73cad505fa125f5bda1da39b94a818785b46f65242d392d6fdfae2df84b37a8dbfe9c090fd91f9648de10908630ec479582ed493f45e3945aa7b2c236e3e6f892ec5a4eee6a583dec971a55782e68b80022203ddbf154c6d856a9221f572491f82747e344588c445c20f8609f813912b16f67185ffa275ed279cd0f13feb8e8a11e311438bf5fee8c4bc5f9f984d07ce39c9a47728c0b29a37ba5344a60ae8fd1d309798ce6a3a13a98d9fc6fe7d4bdafe42f7a98a6c9fda4a378df5b2b1d384b0b316313ab645eebf3090d8b530d52149b2e9a012f91e0e4cb2c58278fe914c68f79c60b3b93ef1b86c095f0c151e24e2aacff25c369d5cebd102578302bad512995612090d8a0848b882fbfe752ae630fd534b43f89dbc323b1e3ee4da48b72685e6aac42141e079295209e94f9b4088c3af7f190f7d738b7e9eb4b6be8a038288041b72b990a7c2c31aca215c983af03811978c8e4eaa36072ebe1e9ef829fdc863e40c7f41b279736c4462afcbad0b5cd02dd516fad725cd7eea1ef7916964e0bd6a310e083a93f2ae2d55c1d0c7024930100c8c117e471777eb14d180699d628a6f98fe71cdafcce84d1a20c0e3f7d357ee1ecd841ba562e66a49d215a75d7d1701ed7a8074670a6e7e3491a115886ddb50eede874d520ac2784e0239ba368d7bef6f76bf88b616780f07d7b7ad0bb26ec9addbf6af7b50d121ae6d967990b8c7439db0632092cae7d3abf17ecd519bd6296040588381aea6fc81f4a2c2a4677bd617549002e263f7c45e13f190d34912cde5dbdaa0ef3cfc7ee0933d53bc069045898272f055fb629836a9d4f7830281f3a05652ea90cff53ee1cc8d330c3a34d024ffe2bcb914766c8ef95275dc71658c082d8e5b03abcc686da7b0a2a629888b098f006be3dcb10886b4f8e076d31ee01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h10a58cfdcfdae45bc8ec38b2c16e7bfb38d89246367b450e2e62c00cba185061e4ad4cb034c2158416f3854a2ac8772e2a4d7a6b1b932a989a72fb66f9e38ba9c3092250e5e45e9321727544ff611c6a8ccae7fe350700e0fa264a233941a9dfeb3887b2d4e9fd84acb3843feaa206c3fbc4f0e3b606fc5a3d99f93c18bf0454b267c0f91b183812bde588ddabf0bb953390dba909c7d4e722f64e4e712d33e1836894fc2e4ebbbe4262d6dac84b24387be9a939f62db1f3c7649cb2fcb5dce4ef7057e1fbfeb5c7800c1de55546650a1faa4e64c213cd14d1383509cb6f4cd1157cf7afd3dd943f81b98416cdc994a6a9e4858576b09275a703f18200a7c2b21ff062c625e9154bcd8e8dccdece0abe9271d37b7aa117d22927ac9a2d222d51c0d7bb549310f9dab654f7efeea4cd62cf61f6d14f2bd3e954719e3d14fb113af861d3abc58274adb5d3563c5ef3dbb5bc1be942a273efbadc381efa352446b1880c5ed33d1bb3df17700d2c359b6efb27a6a9201940ca3f1a89e8764dd51ff7b82819c4a529791b59c9ee7811d37610e0f73ed84eb147355f5050b1dd22b70b46f9357a1e5bce9c6da46f6eb07e02bcf7d26b7515b80124516572e9ecfef3952a61f5fc2674c790b50e4b90bc245636f0567e97ccc9ef844acdbcdf33a631745edd12b9398481208d75592f9ed1c288d3a8d36218b5072a2a85c5c282525aa01e50e7f56df2da42dc2051c5e168521c67ecf336aaf8dec32b5211f3087c29101916a0ec30e5accc3d1c0aefbedf1c449763cc61ee385db230ce1d7c89f4df216ee5b1ec0836aaeb9cabf96ae28f845d7eb049685d451b1a509afe1d6ffe649f6afbcc2b0a2ba58ebc9c964fc5e8271f298be3fd77eee50c3e2cfc2728b2969ba3f12c51ddda6c4f33d466bd705060fef6b8200cf1c7568b419b09e9355c553d24bf3591d0d64ba7491555762386a02d96127d4b61b7e014a06eda3778fc507b7a79a99d54868ae2803389145bccbfa6311294247f2d810ff54fbe1f9b465b5371f9e4ef4a22e9ffb45544593f421c43b51c14b9a8f09fbebffe07a6c55df3dba47247ddae5d6d6694a529ae7872f2ead08641ca0e54042dbd6354a8e969d5603ab9c7495660491d1262c38f3d6f35a9c647af02eacb2e8ce68bbb3d79782ce032076d12d541e23d71acaee0d5aa0f1fa4356fb625a4040f45dcb5d27b17a3876aafd1c2a595c2dbd1c9ddbc514821177eec665ea09c8b33e5480dbd4d363501f8cc262220226bafd5604367640970e3797e26f29738105229ef5139518160f7457aba1ef1d992a457b7e90d11f6eee82d5e3767c85626c1bd4c072c0aba4a8e45454c16ea84a84cf07255a9591c950f33c1d3f18f18d014e2f6e8e9f47bff842212451a4e036d592ca9fcfd6b38df6f7b57742d90e16d5fc851c66686e26fd63d8cf58d52206bebdb0f10a3cd7f359b7686f91fe55ce834e187cd10d4c2031d31d13878fa9513068e19e95ad84bad4f08de561eacdeb723f0d08932c7602ce7fca09322a65bb752bf82d7c0f8dab576d3c8d91dac8ffbaeee5d45688d2dc48a432fb1f05c27ce80134499a22c20903a28da4fce591e2687ac4bfab070c35cfc3cd52be174fb9ef23b4b8be8ac135dd34af380f5a30ec0dcdf56a03e8ee660d0584eb4bf2f3d40dc18dab4191ddb6ac3d05faa5a5b232d4f2e0690a3f15e30f4308ed6ce54c43c69860de9d637203a89c7e75cfbb803ebcd0949349830788fbf5087f0178018336312991369915b5c9589dfb36732dded02e9946f41c9224f837a05f3094c95e20567cd99f76610e3a1823affb7d3d65f2c78299390fce0fe3b3f13f297623087af7ace16c700e614051622739c06555b2573fe32d77882da40f25c502762929d9feccda5d899dda2ef5e3103734fc952d2a8e514e64fcbefd21369a36828a8651eec7901887165a767e7a356c92afb989539cc29b0668c0601fd652082a6d590674da38ce68ef6798acf4afad4c342c607919ea15bddc6eb2f8eb3e087ba179144a33c0696f5a4c507ed40c3a9a116881590977d75294d37f07cecfa40a3df3630cade0bca1a0730a0fd51e4e36bc43a7311ac3a6404d937b074c1253dc159ab8a07e8ed5ecc7269fe0583508a030ec210fa8aa0f808f0ae8ca98331876fdce1d871aac3d59b4b262ca23e3a706b6ed6d23cfe9808c07155d8f9552c957067034e2bb424347722ac8a03aa2577999609de05789e2d75cba4cc15f5d8ee5ea19cc53e42b39c3360aaa0f22989089b347f781a0989541ef1a2f261369daccb9ecb6aba5931b3204df9ead2fce83bcac0c806f8d9a1cb8afa6ddb4f9ffaf39fe561b9ac54c050b3994fe535b4ad81084c2a1a7f12e033c70cdd36cb9e35d413ed20539c76c94a01a2917a11e91e03ea9d67c40190fa007e27bc572510a65a0132fed5ee01dfa4a236f20f1875217a3f387cf39ce4215c31c4ce75b3e6c1dcd09cc126826e98205a0502e62627d3a4e28a45019998a6a701fb02b0ba44a8af8c704faa54117b900ad8f893496a5393f7e7a30fd8dc53f3ae6790d000d3d0a10261611806b39af0b252eadb93346f30f7c622c133f5dbc589a5a8f2141b7f37a92162fe6e0f5fd545234fd8e3b2d8e24c6ed791b2cb3093e882dde5c8980ffad5e887ed90633bd5256c35e1eeca8189e291a1aa86eb97f5d0ac8d81e01b9a813b2aeda1d0d71a135a2884a944648faeee7f3a3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5296163c72c669f846bf7bfb825882ebee2ef2eadafe7dc338e1e2c5e2467cdd0f720d1cc363b59dc742f1a5a54df27ccc8fb6973872d80f70d3f20a1d5789567c95587d676fd964f8b02a4fd335a15fd519e6546d31c31705a8883f3d97a67b8e62ec4fe6f481e104e08659dba1191e3404d8e6cb44ae5e92f7ada19ce6b8edc3d892d93ef2d5389f8b70018c7c71e0e65e2407e5b116820a76e5459ad0e594ab8e344a8cd6008c55f16d41d5c5e45008273e79b29baad2e4a551e9144c186ad28fade375ff9ba5b2559f065d17068d13819f91f3afb5e2d14a88974207733e9459e788a230204c44afe9f48e99db291c2e407d7bfaec1db1d4073c45047a580ce252c091d1430bb94059903466f99faf0df14a2cb906da445ffecc320d77fba6d475a0c7f76d07767f4e6ce04f3c7e86daa92945a51e4809734542dccc24ce3352b822e17c27aafde3d179b9ab72b4af342e6a7c4da65d9a580bdefde200cbac00b00038736ac6a4a00aac5335df0277dde63a461c5bbe42d545dbde0a07f4178ae579164df1430270a519e655157e2a549c3791a1078ee1e5214e500cb0b7a4a8609a9cfd1b0745536973827c04fcf41daed39a6f0dba4ea59af9f6fd96942df171dfc4cbd9b336769382388d7552b7faf90cca6c6a1adf9f03911452acd0f0f57cef0fabdeebba96d3d9bea6c7151e0693a5f22271845cb400447a8e0b1004bf5e459c8d844d8f6e66fcb36f4578cfc8780661b56d1507b9b9ce40aa5e8afb96779c11d946aa1480f2fdce06307a6d0e1b08d6ba484eebada8f39a2e4e14e286df03f87405b6f4da2a61133e3563aa19372f2e8eeb4540fc7cb2c1277b5aedc53ee0c912c1f96dd2c11f8810ae30d9a479092839d70b8262077a70865dbcf8e54ba668a8849eefe56a569dda8d0cdb39a07b0d7f0c43e86b2d69392ddf75f0213fdb4169834064f2128eb042fcdc7bb9a4002538cf7a17ea23641e0f37f49c8a0a318802e3313ca2972c4516d76cf8222b0a3fd69827c06ae64da7889e7e92c07f866f99b84c42c6c3ddff5d40602391d8f86ef22b07a548617f1a82b98256be1426ed729863890d5404c384a67da292c8987dd0139eb13f67a4b36873bd17b2c293d7f156118aa1646f33cc1cf1f8b97e8f260ecafd5a812eb3ba1cb3b7d0ac945a1a1001c044f5e1fa4a378bb82761375526265d1f3c2f4bccd7ebfb497ad85c82eabd4f99bc4484ed51f14eea67a3cfa3cf7c4f91416e1ac3bb0d2d9f1482955d8fc6d7d2f6ad8e24b7bb45f1106915e98da49fbc7f3daa5069b9038ad1a8c735ecac9e34d126e914d751dc8c8da29bf4d1f69c3a43dc3ccb8c745d81dfbefaa680fc3520ffe5507cec27be993bbc6dbff47f00532b9081c14a48c6fbc2c274854d0bc79a7fdcc4720914c5d2a008b9da944620414ab6494df4e3c916f40dd616d32ca30c42ac8556ab7a177e956e7ad5586c329c13715abb67ee75a30cb4b47778a57bf1a461fded1820eb450234e0be25d23eb5321dcac2d9849b68f74f5c031bd9e4ad6da186e24eb19ab567343cb0513bd8543bc39d47ca4ebef10a33ac236d47ad938f3443e57b5097f956649a51d8295f537b382e7eeeb7d18c968c3993354db88f26352f0fa373362a28f237c5b7c049924d216e423c44818d6cc171be2a140cf9df4438e304f7ea4a999ddc330ee6437b620ad2a75682d8ebaca9291d2aec7e5eb6139e6c23ff6a54127e3704a05b2e40cfacfa182cf502d4347ea1bb1e50c895c591b9911147185bb5a9eed3f7f65cd6aa4c41f6179a9df0fc0f3a2ce3d261674d580214cf7ee4fed534c38cb067c1b49ceb5b1b9bd9bd9a9ce34272962d84ebbf469757a17172f728f4128c5308c581bdbebfa40ae86194e9d68b1ac77155de9bcf13d423a668c6215c745b61cc515d56398b84f4cc9f630574097cc1b62a985b1041508da8158a0ea70e4f2b29d0fdd1496dd6e11a174f8a281f3a2ae53285590f2ce2139d7cf17574dd809cc60cdf673573ee829162d9daa5f96b2bc8aedcc9ecc0eb28a766740fb2fae008d46fd14483ac8089f5e23a3ebbca3bfa6232d380983cfdc0fef313d4fc9e397b29ee14d341c0369dff4ab7ddc98f8df6d49001ddd9396918aeec72ca8db519399b98f1410852869a16188f54b36072344bb45f7520487bf145610b27fd3fe24880c53f4ae8b1355cbb1bf1bd2f540a044a3130b18981e5c2378cbb882819e1a573a195b90640f4c7b432bf3a51c4907372a868a6af5482dd90b2127bb8d397be87ca2ae46f64fa64d842fa979a784073d1ddeef95ecf7e85c2fc591a4feef5c3e5354e51506b941be7a3c3031582a3ced18124e24a43145321fe9725c23716ee684c2882b814da58b9e7a8e7e5ae3e1053638ec47e3c0c566f491e6fd251e03db677e0ba8df62094db7d8dbc64772f55707911b9545a4b68bdf5b49c8d3c236d5f1caa5ee2293d3b9c4ac6aa0ffeb55f73f6372ab893057c122d47fefc4c324576b77928238f9219dd46a77de0886c94d834ff606ffaeffbf9652a54ec1fd0251855a4124663a76c88933e6cfd5587460f512e0e2a30b0596e6824ba13cbaff7829535ff9740afe7c0045a11c8aed61016f44bbfd7ed760184c0a63b9514b36f4551a8da412fb4accc8a7ffe445358d705ffc68d4255f06aeb6e8feff819dc885e8fba527527a85e38bf360c53a9dec15dd3a5bf5a0666e47471b7e66319e126ee1567;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h639940d8937b7fdc9de1aad54111d1fdf46d0917f1c57bb886146b4b780daff0ed9218428d320a8e326703dabfa1ab027673d52dd4b9064c8cf214d4b1fafbadd4845a67caa4131635a4f9f610ed7b026d9cc0ac4d1870838c8b99b1339288ae28d6e6cdeda96df93488f1aecbe334e6f4f947d1c0433bf8579675520713915bdd8985c79d601120becb5deca8361c22da7d47dad3a60ad617ff3b6360c01816a736808effd3fb55e9931c26070dffc51026220128e9ce258aa8ddbfaa1d3fbc084ad0aa27df0f31d35365d4d28141ef7c77645b169aff82fb606299c49bc318ea0c4df7d8b1f1d96ddaa0da34c6649f8a8019b5308919d94400cda20475db0b6672eefcdb56f1eaa75c3b56bc68f1a8f7baeac551d4d49d8ec409e7fe00c5198ac8f0e5a9e19d3f947230f90d0c7b14cac19911ca7e0bfa29e32e3a4290f6b3d1b8f9260670645fc40836d0384737e2cf8ef388c4bb46b0821af05b8644408f5de633c718415d8ad563bec7c7ec4c2a9a58f86dcc7e6c60b15cb20e5b62c557225186f71c7ee4298ba903c2b35b0791dbfcfa9496c48f5969f672398f5cf300f5294a9a679176380db0d8a4d8810e7be2cd921541c6328327dad7837ab4d729b7a661bbc90c4a1f344e96462c9a7e0f9e1d743526c67bf7a6867593a60296dbbc7715fccd9deba02892b67b7a8c2f7c5c1ad53307028f6a0d10072df1cf6f14001f7920380304a4b94b0cda123c0f20118d0c54a2ce2b6c452fd062128d76f9c435a7396d7beec375cc0be842ed0f314bf0cd05788c67e99e6556d9c8f770ee6bd9fc55d05c914e38a1f926589c16385d622411b386be2a111ba8f8755e8f5ceb1c36bc33cbe0f1cf76d04be84c65182a81c990a701f4c69f1c704fde2febd7c0745ede4b82605f97a33f00034433324d994c17ba8da4310abe6292fffffb2643f24923fb27fb05821adab8a73130c27f5bb6a69ce886032cae4e8261441fe66ee64cdb0efb01529d897f45e2031586f1b531af163d74ff93605d0ea9aa366200d71c4d006496bf0f14565f01e0a5a3fb14239d801bc5e0085291d3f07837644cf4c7782b77145f797baf2c6d4f12a0224f66e65ec233039e668e7834805bec178e0a62593453124a5467e3128eb8416c1acdd6c2251322996582a5d66faf038c769e94f3caa8f86fb2e0e82489e10229049bcea29fa1d75a75a401aa4c24c6b5d351678d32ce763925869c55436927035d8c60173affa600377ec21a4a96bd8a77f70510c718e2b3c1b7c54b09500c2c2297c21c9263407e07699a1ed9fad96028663b441efe652ecd3fa199274a0bfe7ab975e48de22bd8501b36cfbb429ff96cb9cf81d8fcabbabf71487bc4e1c54c39ea9b07ff84a0b9dc1b25795ffe9e61af23bbb8e0f31837cfb4109081e819b5a169145a663b2db9f031600559740dccda88a7a6793db023b2567a71771263e308ba1c8ff11e28529e589f161f2832890b429858e8d35026bfda268d5d2f428cc468b2cefe932763f7084e2d925499f0b76a49389caa8fa5ff937e787534ac18411840d12853af55583930bd46ba1fb77ae310eb2e8cdb285e2d381e30929cea03761884f2f551326f68031ac1d58c0f4f574aa3c7854dfa4d3388ce91c332ae1787bfa4e689b6694304d3af09f2202c473de5fbd799cc05c0663b517006369b72d4fbbf901b431a821b27f46706f5e9c22d9e30dbea989a2aac8197ab325fbe1d71fa9803a76539ef4a545f087f7fb44b178bd7028e7eb6637f73b728b408bc0092a4d805224052e281953cfff0d3c5c0ef713396afd8635ba7e117a7cd0488fd80d5b0499657c080a7f9a679670f62177dd3120c0f86a74a2318b0f79c503829eff188e9e0cd776740aaa3d5b746a424b5d2457e18cc16ed09bd0b28b47fd104831e8cbc5415520a7b9e9469435cfc66ee06fd9a6be22f84774048bba234cf6776daadc106002bc37a1f2233cfc28741068ca6fcdbdc0f8eab675f5f8081b125317ef84729cdd1193adb72cc139ad225a9bffdf6a13f87f00faf7e3c710837365e3bcb73b6fba4c3fdf5511206080da08e9469e19cddaeeeb78b6186b352ee2e689b5e045560cc965b82f4f533c6fb73bad5a028a510fef1b4006a908f9006ed38d9e0a694f85b04642148706c37dfef6358795e560a483ffaab37b3ddea2bc903a4bafca21176dd70afd7a824e2196b096f3779267517a41f653acee259dc274f416593da9488a41f8f9886c19fa07fcda6bef08f9ea436846a6febc04192fc1d210317b834b3b1b3e415ee5aa547db9697f025f810272546ec66ee24fbf271da806e1a317f62526ad8ef6910f0b8a6f7418089297ac92df67c1ba60fe5d09aac4d5c77fa6fd3f9f9e997decbf0ebd6d2a8d67cef0ef49876626f214fd446c79cd6d4abaeb2335dfba633796f999e113cde45e5ac28d2d8c9a6bc82e8ec7553ebccd7474fb03169ebe4ac537c256a151e8235721432ca0dbe051ce5ac798bd352ba7b3df80f9ad22fc596d829fbbf2135b0c144754ed225bf9e5c354f7f60c8e2d37f24b793558f42609a2e463f1e1fec482533a993c1398190338221cb7815a8e2f6d12f5feed83db6421594f78db6e06d90eb0c1602bd30086daea436225e7efe08386f75a1c3d8de462e9e43b7f64a26dae196d8e45e6e82d901d679aeae559eb62946ca786266eefa7a3fdb20e760302ea73ae70a8fcb74b3aab7328184a736f8c8c996;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7e5595c679eb6b10e4984c5920c88c01d9551a5e45ed0c22fd463b721b6c5821b4690d798980a24c7670bbc1b5116943ec3fc27af3303276141b1e269088e536d5828156b225f9118e981899438426ed01ec0d73666dd3dec138662176c42973ca978b4119349727a9c5e0358fbdd43abdea011898a596ae0c54ef99a79dd2d8ed4f96ea3864be2237daaa4c1ad6ed154efe67fe454de4a56f9b6d7e9960173746b9deaa9d8bfbaeefedbf9045c7e8cd0476ebf752f3e526b0450809b72e56dc42f3d346abc9f0466bb3645f862e62d209058ba4e39043d15f9bbf29f6694524da5c61a328e3eb6642cc24e53ccfafd2916206e0a849b814993a8794536fb8c0ba3228d50f9f4d136dce94a4b500b3c7ecbc911ed1432d5d1dad550343ceeff558749a0a116845f69d7a8cff273bfb31ec28114ec645aa1b619e8c98851ee827e536dd0ee594c61ac14babf35d1968bd9a26991fa80559e4879f9389e4454d5ed2b289623ab75d4263ced13859b8dd9934e0f3411b9ffe0d34e6b77fc8a81a883a31bad27160ab9caa91856704bd938173f405c34d5f489500b70db03407be707a2d9db32feba59df0ea50b155a9f482caa017fc5fe32567e3511eb52c7bd99b2ac49fbd354f55486b28fce4e81e66433e0f3e7b70e09f7c2f3e7b4a2d03e3a0afa91233e2cc80ab0cc237de5103e18ae388e72c7fbc6be10dc7f5eac65c48b0e7c40c6be292a7db2e65d2211c7acf5e64a0c785caa3a6c26b73bed29ff52ca0c1addc3201dc3319e1e5e637dc79b28d280772277a46de331af25b6674b782d23ff5ae4151e0d56ff7d3add74fdc0cadfcd89f5bee5f48339a10a1cad54ab6ec46da81ad4f1d58bb21f60b94eac1366cfce1251355f0d4414f32838555e876c7dad3b208f5f2102c6eb615ea899799046ab75e0cbf3a774f223663976406c46167e6527e4891a2ff809b5c74fbfff87e44775edfcd5839ae02a3d15eb96494d1e13f1a3731388370894bc1ca24a37d390aaa50e0e918cec780281994d4e9b66891a0fbc25dc1740166e7b0bb2d65324e93590205ada216e1e73225af2967825e92f0ce3529afee8e046fa5696b488e6d230afcfa3aee7bfc1b8ec3ee1af2100d16db1dacbf71965524e1f5f93cdc4bf05c0bf2a2de28c7349d0cc1ddcd3de51eb73cc257e46a0f93d94fe1bfd8671fd5f00257d7a917d7aa5d5d8f3cc7d953050f9e82582e0d23b2a93f2a92fbcebdf6be9d77b1f3a936d14580cee402d9b380d77893d7d6c4170e9fb83cb469f3be03fb1972caa15b7c7a186d42eb067e64939aa7cf50586815c5288d70e6ba6dfecb201cfa59f3ab9376a62d7aba42d6841acbbd42fda738650f812929e823b8ef09be326e0f8424ad7e3cd4ec41d23c1e690b5a35885a8bf8b44cd2d4b539eb7d22a1b247e2a48a84580eb41b2afd0cdaa8d50d4218ec9235ba663fc324dcf66fe38b878b63d614c605eb9dfcb13644c8b3df4c87ac89a4f682fc786b861a7ed4460ca71d96e3d6c18aa0aec86a15e656bd596d18f490cc76a3c1a1ea03b099b204929d89f8356a050a851e0dca1eb6f4e9363c9fde08abb28886c3241f8a8055a0e518c281250625a6d51d52b376858abe2680f0b9fbb368bfa2c4848ed01a1bdc5beb37538f66680062ddc7d70c17a0aab3847cd499dfd1ec444de656575ca6a85dffd35fdc596ad5f12c05342cc37978b6e138d5b971ccde21d27ddb8249a1499af1ed8116d2080afedbb75ca9d2cb8a499617b38740c171bef8ed2ef575261dae54b16927e77287dbdfe240ea8e2a60fd80028f6bc6479580e4d9bcd3cd1f45979a7e1b4769b077b450c464b1693f582794b309bb18a31b81777e6e85a98223087725b30c86dc1e131c5758f37064915e03b7cd59f1871135d574064f466c854443f18090fb9082b4d5b19eb853fb8f67a082ef5cca6103a185451026112c74ed25c95fd7addc4dfd908218334b411284f384a2ce8e5e56d192d0aa26e906e243998f8a932f100683e56358679cead2f07e157e24494df285f2644579257883ed73839605dd1ee0a3636adaa016f42bf2251a7f4d4ec10c16389b1a34d6a53cf7f55974436e44fb9e5adc772559a9c4c8e4b8545b461ded57d92aedcfae95b1ce86efd5012b8dd985ea81bc9c5af15801d82cecf928db3e195953160716a87a4c8eea88934f5a398cad60021f823bafed544719536d3fb39e716c02fe76380e2689b03f61bdae1bf42da7c8856ac42db404e8159b63423b19d193617e555ce74ccfafc157f90aa4833372a320540ce417c925f90ba8065fc2dffe9f3225d8668902c70eb5c37051c951a55bec14bf467ed6a4bb6330f67a4d69839ae803bd4bce8960bafbc650aeb6dc26b7b6705cbce1a9b86117a63def28a1b9934e6551a2722b55ebdb72b2134798f1a6d8a8e317c55af42f7db87667c33a368fbf9047d6247a1ac69533cb521e3d61dc9e2060b1202c6b3ab6435a26b2645a224794d0cdfe6da753477474503a1aae8c57f471d4d4e1c46a1e4f4d20896a991f049c21f3c1ae8bc3e7778ed1377dca83c52c7c576217bd275b76ceb6c339d11ac665b1590c98769a3ab1bb245ef2f2aa9843cae2d40ec973ff938faedb118dd7a19971fec21489ccd031f332a91750573aceb39e480b1586d0358e1f7076eb2a4badf2416343f6b34bf3c1b328e34802e34393cedd6f66a07c515f26d9578633c32b90d152e7b6fd2131a28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6135542403e309701a5514dee787b8a062a451c4bb75c47c9ca19d0003fd4052bfd0918aaa75a701bc15b07785aab5c90cc8f44b381e84b29a56b175e8b7e4b27ac949deae8a81bbff21fce7bd977a9a0e47b38636a10e7d54f3fbd6d5d83467c05323c47a42b36c7f0a403b1011db58ef713af1e4b6a67fc14347f17cf1bc5098ac4b400288bd4daf7d9a58249ba6daa75c6c017c8d4355e71b62b28d65f42780766fb34aa3a5790e491e3f1f9f4c38f3ecb2ce62373dbeec197a84620700989333bb87a53be3b5e76315a0a7e7d233027ffde2d0157ae15557af273c3aa9ae9e9913cda4550af44d2be5c447937234d3ec0beeee19d7cabee2a81153c63c58cf7e4e3d344888874dd742ffa4b7aa72f58dc354dcb90ac47ced5658a489c08b41b2848ecae1d16b8df9cdf4705ffd2442d45dc9d387e7f908ff1e519d1ac0a5ab089537497f702774f3f4fd9c3c74b5277c0982d16a91d6551cc9d46f4534dec9e757cdc590fc9f6dcc8a0df83b459b16b167eac0a5f6c72609d34fd4254d3bb42b170bce520e8b9072d4c046cf5de4984568c58b2985769e3efec4b760e1436c5e32e29b8d9ac7a0965c0b525f9b02b69c25edca74c7a6c4f62fce7f06c520580ccaa3067bd5502aeb2aebc7647d217e543a0e1dcf1f6e55e70442ede893b954f7ce8ab3639122f6e07c85192eb1ec7239d04de824923a10a606e71a0526b186df0cb2b1a06bcf8d54e2ba58a43b9542fdcd71d65ab5929b2ad3a592116f4dc1383be39ac663c35d1ef5084a1bf1ef8f6afbbe4a6117daf3b238207a32c44feaebc4335b3d459a76a5e50bed02ba097a72be18dcb32f1dd1ad5c9e6de5d597abfeef155a2e00cb78e66e3b728993bd2aa625a41147030455f113351daa9ec6d750bd85f582f04e7f6fe194b0276a37901dd9a0941aff2933545e61934943ab0859201eaf56baf1ca464de86f3db19ea1dc48d0d69a5360551a0e6c46e5dae1bd314c30ba5b1b47686cfb7b488c7f65d097b5bd23def7a154cfb948e9446e71ffb12f2b4ec4855750a39e7bb65b27cc71d25e430f5b89acf0ce57c8c3432d2763e4d1e377b0a593c799a8721ca366d70c2f2b8fe4a1957ad8477b2cc7f2d464103532bc0d7917dd1dd3a7418efe687aa11b7a270c6c0283decc783f856ba768d5bed7eb6198185e49e7096aa996b31dd7077c183ea70676c330d3a72c764e26ed40f0eca02372f07a0173f9427d78e8b1460cbffcf7d3aa49cb4bf6233525c24ba7dc19668be35734221d98503cf30d5b0d6219f3f16b4587d856db511bc9231ef7d5990b4eac1c39327697eceb08896464b4cd0a748aa787cb06ebbb45072b801a0baece8b3b78ea6988d892520a71a230aa470b66bf20c0e074e14458d950bdda886ae70100a86f8b7f2ec24a54ee4adffe2882deee3c1eafc9e51ffca47722df3d21057b02ae37bce3e88937537a25429130d2e5c4d52c619f99f24737704fac980a8c44ca636a91494769095276edee5a13c53d5fbe09bfe319db10b163f3ca5b2c5a0189c7ec809f2ae140cd66591d2b2ecc65d160463291cef5d62c7e1acc27bb3e9f56b63e4e7e3a4a2140fee57cab5030e1aa5569bb5fdb158e07173de604d6fb9f162fc8cbeeeeba5f04bcc49a903635dcfd5211ffb34f230bbd58ffb021432ab0c1f257d4a4e75908b0d54068f47d6146d3e48d3bc033327955fc773ddff1e15cbd7aa35535e1b3859c9068c8d482fb110a4310d62b97619abebb4837f5108f9152c229258c1f11febcfbc6fb2ed930b60cc919afd91dd27baab8415a9dd0a521bc6206a088b2e70b3f4c32bb89a626a824e9b822b4d401fb0331a2ad0962f4763b46df260b7703a9b6df752d4809c2493671ef32abaf52764d92da3b3d5f785d963f4cc9d64d87fc96ec253a5ff9d98b940ffb899b89b9efa09cb239a571aa32eb7387ea3adf7472c051c3b8c0691419c66e7def86135bde1031691f8aa126d1d608d9e126e1f94411179ba1db21999a84242e4160b3866290630e317d839c9eb04a6121381f53ac80faf2ffae508b757488d758b1879c7eda1870d48d3c450715a036cdeca33266b88b88987076924815d44ec7060963d2c7e744f20bea11fd633c5e5d8f810a794db541fd228400805b836091924c889d48a710833a6bbaa0bb9a1601f6f8bd8ef17366625f4a7d7acbab65f8db1bda003586b77083543c0873bdf1b1d4ce40b4aa477f80d6996a916bb9858521378f7206abe0d70d1702bdf242e4f458aa377affcc08b6e3308ebefbd23d1f6e92049677aa61835664a2e6d1ee952940ecd52051e05ffdd8729b0ae55dde9940610eb401ccf7133d7a729e2e9ec36c21b4e024f80d12f8aaa6cdff8b938cbccb83b92d703b7026092b56f1ca5d0747c2c241ce38c035e61fb8999fbf10ceb31ad368bca843e91196b977028a292022ad9f063795d19f93c7e4e503cfb1f5fb18e9a97bf91eddde6b654fb33aac0b6eedc72ff36d2ca60811d5498cf53cd3cd1dbee59079b86c4a1e6ad4959375f1f05f6392e33a83c6c28ce28e4444a1e464e62d6ad794a9fcc9d0370b4367ed96e4fff411a5d0ba94058a1cfd09c32d6a65a86a3fd4d44c5b97b4fe7b64959fd25ffe29e4b61756e725058ad94cdee089138f9a5f3ff027cb7e18435f6c1504589149d0afdc4dcfc53f62ccc3f902d1559919dee9ffd1ad54921c9124a966b456a4078ad501197d3eba8fccace94521;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hedb405355b95994d58cf5780f08b16881440bf9a3585f73f218e2b19822eb6db98bd6e4a50e00ddef3dcd3e49231bc9d7e2aa1efb6b529633e744d11b7a9912aed280af78b6329b37d9028ad444ce4d9a8117c478f45c5521c460739f1a27647940515187637cda1884b641a51f4a74326af527d423bb92edacd88a56b6a7a220a7667a6fe4ebfdd8d0bb4f864727f94e7e33b1802ab99358eeab9712375a31b43a6143a3ea76ab19f1406de2fa5c35b6d58c4f7601db61ef01355274d197de5d621bda90c17801ce17d47a037f7b55cb76698c407e710c576749760415a5cf0a67f6981aca60a0af56a0953dff3d86c32aa00c5f9036a9cc1e7060c3d79eb7a41c63c9c8f23dd0234ecfcf5953f0915a27e836c1f4e38bedc56eb58e3096e6d5d129a1fa0cf9b81100468e8233cd2d5a7af2b38c5f691a7f69cd541f6e600e8db62743e5ddf30ab0609d2a39ee767dcbec73dab51ed9178d2a2a5ef3a2b17f0f45f365b40531b2500c67000ca48d587b022d672c86f7c506ed87af29302bdb4a61dcadca82fa3803e57b01321384964e6f96ddefc71a9322311d6c17ad977772fbbb46e0bc1881ea3d2af5671255f9e898fcc48b676875a4f10e25fe2cf838423a8c69b05724655fd21bbc8542eace19e22d39d14b8fe2541624475e06f21d4334867c8325bcc6b2080d59c60ad1fc660f992896cd29a6f515b7b9a3af46f218e13dd66d0cf07a184d2c9bb88e144c98ae24cd8ffebcc97f1b447d168c08401e643da2655c9db1883c4a34008fb2f43db3736cde4007f93b52ad280f6c120b6e3ebfcf7ff7f6ae5f00e1f6a4a9621a0ae0504b87494e48a0d5728c9a8e06a8eb75b60b83c42d80e115c3ceebce8b7820df3d9fe756a04c3e4223e17e5d0d363be78a19b0720cfc407fd26ec1f061de7c858a8213b34c07f17e468a0901c5e543cadf9e3ed333bb294e3b6b0facd151cf626eb2e2d9d4295eb478ff7d7f3e30d31a14daac202f803fcb291dd13ba980b281aeb45af428e6c5c3974af0deedb9acf5532e443f986d829f93134be9b9843b5ab5cca5d1262d6622dddc71dd850e5a9f645adf70be2b67b650c72cf943608e90fed35a2341c16ebd3b0bec9f35091349d04ed2f43b910fca5775c5b3c407dfa72cf3d0bf16c16ae78c370358958c427d1282ffa75cd887de5272094cdb317d6b608cf34361377c307d9241044945f91c118d900d6db22781c423f3ad5bd00c144ad0440f94f167acd34af89e6e7aaf47b5827627772af165b6b67879c866005b525b5de36e3905ab160bbd84ef9ab926ad9acff71fa894a722c247552aa35bce43f7c44c42af3f79f405b8f82ecc75b72b24a2e0a357d6487ae5f401f3bcf6bfc0ab474acc72add7f60dad4d915b33c731f75afae98a7cdec5c82da0ca3bb409a3a5448804f86dd322aedba6517151addebc0d04a8e5e05c2ae74abc50b87e6db6d23b1312d43d3d2b31490ebca0091906a51f83a3499af3931a4e823d2653bb970173485d1c3872f5b134d18bd62530d90f1731d4a50023c9975b3983d64e22cc96106d28fa2741c340b8b4a9b141aa4ce28b9edcdbb4f1c8c5a30f36c2f9101649ce1b9a5adf45f3fb86a0ea3aef6aa7e96b2dc0455a104daa996f09e49b7688cd866b8153a6cfb43c696ecca717d4444f0fe84706309cf4e0cc2d338e4930f9b6d7ebe4f4662ce075c5d0530779fd58349defb0364c0114308a752b6a5c76087784b0f0b1e07011d17a09d13cab5495bda3d7b8692c6e2df851d0ad7760c163d4734f4840d5d26c35d215fa98978346293c23d031d442c1f8d9240f290ae43e4bc5ca7554b413e51350c4ba1d12825d4ba99680f933c925bd1d30cf6973472371fbc11b44e7fa7520c01d7bffb5043bc6b4ac3004e0b90cc703a7f032928675ced33d2de5bcc01709da2922f3e820dbc0deb514d170181286b4dd287259a5a1b93e135b332e1643fa6abf2f47bbf0e9ae77ff46f786d75a771af581dcdf69b260d19e21fc6d5e52fdbe212eb19e5dcb46b8296f622b701b9e2ae4b8e4bd3ba44e77cecce0fecb9f40154abf3dec61eba68ded398df7af26bffaa126b44d6bea85d6f069d7535db8ac848c255ce3fd51c2cdf3ff3c9ada277e48e4b22eb523767f7112932d4028af0868712efcee0ad70e02bee4f35f516bc56eb54670e92900fce2bece4a86bcf565ee80debc73f00e9e8dc4b03fc627a96fc154e1f04eda4104137465dc39aa43c37afdb6340ca7ce0ee334113ee76b38d7311800625b99317f4e74d4189ad491fbc8e2be1f312374d0a128e0070333012bef2bccf94b00138337658f3982078c8754f56e0f16d1c08b422a3b58a62fcbf4b0e80acd4d3ecdc624b0933b6fcea19c46ec136e771e7661a2a25257bbd9cd584dab93b8542476e45f1aceb6167b670166c1acc3cd81265d10c5b94c4a1b5a378fe1d522a02b9ce84331c8505bec87339fb3b7a2f0702a60e065a7cc7365aaf3b400008135b2e9a4bef573ea87234e91b5411f3bccedc2d3e7c303d08178411462d20f0b6781693885a0108d313e9187c4c9c320116814fd72d210b37840524b3dc38e2fcc2526ff106bf5ed60f123f65a2bc05c2833e8767724087f0a11a3961ce6b7aaec1b4cdf319ce78869bfe172bb1f96cc1ab014099198a599adabd836a36e8b2369092917131d0c63128ea2143ad4716ca543feada23ef4d28f7244446b7e862807ca643b332507f41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h86a6fa18773dc7be131ccc56b8b9632540ea35ab281a0f47568b3bec3569eb83097df771e91546c1627fe9470ad1eef2a098e8c706650dbb005221bd08c5158aab5a65ddbae91ab13acb50fbd6e6cb7afb800cdf87710783f4cc12e8096892f873920c5bed5d4ab49a602dd02e4f81d10a3778a6f8577fac423e72f866978edcd226a3dc3330aee446276c7e347d8bfe2458654062177d417b24d4c831168bb5ad8d34af14b81139fec5f9c96a0312fa5edf1de6cc0a3f678bbe11eedc27df56d16129c8e1ba7b1a0b1c53f8810fd8521d1aa2915dbe0dc5b445102f1c9606a90f520d5ff94b09d51652bdbe0f60035efaae5244472832b20975423ecf22158c9e51318c66692da4d745864aeeafe19d5134ed02bb214a58ac29b1029dc7dd4171023bef38ceca7b9c16a5f7fcfbceef80b7b425900a9694ec6fc69f4f7ade1e5dd59707758c67d79e25d9e8db9d6c2242911df793b03b15d8c844ce08339c180bb793bccf7674d05424f278da36d67b943a4ba000dcf4ae47517f49a4d7881f01c00c4a5936245cf2e55dd8793eeccba361bc2212bb667c137989a585fac17b2d34affc2124a6b172146dbda7b0dc8d40bea89b682e627cfe753b5e96d8dd1ac339bbaaf367c5f1610568add5f45455462dc44d5ac723a9e1bf895679073b818888600eb6e118de710c6b40f334232272661748d7ac6d50650d5a5b0dfa83f0bc0bcafebfc098f8e8b543e6255f42da222c6a3cd9071b2a80d153c08f94e2bb16867f02918f28e237dfb42dc62129ca46c5fb97a852e0f2d5e208ca32c05c22644935aa3292cffe92d871b8b0a5e7549e13207c5a4e404ec1681dae4099b3c7179b5812a26e10f4ac499c2536ef0b9d1a87bfd3d85485ad84f40ad806b2e3c6bf083b57d659298e1ee85c36c17d0ed738ee03cc8367e02a85a7e6eeb40f1ad8eb81ab14d07d97850b0e551c9593b0a796dc1589e85c6267c75d1092b93fc9e7c8f2f5f1f640c435322da492322944f1025d3fd4d3ba434d93b0f42097ded4d7e1847f68e124f819338561bc8203e1bb2654aa6a08d5eb5574c11e7e477aa60862d9671ad6877bed697c634196efae26a615613e5d533aea67a4ddeaf898129d1ed79f0a502ee53ae3c3f9ddb32d65f16d78c50535a9f2e17381caca56bd1fc48d154665860b775b7a263a60ebb7c400947a6b62012d2dc39442e14fccfd6c0bdee0087277378bc4c7983f1063e5bdbc94ea4881d9edf041abcb0001c9ab1b75fd8af4e9a4517a4d79b74ff6ef20d0c49742a2d46ab86cbbdbd8daaa4daa43acc5f943474efa1352fec2dc09ada66f276a8aae2519072572f59f32987e26b9426871b455029f5be9ed799730af1d0045ecf89a1ceb07ab088743208efe5b33c278f0fb93ac62d0c66310312e97515db0cedb706e991461bbd527806dd80dda41b17ef7675fdb1b6fe49ff82fa20203dd4a4bb4c4b3aea3477e972e27c05ccb2ebacc6a022ef67183d5da5961b5576f9ffdf78cb96bc12a5834575be901be90e4303444e088dacbb9b401992b31c16c14abdee4c97471de0695f9e80b05098e2ea0a9625ef35395f96ded14fc38d56cd2c9d51d40d2966395dfa6e2eb011372f00003bbce1b9153e79b615ccfb6710affa67a6d2819f05b477e8f96a4609d3d0fc0ec802c599355a832076b908d27abdf207df1b5a9026ac9b22cfd36f5b049efcd7a9b55706069ac86efa21e61b31410f1453b08e85ed8512d0e5cd68b63fc59b2ce723f9c5be28828fac9157b873f19911d683cb7d72e2318c048f78f9fd906c06cbf9130f3508d945d7624cb62209bae9632d6ba4805ac723b5a19a13d030aa792720aee4f625c2ec8b16a4ec9d671f2867ea1eacda0c9baf236a2090d6f807133377750650fa14045f617b9ad1aa0bbb1043e521cc21b503ae033e89febd2c2598aa73eb2b23d8291dd91807e00c49544e8604aa2bfd989cbff14317c5b22dea6f0d05c175fdc56f8d0403eed39ee7610d918a075b365b2f4547880c4d72574cb9937473ee23e1f74f0efc1fd94bd8967381cff5827468bc509bd4fdbaf8d6fed19c2ef3be791e416a86690b21419d3d6bc3b74983e2aa3ab7f9d90b02b82750f115cba14d355b340611bf8021c51e41e381b164c313d4b79ef6d4fe7731a9d37e93a0b211811fae1c2b0c86618e497a30ee8d9f37d71870079390fca5d6d2722ad39f08440e4fb66f862f610db12b2704685b06f9a83ff541d204e22a83303a01bb5da888b65f20fd4010c245644891d4e60fe071af9c371450b5b2f410e36f4e289e89b02c6f7507421d59cb656aee2ec53928007973bda8fecd7a60bfe41dd67d56f860c101d5c47f20af6fb0b645fdf49efa51de139be97ce137d6d6d3853e8f7b7acac1c0bbe2890b700a9976ca6750c0de52565053afbf96c0463f933ac9e9fa8dfb00521a096db3eb30672bc77f8977dede4d769f6f0c8e046ba976fed8730dae9d3524c2b140c8890b4578117fd6d679e8a066f145e3e3f672ed6f670d46fed97fb53289a40739a473d60aea134d22e71f72b2d6d7dec9c5d633b2be5b53e38784b694b3366f6a6f427ceddcb54ba6473b9e1913a1d1350ac4d54135229f1223682bcbf50a859213d4108238ce41e5c1e781fd77323e8bbb5c6dd658bdf74f03eb50efce6d5c9e68aeeeb1356e0bd399c8c8014a18b05c1d94a288f917345f77b54fa27903d6cea5979189a86443168cc4b0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h65bf6c9a68584e743d7c05d25941f553e6e0898daba8d0b3a5b34154337a5b43dda080916aaa800c52398af6a0badef50111be9ac3c46b176aa5ff55ad7c445065b212281a82ffdb82bfb324ae5d6efda6bd95c4c297faa8a0eaeda954fdd3b01aef4ce0e37294fa2278b545cc74f2e78da2cd14027ddaedd3ebc0f5cbd21e07dece0c3caf6d81220ae459aba705a202b6456418511579021a353844efce8fe1909aabbf57834a8fa6ba6bdaca7f61d8c51c1d8b90f8ad5419dc220adc0d8ac9c1f549dad2c2e1efcfa66d1e2227de903812137a46565c4b32a07821d4acc8c03d9b5849ff906fd2496e89b32052520b4bebe87c86984b6344e9da309883a37cc159c41255da5de00718697fa3adcd9a471c19fe78ba4c0eca267541e429d82e2d2a87454dcf38d684617ea458769b00df5b65519fcf05c311bad5100d0310d85b11e607197b561e55467d6ed029b8ea16e676f2836197e26c8b65aaf585e17a1d93271cb7f7f8eee90b125352322ebb7e5fb6855cd13efbd882290d239332b0156158f0edd8d5fc1320c054374de4011632d54682515b50953327f207c40f936987071f1f47b767b31f81fdf249187273030d186d84f1464c548525daa7c436c6bedc9cf438df2737f9438cdcf5823827e72e7f5b1930b3c6a440502a4ca48af37743121c84d47ddbe294af09a230ca02eea0fe44622539977cf06cf0d27eaf6cb3dd0bdbb42de7fce5ff0dd4276b9506ee9fae766523669a36c62cb6fabb10950ab9616578374579f3a10c5176f2db648c430e723accdd494c287d5eb1f1bcf39d8c421b721eac1f10891ca16850b2701609b65abb447626e1d8d4450be914ffa425b13c2cc7a75fef0efb2f82f7147e6739bba3ca7f84497c7731f6eb1da4d1c1605e12d0e8230b7ea571edf67a2123ad088270b9dd6e843f8bdc78e5a3fe95b04c82132a6f4d96604ac169d43c4f55b037f25a89857e6fd7a9cfd936f6e2331e78a7e11721439f84428fa4b1b7e54eea445393248cdd0a1a4a948a9174fd74103a2be5bb1d24923943be0d683372fa512a2151360136af78a30bd7087197b23dde794d0b4cf655eb19ccf94960b3d30442832cbcd616742015de4d13a22ceea826c5d24545ad2afaaa8b83db419af72fe98ed3407639984929c2d815b144f5ebfbda09594f9b7f453d989c22a2a871d224b47d71367d11f446fe2604ba065445afe3c477129b2dee67d0b8d2e5b5df247d6be0240045cfd005fb04e829ecc69d99c6198ab3b46b11e4dd9c91b20988a22503bfd2585d0b8ca8088ff16f5a1add75545a23d9a0fe7664c9db25ee254817bd8e0493211245cf7f56493386274ac1a23197b17ea3f938d8f147d0c94a66f11079e8e61fe91e7c1d2f3387e5fa84a9defb00b3890d0454ae2f934661809a5800bce3b81cbadb679d2e3f32ba8ba08ddba130e95a36a339cb102f8450ddeb07257525962c58d70c24211bf98fa16d2546360e8adc896546e3def3e5548f15b06f913692bf9c0925c9f34aff045b53d5ee8ea592813646cd49a0bba8c1c0bd6c8e2c656b8443ac5da41ab5eae9726406f86f0b1e732091c4f7f14c4b47a277df2eae9287c646ceaae93b63009f92fe517b47d8cc6ab184366b8549f527a67ef696ba9158c539b7f2f5d9415996cb34a33544a29e8cfa462d4d5ad0b042b3c176a4d42bd25f7cd6a18bca5bf17e45206bdcee9476a38c4f6ae2d8a88c60cc1ec769fcadf579b914ea2a38226d01cdd37cb9317e80e891bd8702353b1bdef28cdb2bc9312cc857e706e239bfc05129491ff08b35517157f738cb307a91d650031cd73beb421699b94ff4263bbe85a69d9974b2ae8c266ba81f67c073123397194c9f8bd1c856ff5bb5c74c8388fc62668f6b204eaf85fdf8055fb43f000cad68592519b4030f07924634a6792eec21c1699d190596e30e2aa797580a765cceb3cf7da31f150516ba3c7cc3cdb980c96c2e01fc2d58f3ed474d97ddd8760b6b47183a53e5583fe01264cbe05b8c20148ebdad045eb8617162edc690bcb45b715fc60ced14149de9311896bb729c2c15d5e1956fd200401dce819e4f8641fc4626ff79500f8d4b38d4ec302996741fbd84641459fac2c5ddf1b085298d7e9560f93be9eaa5877de302e2173d3bbf2716b7e3ed9ad4c8f51f2ea5f1232ec22255e92fd3735766b0f6f9b29efbf24e7de6e180d924b93ca1028c4da4559760edba553729108a0910006b1d728a9706f0b393c802c49eedfb0b0b1d2d68c54d9e3c1eff99f66a1176bf5359b3aa9d2aea5e633a44b15b016871315b6a7609e3d75bee7cbdcdf95b9c3f3209054b87c4453d765550f192980af8658db9d4091fa4c6c7d793667e06af121aea3f33bbd779b784bc2dabfd963e3c5578975e3aefea8927de4c5efd36b8b24b6df91239897bce86dcf859d36eb91cc5c7038ab76ecf6a1119864a852a90d9e2666cdd65c9fe23bd9e2cbebae2db0852bff1d63d2d7f0c9b556036f9d74da134b968c5d9beeeca8b308b3c80993b0b9320e7dd6e4950b11b81968ef148201b7b3f690328156405b9d7a4dd3f656194c2754b8fbb3ff07033511813db1288a8277e312016b80a8b95d655c5924049877310e6f8f5992e28aebd7a089ce2b7a247da3969347b415569b10c6b0296a80cb913baa712dd219d279acca2731e4df9f6d270db029c26445155218ea84664932a2095402790b45ef4079166b0c1753a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1e8f13a8f8ce90c0cac6d94164cc672216af3f021c30bb5595a0126540708bbea73596d718dd4a66869f57fe00d8549dfeebcebe3b1610627d1067617fa322b01ae0a9e2b2e99bc190bd999dcf214850a518bb9659a87acf114fbc5d06d25abd4b2e24cb1c4c887b39578b3a8d7ed7131b3fe481d816b34a962f41993226b5ec7edfe547964a5a43dc1a994909c0474fe60c0d3f23101a8499dfcbebcd833991102f0a98592593d7fe7f54d340eadfd8875d8732d1611d3af1a9f41d22dcc93722a34ae8c46a3a1b8497ceb278254932380c1a5c8b5cc23aabb8662f0077da36a93e2e720b758a9c9628abb7e0396e61fe02fbb33eb7c44f8dda694ad2c9d4403ac17ee47eaebb2ea2fbe122c6abf3e3f2d6bfc27cf87af44dec4fbe7f0817563b07d9d221a0b0514468f318e4996aa0597b3bd8dc4267e9d4185e7c54fb72f53faeda3b2272ef8094890202d971a71e5b047d52c51adcaf58b085e38e16722d1f290e4979bd62d5c81f52503b29fc128fc3a5ba36cb69f48ca5823fa789417b3add88458d3be33d55c3b633b1d99006aabce340d8d7b7cf30b1931584f8e41d265b3ddc2c9eba5cb5a3149fe053e2b1ac453002408a5bc74e0e4cff37d69e77dd67557c918e4bd22b65249b5854a2fc6afc5332d1665b5cb443c099807e9f591b82a4ae0699b162038368d0ae3622ddce5c1fab9d2ef5b601bf39d9b988932cd8005cea60c4e56517b1c40f5fba48acd36d4620387e148ba43e577a3bee59940b8b6004534712de15ee659030b7591f527a8f09c9bbe6f6d976e5d8122f4a5712573eabf02516e614d2adf0079ca91c3fa2529e1234fec0747fd28fd0858750ed5e637b87ecbc6993702b76c683ea26c28419aa799bee409bdcb4bf21ebc0f743ec21b469eb78d1e5bb084506481598237637ea52313adf6b091cb0eca02e61f324193cc9b4037d027a6f4423ad9f8ad210beaca71f97328cd93472fa140dc89a8b2da7b54b7ab37cc4c2bd524dcbde6aa1fc7a1666786e117d13ee2af6d13e1ba1116f5449097e7398df0d0cb0c174982d430d312d9b9230241608262e6cd3736c3801109665eebe12f934157c3080f3b9ca00c6a773e2953bec2eb287b1d340a1de6a51450a96b23ef0197ace1ffc5225104d4f16448b9f4756a65ed2ad50be716e72d4cb5b1b491448cc93cf907ebea5f1209d3ea7c9f7827763c0c670829800ab7c1e0ffb74137c85551ad96fe139f2b10ad518e72915cf164dd85a3573616fb02fad32a7b54cd5312917f07726acbb63598191482cd5be19bdf7e20307815e15ae2a45290b351461efc1f25e740ae25ed1930121f5bcd9aaa0b1049b5ca7707f5efdc623abb4462cab12a3679769fce0528fc852c09f6f1f39fb74e2d59e07e856ef3f3dbf1afd1d709c0067de8a73de7f1031bb346f874f4a7c66906a9e721273ba695e6828173c43d664821ecab3ec370bb33a061bf98915e93eef758fde58100e4feedbe7c95a94da301a2fb5fab0aa07e40182722fd904a50729596c4bb6335be52b4e840faaa6c965df07f177b5f9b3973ceadf0ea5a5399e486b378c4e3af50320ab49690a524ff20673cc5f798c85bdd1c047a7f0b6c0d0dfa6d9c7ff4f6cbd60f815e0653ee7ce3ed0c30eb4916d33af8a9c48d9a42e7786c174ff948816697ffe04a56f141572191f1f3f4850afda6890228fa4bc1cbfd380637761bd330593737cb060e4e94ddb336db80c31db8c2f56348ab9e0f6fc5bfd889417a3a009810af78298eabc55cae6793298d4e5b98275eec7bff656dd2de16a0dd818e2be0145898510627a54ac1fac0791afc26feb7295404c5649ea99d9d65329f5604acc305306f65e77a424ea590d7b5f866266f02b6b44e9f61ef336134d29de7b91b58915fb06b1c6b22d68326dcffad4210057fe7bdd9fc007b75064bf710039376bff0389418edc1bd940e16bf7d1cdc50a67747ca198c960fcbed9e74e132fd6977b7294c5cd95dd9ce2d163ce593ec9b2d6661fef7ea715a649689355acc1e2c7501528e0575b9860b47cf78cd24a592ffdaf8e948dbbb198007327b7d406f4a1b7f1f5c5ec52a507a012534f482b38abca751d33e432d9bc2c9cae35d5aa235959cb619680329d376b857f674514c10fdefc82ffc2f793e4e5d056cd44fb113c97fadde57da3a149d8c68ee12f320c52c9676d335efbd29e8eb070488bffac2b61596ebb0e7f94ed6a3a94adf4b7a8af7840076e9e2667d09e6ecc3d24bd666f1cd76dd7bda0f1c9070ab097dc7a17d5ea9b751c8a222b77e71ec51d48497014116528e9e5873823667b3c492b33de5caa38f7151f8b31847d6e897f56dabb299c504344ac2912273d38ea1915fa71ca46cf2b657c2e9610ee8bed85ff5df17e8cf649eea03e16784679ffde13230129ccf4c891c2a0c507fba3591a1241b144c0b4bdf67ed328060cba77dc085c560a6de0a542047649eafa09d0175bb28d5e065853c6b40c674b9710f588575824804dc02d1a67d9ce0cc6a5c9d5c68f4cfe5820f10de2c9ec80d30113a212c456019519b75b9976d71d4c5688089cabaa834fad47f43e71d3dc46ce702f085a8820768502016a35fb25e9e72e591add74218b623cba82ecd5f25ede93fac16fa537b18ce936da4d77beeb647437a70228a7a36b9adb1b3591ef4b407a5f38c6e5f7b32cca065efbc5afc7017384330d9b0246aac4f8381a8312ed8dc46565abc75bdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he39983f4a5b0fd7cbebee25a6b6d22a3548b490647c70eed6c30f19a5a80b0d0b089a029fb8879ad055e282729d831ad86a5b1a392dcc1c02af48b496c4f7252a6da1ccabe4cf8fde30b0947aca6cebf514f42cd462e1c6880b373cda2a78a24fe1ddb364a359493d0a4dce341aeb199bd1288d2a591d42937c3470eaef98659e9554da313b8bccc829da8f01ddce5f83e3eb1c9efa4d5f18bf8802ea0749f4593b2c7d156cb9ae92dcb01db1b7f468beecdbb4e036303db15b23b7ca37c0c6ca829214c42efaf6cb117bf65216005d7a1fa7ffd0874555271ac4bde894879ae0b0715d90c31377e132ad75e36fc4124f1e5a2ee9a7bc7b774efec3cbeda7c848960d2f492c76c9db113c9d85841760948fb0306aecbcd4b50109520e9caff3d2aa02484f2665154d1a71b06ecdfca6244be927d553d647743ba79560608f07551234bb104fcab384cbf624949a1b0a2f77378c68602b6723915d1fb8401e25c488970675bda5915a41ed841eec06b9a20fb8edf65db3a7e125f2547b11b27fb0ad74862d90f4d59eaa07bdb47d1f7f9a2ddb84893ffb9332106f42b027c12d2994f6c3aa6678edc153c864ee22f216fd52889c10d876123f923f19430c834f2f0863116425b346ddbfa3b090195b855b98a09c39cedf18ad464b2f5dd07f6f3e216917c6919647fad9af9a0d5c0673fb35b07709e03e2c7cae8cdcf8c0e35497bd0670419ba6f5454c1856c0db9d03263f04d93d394a52458bc32a7f73f4957252f4d1e46d077df8f4d91c475040497a1290b9ff66f5a7b957bb70d45b94368940825d9917381433b0e1e36135a831411a355a88829c58389b51763cf840415e19b9148bc7c418a52bb8b4765b310b484d122ca0433daa691fe18193874e46d0b28d21b88e62b82df3e0aa8aed98a3d0919bc8785cc2885e906ef20a04e6d925f7a83671449d89895c643e425bbba190b2009cfb5883d49ae0aa74024ef36539fd2415434bdf0fa30640ef776a03d6085952c850e9dc2074914fb56a327b374677e46a91113c97632ef58a483e6c138535905ec5db45f50a94542218286e449c957b1bd6163bfdfbd99bfefba1eda7f39205b423b0c439bb05d4b43091c4ce3a141625c0223c1da271f0886373a65f3386be82a1978db390f79a0fd88f7a9a8fc3bd8f19128660bb7711ccf940101abdb6fc2af0a1bb3169908b47e76d7b165c016df3a3b0566efe27ca3d8fda838685139cd82625378acf2bcde4dc3cad9158c8b0c120c26d8a57c43c5ca9c22c1a0d8ca40e5de26078040eace5bda7962b19a0122998985353c1a303292666d050fea662428b433b45703cfa6dc5c3c2177cce59a28dedae0c3d9ae2f9b97e63593257321327256970c2c2462dcdd5f158c6012e474efe2e474e0c17fbbefb2b63a5daffda9f336f11bad5d55696ce11bbc8bdf7c530c03d6478d2e210161e220341e6ee33189d13c0799a5a25f6f833dfb5633ece74f0abef901f00a8b3d6408a68c498ab09e3df7a921e5038267468b8c7aa77e9102b72c6c84d528875798d4a336c825536183b2757c0c67a096b5812daae6e25a2bac701e6ac327e072cd2d46e4826d7770385d8ba4b0ffd1f5efb4521f7fa25a395f96a9b3e038ba8ed5f1f1b40efb8caec385e7dff72683464f6680f799a138f87e7a40fdaf4b1f4ef1e4e76a1e3d574c80c4021326fbd3e2618187b6e4e80b871eb8b74d081b65cb9ba3e8f1b3a099e35969f5db15802d5c65503889703010bda8e18294bd9e816a99b1d9ef52fb42a2e698b8745440d22d6914408b9e7082687e1926cc053a03d44bec30625996c17b4841742bbadbe7d1b167aec4f596625b374dec885cdbddd897778d6bed521aabebc5a6ac2c3bf99462188c58a8d5384ef9adda4a4844562bc560a4fa408553bbefff2b3e6f770d6d61da48c044a075235f2dae655d36d532593311a041d2d03e5057f1af24b6ccec4b2e708f20427aeb565a95cc65034ececc2e70b92fe1d5bdeb825cc55429d16805a1cd0c32ae30077286532738f95ad42f1ac7c54d84230356eb1976c1a74941964b2b93e23f963115cea5cbe742f927fa7c892987ac020bb09e1deddd22fbe67ac9d344ae0735a61c4cafee3dca7be88f3a1292c27747268562a2a78c4b6a28ba5f795aecf3bb3c02b4f414e87ce417905c2e84c98cbb846b8623052d4b68d9e6bffe80678495f1be1ac128c0ac264a5b629f3b9d703449b43b1ccab2fc22a83e8a2e12fe80475e0824e8e25ef1175e76df37f40c811ba645397a2749526a5007abe4563f6d6227861311da062497922c9e7017b6acaac7ea096d749485211c89e2cf4719ec4f4abe0fdc43b1d915817bc08fad293b155acff2b56b96925cd22e47466d32f8e9d8b10fe80a12f271a96342db1dd86ad2f8943a0a0bd855a988755ddda8aacd6b7aec6cd879dff743d3af4ec35ec85ee38ba4ea4cd76022999d00743190be4cb4af75e662b3b30b866d3750c7d5a2e7c898935c9e594188d848bdc3eace14d40f452f149561535775dc68dfeefff8028fb16d3406a3b2e1ed30ef3f9233c70fc4ce513e8bac2f481b4c25a7dea808b8935edc9b2153b834f7e77f22c9cf8ebb3a5bbcfa188a04e83420d04093ef7f010211a50efcbf93d368d98f6cc94cdaf1116232fce195348b5616002451a2a197849a7a2939427e61d140fe66f209fd254590c8ce0ebe7bb6ee770da1a5993a0c85afb1df05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf7ac03f68b51d1c423608182d336d5b0d0d1dab6ae5ac6f56b7408fac455927a7b74650b0ce07aa084eefb91d6b76485b3b65c7cc52c6253c311f523317f1b9aec583569172bf2bef4ed62d8fd4a227ba11849c6d4fce06d75bea1275da57b020a6663fdda31e2e275a937a3d7b42579f90d69a31a3bc0e9c599cb72a72cc41633768f61464f8f6d8eb57c065393eee4689eeb057063cbdc035c281fb4f7d1964daf37d77de862d70816384108b4cae5f337aa1d884f9fff814de4159eb1ff0411e88bf4ca1a5dc949ec53516b0946e5e58466155f9323e99f1bf06486b69084062a2b92ffacf4b69df04fac2d62edf227c0aaa13f153724bd560c19f4fa1ca8b70990a21be84fbe55b47678a926e52ffd4ded243f14a510ea566c2dbb5cb517b5665463034ca2660c71c855ed0bd09e43f1e26a10fd08872c27e70be8c9f836ade9d0d304a1f6a9739adbc679aef44728b823e5d20dcc596e00f2514c2e73141db0ce729ce283472d7f5fae88577b5c3ebbbc0a868fbee320d35d2275119a1c3d0ee0df192890490334e1eca0d252ae2ea4a0a33eca2382a2cb8a6e41882b29c802bf5d997096a4426d58ed29493f870388f9d53497d728c3a86b0e96826f3126040bafe92afde317add7b37bc8e091abedb2bfe40265251fa05a9bedcfd5376aa098156a1ee60481459c236fb382600c3f767c7f7bb436831610e7162a88df408adfb7498208868fc6efdfdd1d0d5a565bd4c78445175cc5372f99e39b4f3e4ae8d02041d6daafd967b95e9b8e7eac47770724c25edb2b376c3c18de4006898d66cf09c488233dd7f8062aa65aac1ff99957f4d4ab6cbd67f20204d92f7655d8c051ee7794768442fd17e7e6f6e3e2de681b63f5c14adc5d5cb48127ae6688783111be50aa6315bd0fa7c457254689d5f302415190101c05c29a53084c80a5e1395df4ab6b674f46bc83eced070091250ca7c65dfd447263612e472c8040b7c85b47d9e9fed9af840fd3225373bccadaab0eb4387706b4415be2a2bc8d969ebe2f46d452a94d2944d146f72044ff109095723cd057f7f3c1b462cdabb31e8feced4b5f9b2d71af3dd0e0c1c1f931ce11e543c266b5759ee2ea7434d8a550c1c5bf73ede4278af70f81787c9fa62233b51d58b0ad485f7a2c838c19a85e9a7c1e1018d7c46942bbc5e7f6835d1f5e37897c0bf6d89969203461b3d89b61d096d2d220f50af1de490b43f7021886695a68848656d6a9b233ddab263da39e2e495435f74cd10fdc98780b925a86215db6ef71c3397bb36b7d15cb9d643460273024cd2fa0bf35c00372d017582814657ebfa4e13e44ccdea335ca6f3bef5046ec2e28eb16ad8235801b1fa2b10ee9459b512ad1349da53a77312de18e0a0d9f7c362f5d8caf82901b05a1043b81ee3d377ba4829a7ced5281910f719b921c690e083d685a362530247a2c449f23d0181d02bec55da17c94b79b24adfb4855877493600680cb836cc9d5020e5fdcee08d7fb3e3d819e55252618433bf54fcf7bd3d496d5509ba1f2e78632acf34a88ef1709f21263525eda72a1fd81b1c7fb7fdea0461542cbaf4d71b3ea12ee8c11b0e89943aa47d63495590e7e7600c800fb54e11aa7427efa0f11b45702d163b2018a2405f46c933c62736c34cd35555bed70a654417a5192fb8d9da03c222ca6dc2caf4f4d4feb9d0de77c6b6e53d164f4bc91fb4147a586817defabcecf7405fcf7f8efa164c4401f1aa53a8063ec2f8f26502f85842c817e49d8107b28cee4f476ff729f75750f45167351cb807eb457eb5d936529b59bfa499b642256c985aef8cb688f7e8369de74eb4c3e4add319f5e8c25b754bfd577feef9207936ad9f26adeb091ae920c1c0dc4e5c11047fa657e6a32c10dc912dd43c6562be0bf249a9652cf08952c22ef1c77c6d0f947f04c59b356639b4059fffa1b8e49e58373f17a6c61a9b1491abf910dc997d89bc809545a52dbcccaa1cd1114a0eaf91f794c3e84f101874259c4031555b43e87ba89a79c2af0d4bcabe8c3488d19952b27744f6eb0821f41eca26c74f481d99d313d85bd2834bcf987ee7a72950ab5c2cfa0522ffeec931317fdb9408e8559ed8a98520e863bb47eb7726be8fd03bc4261318dd87b79c9bfdae746543ae23a00b646530fc843fc32f5af1deb4d8af9dda2c335a45049c4524d3b2e1131d861ebdfbf6b83a007810b3877a9ff94d1558f0f48207edd97d3a16397c8692ba89d7cc5b7c78e19b0dae46439bbe5b2b92bed7d83ff7f20a36c35024b360448017b7fc7622476b46d4401028d97187f74afdefe9bdbd002005fb80e6888ad937874c659402da00f78ff1b5e89fa179c3dacbceaf931863cb33bb6231b11f18d204ef821c58357f7db60571fb8f9c5bcf904999f41ec107871d2b2844d5f36dc5d4e2b77720b8f33cb0c13c4cf4a024dc139198c9d4b635a858ba3a4cd1bed58ac2574c12cb074258234c1c0a172291bfb70c3b1adbd80550989bc2c7732138a35b8d1dc2a4f75b705e7c3a5d9b5608fb26b00142c930de03ceddb05329a1f8d9d3bc2649b8d3504a97fe8a5630395e7a63fd1ff46db1220e77fa6244f2c1b2c2ecb5600e5efa48d61c258884ce41dc4332fcebaddbdc29454d1f79bc92307a53ed91829620632a5c4f6acdbf7f75a02015d8afe9571c61caa86032d99be244c483a93ca2e05456ce33dc3d3e8fd9e2c6f01849fb834689cc8148ab6fb7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf0560fa65c537dfa05674bbd637868e714e6a19fe6642cf189db2dd390140cfe90e89530a2ff6be13593fe2d88ee289e2b56edbe55885bd2379a93b904a33d102d1263f0e4fd908803abdb6a7c37d8594a654c082595bd49010805400d66ffe5172cfee0c4fae5375873b97b95ed23c7822d7c91e951836388b799135b7cff16278171c5aaaad37b89986273777ca95d52e5733249ebadc274004e93ea89c42376a292528b8a595007ea6a218f7e05a028ea351075f783544841d86c88bad014ab1e9e2a90b07a34ddf269b8387484e1e3110274bcce71b0852153c9b5d6592f6f36cc212b835be043610287e3a6e433cfd7f98b96c111fc0f51ac2355e89fc25d6146a5690fb7588707b2c8e0a5eab3d5cc69983c97861bb5aaf24a285903e2adb2204c47ddd678c7221f46cae40482e568854e3c82675076fed289226b8fd166ca66fed54fbf92dd650b1cba42223973e8ca161f2267c16eb8ece8a3decdc6170435ac126c731183285efbdb7b17c60105f19ce6410259b084678703cf7310fc56d1715eed9a7a4a6423518a74565af33f8c2031680c6e83450c919e60468350d0d57a5f9672df29877d8f5a4a407c6bdbfa12bb2518fa4a5a384689a3be249fae5302dbb629ab3ddbfbb0788e23a150d69d6ba9d7eb3d410c602c00671801d1a6d248b04f3125a784d53867781b754cf51b4f433abb1b6f25e9733a66390411e0c7216b7f595659c292d8801e0655100707a969a0ed4d6843990d423f45a878874981d429dc99234de9c6b2922e6eec08e1c0d6e7c80dffab89964f0bd40c78bf8410f0398c5347d0a389d805188c2cd7d8acbfabf33d68f15f35ea6f5d5e670e9c5cad24b14211bdfef0457f39bc75b7aac5b20051ba56ca7edc933a50cb80a9c8860a9078fb94979dc54bdc7a5f69f5d98a314fc051295e97b384badfad59723684d5000728592e1f32ed124a6641e33d9446be02c27a727054b65438657a46aa0da05c29ff400a56023d4dd1760ba6d95b0fd8943d494f9cc1cd7b10c208b44eb83895d1b01ae5aa97d4a404f84884b1f3d7fb2736448c5909cdd68e04cfdd4cdec71eb7aa583142756ae0a2bce59554b22a9b1b763aa8515f592b5f943b140d503de39af21c075e194a4b99c47cd7e8b06acf10f4426a639805e3ee7bc8b1bb0fedb62b7ba48dd10bf058b4d25af53b91b47145fa3676e348b4f9bf8f646614f9ee1fe75be6c629fd50e54b69fae3b1fb58c8084c1dc8c6f17c281a61a46b20df7161c7d1a9573d7801585f9797117d604fc0d2aba4ddd68d0f4f514180a6338315806f1e63a7dabea0fe2daac159982b69cd54dbe63c5d573eec92eb92f76f06d411cea7c2a23635a940d65aafa749a5aec65a80412b3a98272036c5a0e1edeecae5f6fca03d15fbe9317f4564f38dd288ed415af67a8e8ba54700482e915055a679815e673e840c7d9ee706a37365b14b692098ee61e432aaff2c9a3c4279e36be244a02a2452588b5a8ba901fb35ded5ec4a1b2b8435cf6f3f9c906cb0b472747e09abce78a7c712cbab998cf9dc73ed4ce103f6a6664109ddfc9f352ea875dc8999bbcbfd30076fc03d7ad4a0a1ab3bf854549b95185e123d4db8e6fb4442235935f85d3447f2494a41974c14d81e765b7d878ddd0f4bdcf7d5693e1b052a8b26acc529ca08ce3c488523b96f917e2130948976dc8e511a943fcbc9cabd79495096760362e8cc85bf613b6e3f4a8ca83a2dc02c4f6e579f24faafe4a36f5a0a01eeccec84be16c412b7e34fa49e04bafab557da98c5f6d93c5f0290823981836c7a38c3484398196a696d639342e50879642f5b4eb4f5db2cfe7670f389d4995d8ca810734f405cd7890c0d2f98f1fcc762cb742dd80e94ee381d7b04a1d84a1f3839ab73ad6ce65bbbc20f4889ab84b12494fcec3a728d534d87228a7302b9c99db5397efda846712f1653347ca31a0b23729acb567000edd8c9e193a15d0d7ad73ebbddbf85198cc7e706e7caf6857126d572af9ac059d633475e36899b93ddc6a26db85df0fb2065b08e828751d0a17acc93587da2977a86dd0f4004ea49a950afeaa9402bf94c8b6cc7364ff0d500f0a00af1ccd7c6140afecb0e0d8dd806edf5d0fa3ea2da4b690a5c60a9244812f0a5d15669e4a06d282155a92c630c5bc8f7afd64c368e9da0a22e4af37165b2264183554ae10cd306d0d668133d9ef641d5aafbb65a2079b432acb921e9ba36325b460065b7cb1856c5d2e2bac4441e81d7c3f40a8c2ab926b0c9d9c92c5ba7be3c06989e5e1a8372bfd3bc0bc17a605ccdc73b0b90c8267f82128e6623d119cf5481c5ff2ab87e68498613e194bdf31888a9dad9323a62792ce11444151c551ab931801d17bc2f7caf6922079d8000c660520644c581a32e54fe576af0bf96a2d92e283c20a9555f3489a00678320995d2c1fdb4a19c1f10158eea07473987d202c12b905f6b25b85abceecdf6604f6a80a25823d7f513fae84f305e72867c5d5c82796653afdde8403264d19e526c1d999b2ed5accf8cada8e86370f77c4439fd1f8960ca9012d30386976e957cd19df9f0abbb7b699922a3c52b5542f8c400b574e86079fa9323991f06aabf8d1c8207659bed1f737c8115502b26da6a3c6ec6b74c6d9fba91a7f19bfaf47c9cee9ab6e43f731203bccc79623c2cf561b699f4f23dc8e82eef57d0f6619ad13ec3de485f4f8f1a8e59074e4aa0f32a5be9815;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5a1ffd00678ac4a54cd9052662c4527c954c0831615a541219c30bf5bdf42ea01144959b450c0dc6df2d1cbb7f6b9d822cdfd288654b28fdb6cf13b5f834e1bceb02563c55068f05ee663a322e1886510df2badcd9753474c1d6cab6bc878aa575db335c935549b9f4fc700d1526eef4561ebff790ea50e91f0541d88554fa7ae19a04780a12c4fa05b1b9ef5d8528ee7a22850dc3f2f41ecc92a88b771947095204d4ca90af3f671d63835bfb8896985ee9c2ed292285b0cc42d89d018909008f50845fef8d80c0aafe685d1229a84670e88f63900fbb7508920e91bfff26572de190b7d09d21cd6fd38fbab52cc67fe4cf8e22fa38c066bacc26ac90d3b4424519887e2a217fc467f678411c59e330cb98e03935ac0721eb2152686577fe7a6e4a6402ab9c7f7668e638e91f5c2b6c9e8896316615adefbeea26f32ad65f1d04a3095980d035380709080ee657aaf509fd9d77251e967e4e19e42a20786086f103d0f0e27636e8de1fd6194eb1e0ce24e396419949004f146cc53d8c9d7276a5d06d04759a41ca757f706126e3b40e76f9663df2d783252c0e69fc4af2d9ce60f28fd086a809da2487b0c6a88b3a289bb9cc95f386abb4ddbeb55bce594c8d6d3b447072c5cb4dde03c94f2d736e93eff6f773302d028d8fcb1c2c14997dd5e16dcd718a9e55a2b9a140c36e77bd1e7e453a2ff7a8fa513547ef48523907514d6c59cc34104a878893c74ae33c1c03713fa5b6cd2c44147a400d03e275ab2d6c030e92c1d6ee7275a84302101fc459f0351042e60d6fa2791557a341bf996967d2e198f0cb38b97d54be72094340c83d13f66398bf7f10e6d9352d631cd367f05642d3056f2b7d50521d155f80b12857e4975cbd69183cb7293585bba06325ddf151102e7bf6c2859d064046d27e69983ac8bbfea28d9893b5b3e883d0dba511a7f72e8c565aa93585cdf98e584d551895ff1cf1cd5771ffe3af4d232dbd1a27ccb3c772c9b4938b782570f23ffd32359acd541222ecb8f72ca55bcc1fecce8324b3ba0e982cb01b51a3419843648806bf199e3445a15be6e824c9480ed7a455832e76504b2b5830efc90050ecb6735757a78b67d8ac11ac358673a3f4e4d0b6cde222e20cd27611683b624d65cfa8763a48758e14c941f89987a9ad8ffe38810915a14b1f63ce4cdae7873dc69effae3bdc2c7e97d95195865a1b9adcf1f22a7116b3b65e2a46ff355b9549b2fcff1fb86633f9977f746f4efa75c96031f4864043c80335683681c5cc9a2087959beda5af2299e56921e3c432634b3d0c7b1413226db55acbe9603e83a5edccd3e1e13e8808f042fd330e1c57e29428e3202e3d2d869c049d2f03dab379551625d5b3523709997b846132f259ac448151bd4c814c206fa85ebbb2be128b4e9191026ab5641a9d31a03981afd75a4d0bf1a474f7e6c7b108e93478e16ce3b35f6fc662644bbd05addc6375abf1ec19d2bd1e33ada85bc8fa07e73ee688190ed48c1a25d0edb794d6204f97229fc30348a398f9e6eb76d78d75135556eb6b6f38df2834e081ee26c356b334943e6ee8abb12d711b14a655638265c9e6c9fab0d32882944314009ac15d9d2ec98f46ec49ff64c55b76704d41dd39460a15b34d52db795c482af2ca2029bcba935cd1cf600abbc36cbe8aa296579dd77934c8946431098fec6de3cd8a08f32650032002b128d6ad4f37fe0f7f65e9ea140e3198f0e0ebf1bb94c4ba2c40c5eb6dc4015e95bbd7f10c7900b1d181d4cbe3d882b0b5bfd35bd6b115e4093ea5c039b9dbc2b69ed835b7dd734381a0b2c2c76934d6090fefa8557a2aec7488384c4a76c8ffb29cec2ed3f0d14d036090b20f0d12030ce2fb157cc2725c0888913bfb6314cd5fff3e35bcc773823ef2adefd429168da34d38970bd11c58df4cd7cd230be6f71a366f0e0abad6e9c4a8775d8d4498f7ebca8618a942203715fe80024ffd1a59a1903d5c5ad23f6b5d4ffaef0319e71d4ae6fb6573c624a873acf4cbb603e357dc3323b5d38d19447249f695a969a0e4c9b49a49009d6b9a62db12054a7bbc265a506a70e1b6c266d8dc46a2ba35dfd69f9222522d4f34f8e848ca6d3f4ee362a17462b8b2cb46ab7ddf71a2ccc4d3673b2c6eec23a8477f7bc49ade725f83c12fc3bf207e0d705115fbaba6cee42c9559a1ef4a1522e05c3c97b440e7fa3cd8a20aadc285be3e777c31c551fefc2c6a6242eeb8c104641e36dc152cdca6b6665a48271b29b8f6c5231a9e6731f1761bad14e5ce376487d5cdef7defc1aeb3b602fa5dca2a6be59752ccd77b510b57a3d6dbeb9eddd4bf346eb614854c3c72630c3d6b6d619baa4d4a6db01a927acf86c9df8b094d04c7e3c17ad124704f65c3e8aab9e0dc35b609bf1670930225cd04bc784fe50c322393e5a93c82f3c4565f96dec47e788afeea5c2b7bbcce7c5e444315ae3af47b2a9ef643539f4557ab1f417eb12638a59552e4a00cc59f1c6ca88c294ce4d6a3c70919261c89d771a33822728f5432cc21efb760b124755a11769e48063a1d6367f485faf717b3d74dc11555a0720eb765be13ba1d38b518c8eb353b5d972b412a23f1ae823bf5344f45608767a8a5f8a590b8c7b89d6f036af7620b2baa2424f133d56d6e0e55e4f0f8ceb99689e6c29a380cb73ecef5e6a860b068e4fd9f8fe98adfbcadc64e8a649796691574e87536c8c56491adbf936f163b728868b1baa02265dd25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb7f0750b22f2712686cc1d9f78182a210631b7e94f87cb18ec855822ae014c6746715f149de79303f1cd0cd262b20570478bf11b06cde6bf8d5c97e57320e7a07bb36597789b769409ac9b13f1890554beeef36a0060b1959ae18b661b02be2215f57c53cdf3258a04ce0544ecbb609bb5d60e1f348bc548e05c3dae1a17021ddd0d395d6c84afeffbad2df61b5927614c7011ffe6e7779ef569fb0f743cb79c8eb1ac69551b98ede49114f6fcd6e00436f405f48d514d481922648b440bb18cefedf35fa1dffb284f30480f26a100b36bdb9069d4c1f2de25b05e98366b0cfb67e2ffc8a24db244cde23e290cdc5bb6a330b23660506eb1968fcf9b2a8ef1538bf8023fc237251f24f6ed329ca2e1d6a7e07f534d0f74df19b7033b2f933bff1d5c7f5f0c7ee43a3a299fcbf15d97703bb862631531667f3974d18682fac100db6bcd13d145a3b4e2c1b8c7edbafc0093c572187c84e8c02c18c5b9be2606d43a54f08b46e0b2b595793029f261ae772770785cd56b4b2fef4984075a5e892fb9a7f5ba54ea3a5123ca841ad4ea5ebbb989344e83b2ef7b22959e34426db7f3360f35a48a2ba9c04bbc4e738f2ec7ad4c5030b339228742302f63610efa5c78ad37b95558f9ef4e67f03d28b4c74e79e9f9c1a39d2727ef027167d7bbfd8591a38cde65b5696b484afacdec61b521448ec7e96edcd7edf973f15f72d2b1bce0424a8bc7d3bbe351ad203fb15b794dfb4507d066c1632cc15e6bb56ba98711c56348f2c471edba6cf816d19a680ad3f3b99ec8628d713d9598e54b01ef5e4265d3a8755b5a14e195d9090f26b6e596296846edd9c45acf741dae4121caa29004ec2adb15b4bb7742f1a6106a0ea4a3132933d0b351f8f982764abfcb2c154f6486423737a4ddbda924e8a87f1b5940314587916e2e5e913333793bc0fd2de918b0d6f0554eeb10dd63599f95f966f61bba8d3c872ed2648fe019770d98eb3f331e4314bf1c076bed78eb909595131cd9c7965cace531e8437180361092ee37ace6f0409cc33370ca1c0df684851182c9e9ae9e0433dddbbe293a34e5638109cea90ca581739aa4252b09fdd83136b1619d0727a9899e3ef3af9d29723e6bb5ac6d9bbd0eca03e630674a14864203a4d1ce92deb8aa6c1eb1affbc37b40842a6ee360085a7e0812586b2d2a6717edf698565936a21ada2c8e4bb124f7f189142f95f57a75b9cca0494b63d8115c4acb36e59683d202a8bc282d75472c12a5fbfe310e23d8e98dffbfd2531957d26af6aaf9e093d699b9c901eb68bf27e9daed2118d57afae3f9c326dd826941f4fef798e370c3cf03a273630c36fcc0152be9753aa3d57568417a0560d70415573ff8dde113d59de73f7c71b6b47ecbed9d78af3bcae92a2c9cf2d45d7b11137b359b02c342af596452fc49da9a71935b3343f4961bc95a775f296a7dabfcb8c66f39076b9310df250458bb27e244ab2b9f73b6d9635b1a0a05edadca0237771c14829d3b832b8b991e6ea02d149584a83d16002ce93ff888ca6592459c478a6c01ef9e28ef3642e22b2004101b9c880950774a961fe5e2969b3e5be1d92713d088fd77cb0b877ea01be6c176b7f312a17a322932b9872f6b7e24db737df3cb92e1898f79fc25ce85d2b3c5c3e9cec1d45a9f7b4cdbcc48a6cd8f933fa53c10a49f0dc0165c434de2abf7f121a21c97aa19f81f82cab7d3c5e08821359758667998372bfdd1826c42ec4409525144f5b220dfe706aa187a80e5330a70059d430b855e5d3a3097d9c41023d50111f395a3edf8b05a120b884464239bc01543ef25bd56d7d99d5f001f221f0960854e2164a518215a08e8e976723ed73fc08ebf6f3c063e2d0a6857e5653ad89bd77347f0775cdf1ad35c6aa1e3183151c0bf7c5b2855ae01b2c2bf74b816b61dd3374de4b4e28947897da35b29581ef75de51b33e7278d9eb3cbe5f46969098b43864c7e4ca9dabe841fe88000128f35efbdb9f4f24b7ac0d2985ca21682d0d9aefd63fc2087c12e57ef8d4a92c9d4d13c395942de0cc526f75e39b69b831ec0bd7f65b46b6747579437400f306e24808ad835c83cf01bb65e368fdf54fd2ae25f43c66d40b0a8ce3132f0bd8884c6ca2381a76116676b80881d6d6735bc4c8b8c02b23fba16a2b9a01e7a49939486bc3e0701621e68570919dc1bef675e39629c358138c79b7a5aac089246ad018ec222bfb3355cb33352e859c890db88d83fc7009d2be0758168105f3189e322779a87c862d034b8ec9ffac3537b38d45ce61aaccecfbd99f968088520d21071dba6c34e2de10c011b3c70ee28806d35ca093a79b13dc0bd16532e585f24de29432d4747433e3746eec22e68a54117656a950d5744c1fd646c75e1aec6f581e36455410ed63f5b974b8c1f0d248a54ec40ba038a9a5162f6fb945afe3c66e028064a20fd0269d5ab3931afe28c0bcbd46ce87f84f1366cc7307e38b9a3a57b06e4f50e35358fc94a00031bf47d489f5230b0776aa7f9d6e7af6822804f9b4ed9da0fbf746edbd194eec3ed82222723f333752631dd3155685eb684f84bc2f8ba0db12634b4550815f6d8735740dabde6e0eed7624c5fab103697c3eb916729d27244a77039d3c943b823961f6aca2e3553750cad155686d54d7c819f90ddb4e79418224f45e664963d26886025cf83cad767514ee3d9ccb3e6112acdd58141e6053534abe84f778d970f721c2cccf8e45c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5e12ded49695cf1d0a10e2c7b1cec5fa7578ddbf16527a4a0bcdc44456d0417bb1001279c463428210544af34e04831bdfd91cefe8c2c91f72573190f41ee37943ecb003dcb4e1aca7fe30a4abcac57758e8691dad1fb89c96703bd6977465cc98028125a1068c51f9346710cbf15fbeac98e6f12b4dfde62a9a8a7e0c3c31023a794b4c9cd3f7311259975a63c5aee4862086ca7e020044a8e0e767f1638954361ca3e2117357f0ac51147ef6bfaaf76237c29fb4dc02487010e5753bbabcfe368cd2eacc68bde808d5c78e9dbf7b7f1faae6792b1dd33d6ce7cadcc87cbddd7607f61f1c8abaafc9ca51d2c8bf8bedba25e5ce9c9d6e2a87fcb0a1283917c35c8ea4f67cef3e8fc6ea40c439ab6ef619d362db3da26c0e1f93bf61dfbd3f7d46abf7b5e7cfe48f49e0500e62ecbe0b7c0216b9b1e325a6a67b6d16d4cd3593e5e780d8688285be15ff0e2d0c905e01322e1b1914ac3fec1febffea0d8c1db751136fafaeb4c32eb36eb22bce2219717301174a03f71012c14704185ec87e83fe755b3c4d2e0f93757216eedcde10fcc0110b73b0cff604a9e81909d314dcecdb674871fe2a8e976221fc9ca7925ff9e1b869005442126edbaf1871713deb744cd1c32eda0b5fe46054bc5645dd635ea548bba040078894898b2e3b388ea8036f5cac2fc5a6a8453328859f164cc208a147bf475769855fcbf676de1e6ee1030338ac2ae96c973cd20a8c3cb92989da589659a3095e8ee38874a3d86c7ea998d55d37332ef6f5f7d30c86ec1d3c8624b1382204ccff6b3b061a1c7ecbb8b6e6d64bea272062006149edb8c5df1e842e87173921805169fbeac50cfc829a18d301b648fa4b8e9f5945b15791b60cc8989c7739c6027fb6869bf5e588ebcddb84a1ecc385abdcfa603df41bfd5ba15033bb919c78f4345d8d84b1b32e9abe1c0744362c68fbe8393703f99949166e036f77ed4d531fae28f8b70d38e15f6e429d221c466fe663c0c4a919a6287fd91d867285fb16b86accf895bda8534ba85a52aa2137a79258ba3f20050c00a183516fccb76e8f452ff8c4a9951ea8adbdf92ae9f2c3009a8468dcbea1427ad50cb70142395affba5cd3a45275f4a9a993b2f7c2f4180f5c35acf9d69270a18db07ec96add6833a0943d96a3c1a0b84ea43c3568b10fb68d00416ff9bcdab95b75a4ee085bb0af719cb288957712d7d2500cb8e1b29f9c0c62e9c8ccb857b814658f45ea9d17cbde4473a0c837a25e281b17bace24ca765293de6f301f7c7436371ffe77071dba2ff50a6c491e1ff904f6a9187f3fc2d74e1292f4f053e8b7fb570025a2a5a0801c634e130a51e581411968dab8951b460bfd4c9a5b6c08747f59f398cd9e3b36e83842362092f8a0fb9c36ecf0ab4eb1c44325155b7b7972239bd4ca8fb8b9b54a801b6a36b93e7cde4940953b7d03f3d245460bf337b5d09227054a2a71838f99df64428ea124edf605e148da1ecfd1153681e1c4e498c4534643b00093cf4aac45c3221a3dfa0e9a60ddea96a78cb362c2b75515e65ab21c6da83f483650d6d75dd8c1f9338e38c73907ae143d30db9700702f456d5ba4171b8e83e225c4cfdcf12676df94d3420683b2109bccc25102688f006a3434535ee1dd48590926fe16255fd900add68c213a0a2de5dd38936ce70bc3375ce13f419ad2838a503b8090cafb5c18c2e4e8831dba7c7999c2c7d8247cdecb7378f28caf3139154437422120b574b70fd7e4b40a67de903351952799c5a66f341318c0547d5bbba07bbb7dab17e62b3eeeb84581958f754e9de5816980cde0234e0879c449317d782ce532b8ff712b460a5b4bc2355efa4916871b08700b949612660d81a8c28260f0e249c927ba9520927631cdf7ddb5b36d845051ce318d744d5346e5f84a5c2507d03dcdacd319826cdb525dba46d4c54a6807ce32f4d612a9b7ebbcd16e838648b4f1ff87b99c4d0053bc5f98e6e702949e8e7fe7386e8e08f28c9a2439e17bb16ff6337507c3a5c4b6cb0218edb09416883a4c6e5d8e6c4dda305bca2b812924150fa1d274389e3d4ae12b429db123e46c93f1ae833ce06c566e76ef251c8bc624c0fce8eae41ce92e515e344b35e1a1aa4d2e89f17e239043a132c60131dd101d8dc4a25c31dd6a272841c8a56935a36f1b59c36bc9e56c79f8d1eef8c227a1a2d5518d5ce237cd21beee3fb16938827c4cc3970481edbfc89063ca1f2c3eacc6a8ae9d8d2cba3e850f25603d5bd1f8002a9c25433c9940f61d39af98a20bfae6985d6143be5bb13d59653b8412de1984421f733fa197c1b67514df09c9eafe4dd4c817d4e9b71a53dd883e1adaf0cbe4af6c998f71b348c50306f374be6b538e2dd06bc9928f9c1ae3d74a437b55a12635c96efaf197f37ae6e8dec6b2137d371b45fec3f59699dbf3c6a37423d0b398084aa04cfdfd863cb57060514b60a0f27ef4387dcec246ffe94aad7ce72048dd53ca0ec231b9572ad0dbecc17b9b400f1296bf5da17dc5026710ae7f4b99743cf6c364d1085a75033dfb6d5bbdb0218b116960563f895ecb2a46e488fb399f5f0c471b12434286eba66e5166d175d5c9ae8a3bce034e9437312f75a3dd17f1f7cf49533d656386cadf1a2d9ce5a5f607f2a87c8dea27f71cb6fb21f74efd26684d431a1525ac3a80cad6dd06f054515c5d03e60eaa292c39bbe3eccd7b4a48510277b18f740f572bbcb6bda7bb65e81e439cc025;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he666f49248c202810386fe91aebd819fb184a272b946be464f48de2c5af25ce0a6ad30d7d1e52df8c929cff832aef0e1370ecf66a586e26667239023ce1eec0695853ebd88aac09cfe8aed0d3a1e9d4b0b48210695ec000b231407d9c0aa75a7afb679611092fc2a153529e6e115b6cc8545972c5276ea26db84b702080bb5787ce7a8572ec67afce062ec10743affa00452df4bd991c7305c1a0ecc91871fe3be8cd36defb285b144d945431cc28c9074407afa2f7cad75d57a95d6c15fb27db1b5ccc2970caa7b4fcfa9e55f1c80fd0e80b4354c8262e128999d528587faca83bf2aa0f5d9286c950815374c89a38369263298c85a24fd308355dad014255835309e8b859e99d2a4b6e040518e85e6f605f04599bbc9916d90e7b214cda4112b26c7dcf769dfa96926d54c39092d5ba4c2db26dcf91756f44fcdf89c533d38d100a8acf90b6049535ba58d9c3231c0aec8c7e4d606b6808acc3ac31dce926c940749b047433a3974379cfc21af0129b49b44623f4122eca86bfc57a6187e6039018898470f79783c676c3ce6d59919abf82725448bff07a585a755817270d88b4c639832ac9546c310ea50c548cc540b20020e7570c97660b2fd6c7dce857617e3b38b08710d10f377a089f66b4094e6284fe52d69d9ccb8654810c1b580bb887648bbb8c9a853d335aaa68ce29b118f9a2609db7d7737aeb40ad5b89eeee64424751d33bb88fb6ce1b17017f37b5af1c3369439f18b02b99f4ffb6a222599935431eead878352833a950baeab839e1443f6975e79dd1483620efa03f7a0b4e2f70c32609f2148c6f4187e3966ebb6bd1ca670be2bc323d74cab7bf0cf02544bde2109ba21a791013adbe429b37ef5487ea4a3fe335958caaceaa2da6a46fb924308ff6fa3b170037690a4debfd5c00f09fb2242e3d57300f8b55fa253675da319d24f00716f0312a4361993275eab2d5b3e146284b82b4144709d352aaa122c2650fae063d9f81e9977cf51226c8628b615322bb839c14aaafabe415d7b29d1fb16ddefd4e54bf227a7394d8ec8030fafeba1d395f58ce05b0553b7d8e712b0d656ecb20d10608f2bba3da59b70b6cc2bb62351319e24ed478da534ea41a4a5a1b4056779a8ce7cda198500719ac4869a509ba0143f5923adead4f788c341ffe21c5391e27e6b1dc49d2a7e41cbb737925e10892c0c2512ed72cb48b4f289233a6ad06174c82600819a83cf98de7c68d1dfa1c3f9f955ccb8c88df77d8f2146853f005a5179c728384f50b1d7719f48ba7059e0d879faeefa2736bbaf7d1ca0eccd6e674b2501cc595728f230ad4acb9f164d0be59e0d9b7ecc0d53940865df5e9b81d804dfc0ca16a7019d4c73e677c3191950efb96c065880fc283ed496b823c6e78799269eea4473a354d70b183dfd7b12f335698aa7b099e7c4216535ab9693d79760b5f6493dcfff2182de5b3c507dc17bdd5605fbec58f4e48a1a25272e43017536722ae9e7e9ac6a0849aeb8cca1afc4b4fa05d7319ad996f22d2e39755577820a3549546056eaf24d6cab3ca3c8208183604579ed1c4ba68fab9e8eb95dc56aedb3aeefa2868d45f9b352bf547965ffcbca1703413512fec21a4cddd86424f5d9c8a859e90f447710f5075abf096c5c3884c6415152c2af8312977420330c26cf2c4ec73a928c788560ef347ca7e2c2d8a13154e9450c1766e9849973e462bf8015f4dc88f2e9402b282ac6316c4535c68fdd1eb64dafc97fb4e3b9901dd7abdc36a12d8b33fca4ffe2bdaf43aba7fdef39ca540a520a337931f063a87153766973c062d73cb7f757b34f97c161bc96fcf0cadd575208749dfd926d89b1aab5f666b326ef9af0eed53b0290f08b90c85029a441a6ff9ad80dd76ae884af25c998f6ffe626d7a27285350528c032ef00eec987d5ea57004bac1ee0025fc43b75d01bcf5ff1a0a531b184902608922aae79aee55c1df906efdbe76c292a677d11997608e3b130d5259b980b8a403450624d87f5a48d7d888d1adfa311ddfe418e8f81e3e13798554cdf6f4e5e92788fdb64bb34c9efb979c37b5b7233cb57f4e16fe0d1048974444e2511a9e3e21cc387eca30e5408509637b25e10d52520dcd770f52051e5272ea5615080dac71065349ee4804a1fb5e5affc676ade920bb6ae17d5aee01f35557523f27573d6f3b9c091a97c26aac76aa4494755cbd448c308f37afbaf17c27d16ddceac4be9910c2d20d2fa92a6d15619b72081e8c0e3d4e9d2aa0c2e434f591d8496bce35aee5aa60cbe8975e7388ed71f71f66020d1b83f6d3d7c669b68ae08c96a4176ccd31ee5b8e2932895142cf056873740b579b4e8d11101a9a6e97b0a4df00f7919bb6956b9f4305ef363f9fc6dcf1d0681ca3abb73f6632bb663c7b954463bc029dd45eee953d21fd947c4f5416e8dd1c051d1505c4d7f7a2f019258f77731bd1135f7b804ac33dc077a83b44d3e19c4df81d9e6c4789a9eeeb2e0d2d5f8fc89b676456629e106e5f9a01d66c8b62fe12b595275cdaa43d49ddc29153b485e9d099a15ee44866dc0c554b5ada05cd3d2bfc602fe5327d6912371882fbfe9c9c773c85a09f7d2bd7a3793b3a44864747e750195c7571e3090e820b4083780df64aad38a1b2ef14565f8dfb4263ce0a508ffd215fd265256790dc18c0f1b2d95eb0c3889421563e9fcc9d20a3fe6d47f4827119f2660417c1134eef759cab0937b550315b377d142;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc2171e4c6dc11d3cd277ab90ba4869cdcd75cd5b960887f448150f0d6c2228801b93bca5a1cfa3752705fe9bde66837beb8611ad8b47111fb006d955d2ed51c02d3fbe8cce3e2c424f616e49b5676f4c96d65eca720de58665964dd592454c75fcbcd7607b86f0d5ace16d3e680f781fd068ecf00139cc156072d8287ebe2dfc0efe14c73d2f793d11edf4828fd68a4212bacec9d5f5de591c171701407fbd20aa47d9130430dac6845066ad82daca91c5befc7be20257e349b338f2ea07a3d16921d4a165cafb2ee37b9e474b388fdc1465b22897c66e5d9d2d15037c4bbc3c525ca478f12f5321e8d1c64e85a65e4811f7d9a3bc6e10566c2ee2553f1ff1fead19067d1d977ead1bb6014461f499804d675887501a3b2e6f8197960c9a53f8c174a34c7e556b0b5bdf4997b1797db9c7c027afabb4770e48a38ea631351eb3d7c080789f20b18e038e42c5f75cf4b43895f9525227fb858646f2d93cd01cf187ec87c81abdb1abf63aa90c73d5bcfe7d2a014445ad984ae1e1493f180fa46b2f61e5fce39e6983890b2841fb0b45d32d518a7eab474e227b55ab381d6df60a4ad5d09c2e7e7a3384adf2dd659e77d4232c8df3bacd9f5b197eb804b6130844ba55afae060653743d6cd9ffc6664941936a686a7ffdcc8102b5e61b0092139e4a8edc959d4ef495e3b72ad3993087b8881568baf3eda018fa2fce6f663fad25f78616d2c28b923df63544d74d184556a8271b8b4e6ef969252d4c1054159f6cdffa7ec2ebb94321e505bc372ff1c895e96507d11e0e67f1a336fbfa96baff92c620445e7d8faf5a6ac2129fdefcaf20a42772d39a26c03891749ee2485f39d983264d524c98616f41ce620011c025bb5e0f5679e9cc9f1bc50a3060bbc47c11c16cab5b27379d05201354f30f24a22afef4746ae66c1a037d7380dade016b52c502e590d6a3e9f930d6722980741b25f674a748eee306e1af06396f8d08b016aa4c8f02bf6e35bfce0c34cd65563a26f4fd08a7a61f618fc15c623d8a933863c8ae761a1f03f55a54803cd26715c14d15ac8a7953d3dadba544c80a69addc4a906682e5a0e4925fa39910a3e6d2040b409e6e846eeadd9aea7c7ac4d62912237c2235b50c64c565905406b9016467182f42933cbb4514118c5365144efad4429830a1a3e12bcb0736290e8d5740bb3020f456e389d68b39f31a408f5c905119e2318bddde349ee112292af5df35a28f74081f165da72ac8054cad85e9da4855fbea66c845662589b0568686fde977eeb7fcd36ae363ac779c256c05431a838a95e19782926626003969ddb6da9ec228b65b43e7e4158a7eca9b783a137f06c8e65f210422254fc0c6ce2772ac2dfab77510a245a93e528ba802d6197e7412bcb12e866dd5ea2d8eb9f846ea5dd1858516c91acaf7e60f83692665eb10e618a3270fa2f4d636d7499725e03e6df72448e9cf4b0339141ead6c08c24d8e40f69f82786e36e8942b477f4eb540a83d7dfd82897398e2832a24e8a0dde83032ab572218c2fb0bce8c2e69fe6b1077ab9fdb3bf07b36e8f63d7c6dda669dfedfb96abab328bda20c2060c03b1a1bdf81ae2304dc3da5e81c820f38c5a9f8ecc59972204b3f229d1038604b1a3a79d3faae332a903aaddda8ea13934589094d30d8056c1d6a819aa5a349c29bc2a02ffa14b309f5aa63b2dcdf734a3880ba8c3bb4e254fe9322be56c16a60f986db1b8887e5a5f6ebc6a81b78f8f8dee519c477b4a9838163f935df3e67473be6f40413ed6eee449ab5df7bd473ac438827b525eaf5cee0eb7fa8b9a064e82d6c585a32ff4253d5cf381ae5666c06d5968e6ef9f5089a3d644fdcbb1663229dd7b6319d8de59cf1a7792ca02655c09aacc669fad03b98dae1fc59a5654e5f0d8c461e08be472ec686f8a81094b983012b07cf95fc2343b1cdb8208a4318cb107369cf3c38a9790059586727892f648a2a42f8978df9eef2eaef4d90f147c43c20afebfb04284edbff5a45c401c80b0534476fc9ddf7e1992a49e182cff1e6054668a21a84af1754263ff759e5d9685ca82bc684afadf6d901df765396f2fddfdc5c933ed6ecce51e72e78a831f79bb6b32deca967a829c59a3bb6a47d77128340907d01dabb4131ed6ad97d853315859542352546db045f48d273cf991a4fd2a06f48e84a71a862a427656e448d7405320563c51b1819d6f9a729cde5272c82c1d572d9f1b07af30faeb1ca604b917c5e3e41c9a14af29169ab4e18f1e02b2a77c0c8e8c2b234cf0cfc82369e0c3f747ca67fa9d78925d31b2d9cc116de2d64c689addbc2926469482d06bc6f9565f7f77129cae30fb180f5b56d6a3defd8f60d06b4b86eb63d6b3412881ea3272a4a6fff9c62b224d76b476b14eebb10709066306b413befedb49b1d38a5735002159a16bf45be927222fadf9be5980d287eeb26c9967e9ce438109728eda6d0d38f637d81ea5b70e19e2f56073eaac6032459704d63fb5245a918b1e3efbed85cdee6ca3f1036b096ea8e28d17a3a1d965be5ce3f7ba7770189f5924a616c07609f07866277b95d21d2836d4e38dd83249393f769df448e8d8438744d7423827e84623e1e7e573352792e963a25d696599495c5f9e0e96110901e135b69ec707024d0101fc61e9a253599d328e57d11fdb51146e93e5fa95b03d9e15fa6781d9fe72fd60e993a78411f6fd8f1f114bebf1e60f748b2898085bc6e08ed206663;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h185a5a74c093498b46177b4013de6304967ea04ad4167900b3243dab90d0ffe605ddb0e89a171bdf6605d6c19a7a8eade8cf6a767c5be31cbf3ecdb25f210ef7bc31e8fdec5037a94c376bed599770e9934d726b5e0115a4186e0aebbda52825283a0a25d1fa8a70de7f52aad327fa4dd1ec1d8342fb24141dedf4ed32d1a72a3e5635fce8b5d9654bb409e226f19bbdbbb29a99f823d0ae754dd0a9b5fe8b9b74c388ef51095254285044c5c5e006d20f71f97d892d55daeb8f481117d744b2a81ebbab434142e2d4da1ef0d4198a1636d7fe372def5d95f5331e0394b829de2dc117dbf44492f269c007e361f2d81b41fc9ef2a95c206031efb69fae47c783f925cb32215cdadfe2492d6e8c263ec1460524b59f45b8f0588fd45c4dc58b14cf2676b5e32aafbeeac98ba983a1388ab4d4849ab0862a39b61a66fdf8065d17f8d3ece20d99dcc8f95c02c09c769178509d1cb075a49915b1ce9d7dca351e7cb45e5c68a1a9c6c9846af5bf526633212499d789549d3b6dd0d4d3593e60c784002689e55aef991b919fdbfacde8b943789fae7518f533b63e7dfa292e91f05b0b2f57991ff3ae72cf1021462789b78d8a39b9090053a8a5af0af2c4a00253ab48b4e128b15c3b80e02a73a4d95ad8c310a53ebddd303d9077ab364fe019403f7f8eefbe935eb76b382cb6160643f5c5dd355dbdbbfbb0ee57959851596617f9915404067f8c2cfdfc9c0da822c7d3795d19c7c806050a9e184618d8230c8e007b83503fcb1761ad47c3d46b86bdfeb36391d88ed0f9a9df9dc2a6c612b769decfb308925a52e25abb642f11e5316f8fab80c7e64f1c41ffc16a75772dfdbf3d3e03f10ddcc33ccc2cdec539f9d88f7f287c15cc9ed3a82df0d4363f90ad99943ccd3557749b8cb1a5770636f7786b26f71c00d7541665e3c40a5fcdad5fa9a144072d35c5ad23dcf17230db40dfbe4eb4977c1300274f51dbad22ce085f5ba3bfd35bfd639df2be01896e3b4b41c3ce4598246caa30eb8a0af3cdf5a76933d7d0f121bd44ec8f86848440548cdf72f4687d66052b046a2b56049215493a3c808be692dc2157f9340f209d55649559bd065fb49e4feeea6fdb253a8625a7abf0070a41270337c5d1b6731b2e10851cea6f90c289622da067af8874d7aaf0f496b9ca54217d68e320a461f376778359825133ad5020351d07c9ede3bcf3c9ff8e3a988406daf927c179e802386c18e8177e0d00a4be1278d1088eece27ccba944ae36eb2301159a1c61da5cf77dc67dee4d9087882139422b360e8a2c198e6bf2f4d50f4b65a9b54b1d2e3d83f8f9e5c3a35274cf56bf328a6dbd80f374eaa039744545c4f058192fab24d6aac449becea3b0d6597b4a4f254cb75760200c6eaac6a66117ffff0a2e3655733b2f240e8b12ee278fb78d982c84e0f9ee7d6167b765484d8a2030cec37d5f9031b7697d003fb0c28f9b50e01f193c1eee7f788e885517d4369866c2904f42c65a7437d5926568e8583b2848594f2e5de715fda3652d62b40f77f1bb133855282fdd9851ad4c62e7420446ba4fd6399cd8bd6fd318fe3dce057917bb79cfd7a7d5437ca729f96200c59a82bc50e8df033e51ec699f42bf9c1def72a7ebff8649fc70962b6a9668fc6abdd9e671eb85869235934a595abf79a87e04947b04a7d956c6512f948180cae134ba185957a4cf330c8741ac824b02a2f1ed4c6e31a12cb23e966ab465ae5b0bd0110035a5778d7d9ac27f20c77987b819d67d40fcfa015d6fa24eb9c5715c48ee24900925a22308982f5657cee474a756994b70d7040083dc81aec04f6c5e7c7e5e0b331cfdaf91a2b80fc7dc7fe2439873a17a5a59937023e52cf0033c043e5ab016d000689348df6304f9e1f6a4ea079459c91d4b361b4f953966f54034b9a51a44055c25d64fe5ea54f4e27d88b9fc1840e0365df9507808a0bb8557fbe6c2a63cd15b98af24d8d971a5311b63b249863e481cd23015706d346f1fdc98ff9e4edee8badcd1d9f972a59995e306aea3e4899b9fc8e9a905f8d8fff302929c7342c39d3e4ffb36dadf646d3edbf5d5be740c567b983a2c192abe120cc2e403e508050e21c63500e04e8291f3f1a64f36d09ec90ec53326536cf0fad916b104dcd70fae1075c746ef437f9b8bb8e953a09f1c845180e14c679d1f838fe713f811d9694828982bd19325412c743f404da023fa4ab913147209a1ed8730eaf07e99afc7b77f300e0c51a90486ad5d71eb6ae9de8de270c1d1181ad22e51690aa337910e8a0402cf6810a4d790baebdfb5bc6d6dc14d6d2b07d05846293dc33bc970d2eab626b73a9e1a93f7c5034f95c84ea4a12cd97efd26d5db0d5468163d587cd9ea74559a7fdf1bd4c26eda758ccdcdd44e453045ee3f750742ef7bc4b8d230651e941e6c268b9a4c62f747bf6c7b3c24714844b231d5265fab6b0e5e56e3fc58c665da49da1105a439b8e2ec44a418537fe82f6a5ac884bfcc19cdd5723a9ca49b59dda5b73c38a381b942d0b6ad08ab1aab879874dfea0ab76c6b83789a23f8cd632bd926e277061e855511a2d8537bf8484285e8213e81ae13aa639fd2126e28b4d99f5f80049a23ea03e9764ef5527856cb068e5e1831f48989754548892b6512c2f8bb91b2c237a4e6c081e34598181df6fdce07308630ee7d17be952cc2684a706c65a55656e51822ba5e2e72a170b9527b71668d2feb2c0a540e95b796a8f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb1af0535d09133dde0402278b71bf71d04e9df28d78af6b685a07d7c5ebdae08d21f8f316c9cc790cd75ac038345468fddd2bba7c13807a217b6ed6487667dda28b6a44ea42abc189ccd0765474cb2b6f6ddc2abfacaeaf67282c12238a688c3739424beb92fb40172c5b0b9ef130ce244ccc969b98dc3fcb23088401f544cef2075151c81318e383b547025257549c61f83223c3d74a5b2e81189ffbe01bbf5855ce17e4fd41593c131e6fe8cff5bff8e041075b1722e57ecd66a90153883d4d62a9af7524c82fa8f06ee28f06aeb215f0637ddbed0bea4c882816cbe4422ac426f30fca6761144b65c6798e382b5f2c179255580c40b802e1d674d6d3c339726c08c6d835d6602df364db1452cdfdc18a80ae2657933a5a7060e3e064d0b8bad4d7167a3bfec06ec8871d727f97d857076791f94de3f87b77139d70d4538ff1429c6d339de9d1d3030c0a4a637736f2ef9b4bfe48845d36ae056cf12779b4ad635469ae9ac165e67f0dafedd22859eeb40fcea00d9ba7fb5de4a1af764bc9cd87188a5e1b58f319bdbb944c5c13f9dda881a8a5a1b90c537bab714fd66447c9c81aee97e1db7c8dbdbaea42500129ae9dff0c73ebc21735dd9a3c82afaf67bc6e29019b2d78b1c6991cb46ddb6b25b289da64a831a3a753c12aebf0f0696a242e5c192f5acf13a53759cc6c044288b52d40d415f497fafdf7449d34e7f40817061f14a3f42d64ec9cf646cf11eeb946227939007e9af4f5e30cc200162d75f19237ca6932c549b5bbb51654ea18f6f2fae511d48126ec62767b1c43f0de4848e9bedc4f75cb3c45c9928f253dec97b72752964e92527847021d92d3f87a41af3d27243a860c3de5de96ca05adefa837d0b72f842af00263868c59db4e9c143468759f750616c5c2e672b35790b1d976a3f45c005c558c08299d715e99487f0702c3eec3bf915e594b3693b67d3a94bb3cdfc085faffd184ea7c478cb54828787c3f384377e8305caa245bb2822f96104a165eadce91cd3f7d29f795c4d296e7606b4602bba5e381af61afc55101691f015de9702b5046be77e884a6ff92fdf95b8624e007724f9382b96556b64ab918c64262adacab584b04df5c167ed155c0f65eab1eef0331e8e862679aac9737a5e451fa0d982503c980c7a59a49bed9a8ee3b434d4fb4cb6cebaa534753855bb31ccf21129cdf6cc601b08740e2da81a9c188cc16e86fe61c5863d295ee4604b68a91963ad2620012d9b817546918bb4ef9072073ee8f2f372ac307008c6bf4974f615f0b1db31da9bd033c13204a1e69d5f4d14eb036a007870c21775b73b90155e5989cc10cbc0ba98c2c166d8d140b6f1ae06f8e4216fd1555bce6d263b3d7de75cbe98c5d3de0af6a912de40d665695ec1af760f60f849be2840a1fd282a56e9b8b27473839ea43399f8dfc4ce6bcb86c079758e47dc52fea4d7c7b2db171e32dfa985d24699d4efa6c5230298a285fc20bb176eb31de603095acadb7d6ab094aa985a4c2a2730009491a4e865b822a21dddc2135888a5bf5b2bb4710936e3ccf7c001e23d5e2d99a573d1ef36dc9837acb0bfe031bb14dfb0259a71f1cd18292da455035c3ffdbc89e90905dc5ffd75e80c96885268d7b5e6eb1a185956ea8a995cddeabfa369afc8162627208f29addfe8986a629c3a3849dfa42785c71255ee6c72381a0f99ec6860a12f537b2634c738b216d1d40eeef73df2efafdd1de64aa47bdc45293a027d72fbd95a12f65f7f67f4b20808f5320edde16f5a1351bfbcf555eb6388800af192ba298b8edfd7bc4eb4747cba5da269a6d7ee44061cbe97607eced8f3d422a0cc84b93e7ff740eea43221f7f7a01ad17055753c3645da0ec8e77ebe61d2c29cc972ffd8baf37e5add6461cba2286699f2a4629f00ce62a4ef0535221528cd7d058e06442968d610991a12cdf1e84363003cfcd71a7e9c63c3920dc19fa6d97d9b35bda97870bfbbb560d392ecc967f1212f67757edbe8bc4deef9e40abc31e3d6cdec9a22075ea13cdc8ed7d5e338da116db0edfe77594822a97ca0ccc866fa0244fc73ecfd1314a85afd229168c451cf811bfeaa20f35106bfb89299f15db6f789f9bfac0ba6ba7b8d64ddb110765feb02e14a77672ca4297b877ec83c1165427169707d802a38513ce1516e35cfb4b1977b14dd031391329fe64b0adf86b97d9adbcc0cc1e366a8ec256cac41850e88915a74f1451feda942160a69629b97de691317af5d22d8ac34853444bbe8332724b8bc83d3b4e4e31999537209ac43864cf8b4f65fd9e2372b2d03ecdeffd072454e5c650fdbb92b78786325d2ca4da5bd127fecd202c84179c478b9a2b6ba68a2c99abffe6362268e72da6e82bd2ebd223ad66c8cce30c32e7e972d9d01b9887c3e370e3b284d73b590ee1958ceec0c2e99953467a2a95ddba681a7b22aacdb6758316476c461e435d7991432178135ce6d67c4d02128f98f804180159298e4c0d21a721fba977dec0d2983a60181d1910139c97a7e5ed2dbe7eb72fc096d6eb583ce765687c5261283496a28bc1697c4d65d2c6f70afa4eb6bc765c2861acc7788346be1b544a32bce098929ccaaf3b7ac076bda477d9cca98e98f4c4d67f1aad08867fa0e05ff64b817353522ae06f52f39ae41c826afb9a52c806bd8772dc7c9977236b1a4ddce2f3db29f5af05e4b9b780968596724ec329b651520d5e2ba56fd461ed54b4a3d01ed84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h96c920231b79b9f3d8061d8ebe6184af643da3d17103d3860e801dc6358090f2f17e57d3223bb023c8c50b6bed6fcc0bc57fac3a54317c07fce35b9813a04d8438a1e75da3d39742d6d8be604aaad3ec55e0a60be5b32244c23f9f03be492e99439733e80d7cc93634b3895939be8f97b40e2c7e93821cc02c0f26f27079d61269c4b56e05d6d3d8f5b78d29c78765aa38c2fe63566de98ba714b0cb3822905244239a4a854a55c7714fa56e3abc3cfa7e860db332e73237fc0a60f23169e40bf008d2e34873bef3a7b9d0c1705de4e9af235d30846d03c430a513cad5b4029d8e3736b1435795ea25a5bffcf04f1b3682aa2e24ca0846720804152ed137e0760b59d118d040bd15df23f3aeb79adf2d60c4ce720d8355885b8959ce2c7803d398a4f50aece62cbe42915e36239898ffbf10af5a8e1ca49dd86b8998900a1fa6274a5a81a7671d845a333f8107266b315184fc3aa93e9bd8b7caf32e356e1260fc5d2f596f3c0986d5720c0400f16ad307285efb1fb3b30d365bf2e233b4632220b7f19090cf6320122c51a62ebe8fadef170eb48b9472c07e307f50c0fc1983d1d203d18f67b631826134b1e0e67fd1795ad4756f8cd3f83c9c90b417498b075307189a208ea17ff25b307747f663fbe8c88faa70f76bad55a5e496b39c38081fcff84181871d1f48f2be5fc6b191064330e884b08a657e8ccf8b077f454cae9b8ff9536a5a72c4f6576a7f36823d3580ac2cde8cc7709e3b021355c852361f2518d7e3ab44f378ed38a47526ac9b6b6891862cd35e7d75f2d37f21f6ab1841939aff0bfbbd37fa3036edb5c3b350968522d48e99ec5f0734c9117d7669050fdd6e21727ccb225a5dc88c8ffff68992784a8b187662a0db0743d282b4bf2a92f24b927b348d1764b0c99b04dfee2e4fcfa53f647b0ee2db7a2ae8553adb92cd34c17829e494d25110ae584128893c0ee8bc74c63b44f1ac0e1797f2e26c9652c18bd8ab91240b78485dc51e74bea9fa2557b7613bc767453804fd4e5da75144d0373736adb16ae0454f31604e0c9e20bd04eaa5e51a04f284c09e7ed048fb5ee7b681e9feb2ddbabe1c34b9437be60293c654d409c7b274c7821615d33b60a25268e34eb9faa2f549be91a86354131d3e15e2bcbfd1b0aeae91bab03c366452df2764b1d18b2200241b48b836e6c79ab985e4129fc6749a76b27c56b6a2f6ba614ce433bbda1b2c0f9fe72324863a0889aa67494708c2353481085b85905bfea3f308e675674a5be8690336dabbb7c881f3b379162bcd00bce58ee4bb0584e452e8d59d3a1b3ce7586d0fea915e6523b77423f0d5b6e6dd4b943f3a60f696ade5175aa14c45292ac33225d410b7c7c3bc37409170dd8bc52d72b100458b784c104d963d6d5890d9d88c281d409c57c8a25f4fdcad39166d79964b37f8d2e12ea35ef06f011f9aaf8623254780b3878010e3ea912c293885813c74d207efd05c85fbe19e6ddb3dd072731b2633e8a6cba9b4f85c164d36ae219aee8e0229453038b9fd14f0fde680f4c7a257431627dde9dc5c3a8ec731b7a0f0846826fa7fc6a2d16cc15600c2a0f858bbb670fb6292c4d51f78334743abc942c89835c46da6af1f8665d0fb6e3122aa5302afd9548c9ad556289c4340d3e043c3762567a20bf2df4c713646ad59432f0211bc4456f480a63e230c87f73768a466436584fe4ec3ad446e24a22213d58d4a06249a8b1f8f3bc03acfe5d9991b302b4df057f0e3e8b80b5460f127292997091f9a709faaaef5e25947d5ff493734659e70f856295f7a91a0cda6abc7cccd738f164dac8611790e6416e9cb1b80c82a0e84c0dae72e9716e2b21f03a85240b19e6ffe81078f5aec1515bde24b93f86e2c80cfcf7aa920942d9224a70db6eb5b9c20b1c0c2ee4750b0d95f0e61ca15f5e9f9961d79f38371f8efb6fa21dba7ef02cc1744b20428c9a28dba1a701f211b969d829a7abb4dd870ce652fd2262c0a453648a3c0243c0bbe2a3d24c1d5df0245cce371d3d741806c889ba2f2b3dbfb75e44b4504ac4192f6ae7e1c865943cb4cc18672796a6c042aad209a97212270797491db9e0580e2ddfb2a9432e6afc639714515c0cfaa93e9edd988b3dd0b10110af08b7dec78985a456322a6ddd4daf2404d7c2f9011c96bd1a6e60cb5f82a8943c51419ea5923126f4e2e441c26f95a5799f0571032fb14490d32182c4db3b95d5bdd1c4d31f2d04a18152f508867741df83a39c752438fcb6d369c0ba92751e1084df303fc7c5c8e60a9193806ceb9d05e7aee45deff3a201a22c8ea9aef099e12ada2fc6dcacde97514892fd136a0453d7805cb52e989aad77b503d0a3be648bc4bd8d1cd561a6171f710e00cf7e3af43ece318a5987340c28af0adedbc551e9816badc8e7e754bd2554f9256a51863d9c3b49f477d27693da8092b0aef005268befd212506d1b1ac855d102c5e33ae4713992efdef5ae2dfda1b5b96ef759f58b9b2ffb22e13790f92726bc69f4ba319257e7be49a9de0dfefa16ccf940c1e0bba64a672e62cd8a86ba9deb03c4a067a456106db88b5a1af1c32729846631ada2b6737bb79512fff9f385f5080d605d3ef446b1dea0c8db736ab75c3fcc0bc123429616ab05c4b7982f409b47524f9fb7793ad01f1af5cb6dc9bcaeb110ede869d627a7f2fbbd82e511d33f9b350e79c3e9e76340a1741ca276e11eed7f5df03701016347df7815c66e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hebd1eed24705f19aa5a8a78192010439421dd3428864466bfb481f02c316de7c723c7bf35695a74a3fec716d9ba6679806e2b7baf3521287e1cf71686277f30d55bab807c29200caa3a518f65ae86dbd87370fe1a56ec3e2c5dd3168a4df084381d29327798f66f1ffb584f8e301f8018cee2ba33765646212f8d398fcd0e83e1f7f45b8c88569bad7d40993856d440b14a15f73ec086143841162dd5ecf807558f36d126394586aeb8ea2785f91f8a40ef0239e4891258be349b5b0190069a589bcfe087f5be98f4753dbd2f5e9632129d038e1d49bfe82baa9a4db981ad7df94616cd8420d27e32054ba9319d6291aaba77b7bc7d2cbf1cd3eb680680e0a579c9edd6274183f05d3c39e315e0a66b5c5f831899b4504f59204b4de604b4d42c05a28a26fd0ff4dc5ac7a10081c2ba3a00c2105694006cc5c2bde69abcf59da77b2a22853caf5cf36b6b1627cb0d7bd256805bb236d663db6913582c5d10bfe10170012a7e3bc1baf010f5f291aeeda4ab2a693bee7feac8b2fe0576ab3c2d09b87aaf4db2f85bdd2f7e5694334c05de28f920360b0576d70698f32a32e04ff8fc8ca36e73e9da69cf658db76929f258547c694367235cbfec66ca5f84b0cb8b526f90346f867b07f5b061548d10292657ba37d726d44000af233b01a252f2c5d90dd374bc312658ba722c2e9fcb7454d426106c86d17c01433209af251e37a6f4cc67390c5ef8917005fe66f128696f33b911b5d76871194e5e284eb54d1a6ab82ef42215aa70cee9978906e4b3a615209e3bf30343574f0447214be25fc19d52e2417a21dcde1b3a27de3598ccd5a13e42d671b8b2a50cd8be49475d93faa950966a65f79364c97c64b101cde9b0ea138154afbe82204bef68c9037c3b5fb702b759984ea919df419bc1ff6fb8ea7a00091c0a4712ab4ee5b56c8e27776e1cd0acdd8befb981d26c60019ecaa3e259e4825a9911d3a5dc89e09a9fa39a5336bbaf14ef156e0913ab3a04e4daab1de639347e733e97dd36e88df12057c255487f18a7633235f405f650e9f0123479947e929b6b9e062e9c44b1f655a5e944592b701668323822fcb7eee992fd95c9f2d28a469649244c75c03ed92cd6447883723eb1546052fd6bfcb366b2a4c042e22710b9b37acf7a365866f22145cfc9b52a282d01e81e75b057519114f27c657352bc48447fcc3610fc5287cdac40d19bef7e6a7b9da10caab64fa84ca6ce4859326c90ea8a74d942c3126d8f90e1284c326c6d2b94bd1767e9886d6a91e19652d438f40dbfe999693e7b05fc01edb3da739794c052d99b2dfaeeb917faf100ef23fa6b06c682763c35d51872b93d904027dbda8cdf37fb2046f97c50b3e626fb201b51a574d43ce2bf1875302f2db6b16adf37bf93ff67f970cbc9bd528dec43409f4e1589f6a5e24a7f91d1f41aa47e3496e2b25b917e976af32b93d07e6fb974f1016c43bede139261c0583f4cb20973d3ae1ee9e8d356e2935f1871201cfddb87dbf87f723e8756f5801ba4d82a8eff13d241c452ff7b1c1cd9396ce8cc72716266636da1d506ee86ee8ee13c792fa9985fefa389c6a346a0317151c521365de771fbfa359f512b3164d5de7d52520167cd5e00ad2a1631ccd5d449ab583b9e5b6fb06b8009ac7a84515541db43c4a247caaae557bc576832274446e64644cea7fc8c8e824fe7d125275edfbdf3075d81837d897d24b47e73d0db25a5602b0359ca46899b18ac0efcd9695994994d4c6fe85163344503278f1d625c80542e9faa453a94d6d94db68de18ec7b8c6479076e9a0cad3defa8852a97147d80b192dafeca1142a10243fd071722ab5e8d0094db61c1e6249907d3560ae603dd9db48454a9bde97973d1b1667e0477ec5654ea5f168ceef49011f4a82e55f1d9943a33b334292f2f167fb394782791a7c27c68e2bb622a63e76a6b9493ec722f4609e17b7635f0a473260fd75c65ed596f6d481ddcea02008dfcec0d1b301ce6fee1a331cb88e7f1abdf674ac758522546bffadd6db3f60aa7cd90a721370d0a8deb0d9f2610c07c54adeccf537ba60a1216c3ddc3f6cace895d32e100efa675961908a80d9500c009494f679628f91f95a287a3b471c8924f9502888c1d6e527a0ab64b7bdfad38d458097c3347d101477d702b9e044b90ba32a6cdde4ba3f9cb0dc3a54e83a58f630f3adb27f49fc42960885629ef2d2821df4f9ac7a1302deb68ecbfbd866a12e71634b23a730136946652fc5c4e291f3d5a99d9c328d71d1422b1f26bd9dbb5ae45482e2e33982a3a67da9f6d788886619dbde4042e43fe59ee663abbd824416d400ecd12ed518570164a067d4d3639ad4a56406e6dc11848a0de86313e85c71d74fd8dd2f449f961a20715c63f08b08fe77c321953362fe9cd773aeaa986c6547972c10e9a68ee5973a7520a3fc5f87b4dc83b98ced5392229ef63a8ca44901995ac4ff14a331056a5a244774df2a92d60c11c9c2d4f5606b21b9790f8b8b6f29ad2a30976b5a6688e5d19cb05a88e8c36250f2246aa6ea0f51527e434e7041d0ceb3d9b98c833e65e0b2bf97525f3361c348932f210869326ac1427d48c9fe081ecd43a3da61d0767c0460e34c3880e28d0ec619cd84cf202a22ce525247761aab5b9e5ade9d653c3fbd70b4407a3912d0ff5c5695a2692f1c842b4e0c1b190d5c04f5be4c7e89199fb557002facb6f9de673870bfb81094729975b8e2203c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he4e323d9fb5f9f92c86d7c696d6fc2a792e05e9d64790246d9e9fed66d37236e1acac6a00ee6c8685bb58e5e94fbf84fe58ca4fd2840bea8e8c8e45e88a3a29ee36cf0c94251348be8ce80222ddcd61471ed19ddd5e213c71e7d9ae0af2617a5bd6f164c47fbfa667cafef222784563ccac197fd5fa26bca95b8da1907596522b641a24e96487603f7ae745d89173e1438916e020924e8da88cfff5c367b8e2c3f7a661916e873ab68db498d4608312f484214a9b1f7660ad97d3c80d8e86e93829982bfe5c1efe4cf1b1e34bc073a2c55eb63a41cfb708225b97fe54788d63b311a7995c349fec316967c9acb16a6aa77daa697f2c3c45b9470e623344f1a734ec48438d0888b7c4bded553f3553c7a25251e90b44ae5861118fb4671582bdc5d1b17b26807c00abf1d1675d2ca15fba52a233299b82afe53e3dbd06c41da52d418570ec9f51ce629acf0bb7c1873831062448275f18babe46c714f72b9f0e5492fe329c85d4ca89258a369378c035f7f2cda0c2a4d20aaa29e1b836c2303820b143439c591ab3ce126f004ad5826edbc8f5d88f66c6ebfb451f7269f76e6dfc800200f77f1b28fe58df1e376bff16366fa4fd21996dc097ee9edfdd6326325b791a67d386aff72adfd609d602878bbe3c2638c731216b56779a54c1ee2616b4b8e914fa6c4b2f7f70b6ec52ead20a80210482be3b3a19e6c51bd0bc2da64a746c77fcef495c692658aaf241a4c9664a8c6a51e955507fcb872077e42a9496a82c21f17c4f360ac2b8109cb061e4a73ae6e2ef1fff5b519113a4d911ece53b08a079635150e899160b90c6bb302e0ab6c6e588e3ac786a71d3b9b62b25ef5ff407d56f50d51bc2a6a754f146f7e1d772695565028fe7d1f017e57459fe5ccb3a5fc1574e65b3f33e73d8fb3c7889d8e214a8dcbb9aacc37d3981f484c7c06ae16eebdb6f4cf992d379fcc34b9b26c938839dad016b62d33d2f7def47bcc3e559f13eac8da025b695745501cab45d939089d877301940c16b551814c84df2ab379bc56d2e3008db03117368acc660321eede71137a5057d1e7662b5ebb9ad3fb29524e9413b859ca2984c11e042a8ac6aca14a2d7fa3cd9743c2a0b724ebb454685b848e1688baca10c815e3a4710008fdad905fe21ded3ddfb05108987177bd16b6d7add2c3516fdf81b723b74e2e9b9e738cd3d2059ae4935dce03bd8719035b98c07250a3b6b9b45a60960496ef07cb37baacc97a35159b4bf9246860b6b1ce622a4d68eb9e62ef4692126066b5f25fdbea4f337a677fd326778a99a53f75649066c4dbe28594030aa688706eea480d1e5b752ee1f6c14e9b14af34f401dae51862d216f3bb0c4fee4b28b654c7e9fb164fea1005a0579239b4aae1e5c2aa651f30aad91c23b2f610650c642089fce912969402857be02062153a55f8859f24bee06321863902cdce201774f34a3f1913aba4e9db9de0bc030b68b73c96f2bccee6116543c69b6f1f61c2b592bbaf8fdc8398b83d66a8fd101e0554bb3dac636012c42cc22909f33dc734f2ae7af2a58e198f3d26741a903200910e340e67fd1bac526f735d800b6e8390e656d8bf9f8d0339bdc2f3e07be44c2bb7775961c235470fa7512ae6cc15c5e9429b7dddcd7725a72c3f67d81faffbd9e0145b6c3c860db7875bb87d3a6ab3053b6b04ff971298835805297f96e8a513435fd88e3bd8ce54a960e10fc15a7431704dd71953ea34930e8229f0714316edc9c2b5b30ae4251b9d1053e3f0b25bdf249a947e5bf28c048015ab35670c261b43c9a6b9e7ba0812a23b51cd1788bf3bccbe303f939a61d88051d43ee6746c307a1cee88091b86749475bf73292f074606c12f56ce050ccf844a282beb8aaca83f2530d501d510468f6e711b019fbb89dbaeb3980f4d35b763b2f3bbe9561a3de33d3d132cd2843ce5b9423f9efa2979e6b3d25a96f12f7b07ee40e2ba514d899dc2652dca6c60fb16af86853429423fa92299ae4aebdc5d4264e487ecb7806764f59cd9cff37214d5538a227ebbdf8c2099146234ad5962aeab43d2230fb449c61900b44383d323474085ed655b2bd6cc4657c5dfa2ddd746afed5b7b65536b9e4162ed8eb3825c94f73e24ebf06088fb3e5718e4b5d0bd8b3d4d402bf26635da30248edc390547d5754569aac015425293b83ef23b1ba94c0ec10dc1fce6f5f0574086ca1998fe17fbea32f08942288314d83eaea7feb93796d22c65b4bab17ce8463641d8c3faa44fdf7213fc1ec88fa13f790cd541f7c0198d390ae44c928d18ee9e1c331fcf87faafe458adb4adbbe36632d974f299d984bf26182587beeff02e1072d194440778eb49692d62dfc6b1b3851049798f098d0f469a3753fc391f042b59797e531ce31e995454e46ea688c649f11e4968d44bc71362b835bb7c299b896d952b8d1f33ebc132c91c3a1aa5d8f75e4cd922a9f7ac5b4bdd544387cadbbbd4ae9525c9f2adb7c6646341054dd47291cd21b85addd0d2a620e22fecd1680d644338d11f5ffbecde779c325f1ff5b3971322d62313a19c5633d89263457c006f7b6259cf625730a4b102251fd35895340b95573aee443036037aa0ebd1c378c15be5ebe2dc7213463556898d7d86ed2c8f849e93924d2101d6cdb77d7c8e653a5f1804f6e489d3be44d6f3e9bf0bd4964c66f3fc43f2f6cfe9514526ad2ec3b28d44166f301a6eed499dc71dcefee0bd95417e8df63037;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha913c04c608f0c77b4f83ba5c82e9a8ecfb573e509bcdb21ae4104adbd864b84524df73eb43c5a3531e34e40e2aa235cb9b117bf6e7c82d81620fc7b80a20153b0d52cc101570d253cdfb4989bed98a5dd4eaacdb83ae4de8cd080fdc391f6e0ef7e5d2ca81f18879880aee0b3abd42f56de930699bfcae22d0d5123efff580b7f448cf11a11b02bc78ace63a711aaae715361c197a166c4e3b8f0eb0e40077d44fb049330ece6352b99548742b0d37713125cf3027cee107fd53acc7f1bd5ab325131d9c573ac947317545713b9f2b1ee464c1f91b88c52c5ccba8d87a63e12bdd83d678f2c53898e8b3f974029c75498d1341d884ac6e64769c08b3d60736506fca1321961dd65a812293486daca40cb2da3c80f2945c54d78f1b0960465734422d45ce2410829d8ed8f5101a85966fa85f70fc7c588bd58fa564f79608a5a68385b74285d7a6a9296bbcaa7e9578a824a0c13229018f6eed80cac5b7ba25675246f004f19a279599089b1e21e39cbc46c6489dd9b0c94ec1e4db0bd700560bbd97cdf3db1b4701c60de6693945f382eefb64b814312eb55da3274930226f14911d35d7c34663f47eb43b327b69b4919527257ca11a59743004abe8c1f21b759c91bd2dd12ae0f4ba27a0db9281d7f6c51de4d4eccf29a2f7d6601be39e1e019f322d1832ff75c2d007c6808b3a045d5f55a90bc45c7c706d168b1dfb72ec81dbbf5ad41f1747ef7ba389e7cb9c9e8310d774e0cb4e7e89a67cdcdc2176bc48e787d1e4c341cd243cdb6d0af1cfe25970fd8e2f1b0007d03c7dc545e1c05f83ceab8b20d416ed6bb8fd440a0075bccb25ee8b24897ab5cb32a47a97c4789b18a200c376447eb5dae712e33d9cf38c1b880066609b401fe0f766fe3d05ef103a91fd75ef4de41ef6180c26be462cb365ecbac3a5e8e68e485548311a2c3f7e329b8157d05aa85661507367a40be00398de10680332233d40a841a64767709554249d6500b4791db004483077b851a097276e801bc085e3742dbadbb6114fc43e2fd6cddad53835ec999fb377f44b026059578241d17ff2e711888dfdb519fa8da71071677df55e509fb85cbae1b32fcd0deca04cef55cec87188241c44a7d9a02e9e91af5b6be183a9eb403625b2c28256cd9f342d1df9870e330b7a351053882bb09e197587f29228700fca53acdff92874f22b6a70e3d1deba0869ebd71138556cb0399a796aa14a22e1fd15f2b00fc0f5b8adfa5a27054a63e068c0cab5b24c619b7d6177604d1da61cac1918c7ff252e408f8ff14b8618ee81cdeddf8c3c6c2c1c530bc8774372963eef644fc2fa66d2c48f33110df25c94c7100a48839a5f071b02089e38eb63f38404c8b882335988229c542b53268e28f32daac8cc63942625954240c842d196867de45baee6104759a2f334532eedb590cdd60622c6e58663c38ba28199272d4b9131f3fe84204a4e8f59176ccf63d825ab30898b80705732275fec5577ad7238bc15e573501c851810295782ba31a6ae93a71c101cee0e7ceff53c8e1e558c2b0772fdcd196d7bec5c2e821c65591226ef71593503b0426568f0175f4a0c42c04b1d12c058b7ce046672e1d8138afed93c81f24a5d6e9d0f8b47195ae99fedd75ced0ad3cce903a6430cd86e22fed3187614bc682a4f43c261a1e3b52109b710d5cc9bb660242024f2b6563129a10fb65ffd887766cf44c03bfcc7aa1626b0f297966c420de8892d7458e1d8545cfc5dbe963eaa93dfd6c48602d6823a549c3ceffba140d985794cf0ef9984ab5e72200571ff2c9fd94790702daf229ea3a0c756cbb0ef71b7e683c9a05bc5aa84f1e27062949aa4e8a76ac2f901a6b83133d469cb2aeff424c4fb03ee265583dabf5f06687e9bcc57661e508359961ecb3d035a4723c438cb9eddfb2884803abbab9e84f4eb4e2f98c12aa4a8e396c605a5301c680e5e28cab41858af1d06f100a6d2aaaeeeba6247d57825b50f5e5e91613bea72ef7194d8ac8451cb69e1f39b8830d629a0a5c2e46978e7a60406577b8f26ea9c774ffc7c903712592db33f4502ad329ee03651fed7283947beeb56674759724ca32308bf22c1d84c8ebf4074b9f435373a35dbd6f092353b4626779511faa3acd2e047d3cf55332e51e294a44d65e90cfbb8861c36d0126c0425e6cc342995e361b1691b1dca11272c598d6dbbe8332b19847ab5442e4b5b71274745dc761a41c7ec544ea5014b96b06921beab3e9b18c21ef8d72c821728a8c79c0c9e2922843b78349b6b2f45ce1fb17fdf9f473ef8e6b4a22bb254a066bd77b15800a83de02d355c98c5608eacc6f87fc97d55a3b8d18bd2ed0d4034c8c316540a135da9c10d817a086b484baf74ece909f46e7ea00dfdd84d1f3f03b3df6edcc40705f5557582cafa9b1ff0d8a1db11ae7d9370b54850684efee7c285ffbe5946d2a50a47007d7d68aa6b56211067a77a47123d09ccb0795d4422d2fc678c39fd16526d1e73a563219345239b1ef810b88e88fc0a1aa128c751c427f806ca3d16707f37c9fd7550b51c36eba7793b02241fee08e93b41507a3561aaddb25cc119d1f0a8fd362a08429cd0f8934f52903cac626115b595a14e8eb51d6826fb3a2817f4e2caa2a5725f3de558cd006c12f7c24bc29c415f6d1389362eda1884631fcbf93acd93b124f146a1be190ed7569da65c48a57605459c530081e652ee6fdb5d09033ed6d24ff5b4a4e88f3b8d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4839e17405242e13e8eac84a96b6c6ee6bd9a9c82682abea0291027c2d0797e44875ed683e0572c0ea4cbeb42443edaa6beb0ff60d76a48643d6833fff4b5482cae94f0319c887746d0edff55416f3e5eeda3afc428a3d31f8062386052451129e084ff5aa668d32e738811bce9b34d11722142de9b4ca59c082025ccdad8240abdf46cad55c20075adf53da206b2d43441f30b8d8b524558ec36e382da65f60bb0d03ce65cef29e2368a43ccece4f39b26b483685c177c2ea0fef3230ee0c33298f2bca748716ec365122dfcc964a4e78a6f238e61042f4f6bdb9d0fbe42fbeb2b709a5ee106fa5a84fcfb968acc3b65107b8b3315c4425d901eb166874c31754ac30f3c25ea24e3e7903837b7d0d8f77d61cabe403a929c6d86164e147e8c77f94f9ca2407d5110547e8ce0d2025d4b57d2c155b0add932dbceb4edbbdd5287af0cfe4a77975585d345b684a1f3941bbaf7e647862d83ce327708af030c3c2881a39ce078f7e2fc87b671d8fb6f764a6dde576f9efbae1fc7b35c861ed87668b473b756eeb5d1818d284e0be157780ea213d988d6a9a2cc102bdc7f7254d586f172bafcb3ce89919657734c6619f0a439e318f39ee52bbe57acf49887826efed26381d497b8284c63d96ea0dc8743b6c86b65c21ca1170ceeb8203f1b0d6727bb6191f9d32605b42722545a72011e7826803db16903c000475deb5455165e981666acf0aa6ed3839757e4119c9d5a5a29543c81d2316d7fa9bc45367b1dbd1c109bbcec72110577d13c17aa693e772e3bb5b7b01c1434b5bdff6e05e0189852cea261bd1d7541990b3f40be7d93f1448eabd4834ea9e431ae8a20ba6779d3cd9f32c9cfe9edd425d91ff8d636c5a849d2196e7c2123680638c39509b70fb90bb80e01b2cd7c3d599f8075ef1105747e0a44a2ad0b5b44da93f1d27e8236143f3bd0eadeef683ef82abad8a70011a02ea1d35d30fd60f6d51ac00575778de9516b74566a53cf80de2d9ebb245ff44081289f4abf8b789ba25e1cfeb31b973b42f1d566f83bc43232fe3f2567cb0c2d6bb7fd11166efe27f6aef51a9e6bb7017667470227c8b3f3f49846a31ff545bfbd33e3cca0f66adad29655c8acad0f81334581a6ca7f45559061ebbd35a243fb506770efe370981a794ce5b441d37c21bfcd9fc5ee65865d85a1321a652422bc2a74e359d249c77c4aefe38213ff09d61b0d2511f13de2158686f7ff7f02302754342484387c681858181b31c13fc3acfb7a58b86dbc6809e7a57a0dea0b0015fa2c6808d907c2dbe50ef30409ef402539744bdd357e1f032f0cb41213b90ca55ff59409d07c6a50e16f909a2736d4285ce8334872b81d45bc4f8b93ea909982dd3cd889a23c0d218c498a9568d46f2f1313c64d5b2620a807621bf10f129cef17d3067c2c59ac4764bccb05aee4a42faf23082dbad968c72cbbdcde4585d11635020425e4017757c47f9392ca3dbe7b5533489726b3d9f2cdc2dd966c069cef6ec1a8ca76eb8660a53ab075d93dd1f159d57f1744946ad6f191d75cca9366c1cfecce0fb2bbbb54d5373678c4c6e33ea7d71a0d9593ddc3ca263b06130ffd172d529c1e2f4a08351adf0f795cb1118a68eb77d7ee0c4f564e26c329c164569d06ba76183fdad472447adb56433604dd263582669324acbc7e843d0399c12244c77d4f15a9f937f1515295dce6e5b3a940573eb8ec0dc7ee8aa599a467eacae583c6a9b3d7eb22bd222f80c5a8f10c14f67b45145a6af1dbf058f7bc8998814694d348d01113b169327002784b1e47cbfcf7b23c722ce92d3e4bc1c886e8b477c5bcb613d20cae1bdb17279062aec0ecbfba4355631a643af4fcef623595bee13337b4a5e3e93a5ee4196133733211bc7bb38fdf65c7c3e44a61d49004392d0bd6edd13a2122eaf77610a013d41ed0a627ebc9c52e26214fc0b8a4a0fc86fb6f5b12580cc87e24573457cdd2759c5820d4a7ae6ee33f38cb71db1356c4394fbc2f3e3b77d7fd9bcf5a6214427649ad33b130a889ac040177b8c964396969b0cd8962592cc426b1f9ee9f850a59676d7b0a72fea07da5f0d85451b88009198cd85044ac764d1cccb0ee325825327df16c0c9b5b3b112ace88f2b1fc8fe6e687612556fd22ef894ebc9fc89c7700753c49b9272f3b02175a9d04accc1de1da6a7dfede06d7b10ea2206ca539abd90ff97da7075785873bac87fa042da521d05865560db0b04e9eda50b398b8c55d9fbc399f1e20f1321c3de1843cafac8a30cb4538b32439ad2ede2b8b15fe1589a763b792c4bd936fc13d72220cfc5eece8755b8a79be3ec8b1adcd575411e06623ac8f14834e52d19da0f37ca2202687ae8040258227f12bbffb8eef0549d5b2ec591acf92a4807b976a1439fa9e54ac0472337b452104f8ee10820b1c87a2171aa3d786275aee861f26e088124dac7e9aa2a6fce63feb8f56e9f7b2b724f2face28fe14f2f55c8a4f6937eca22a5dbf5d3ea51d6520de31395fc7d69727fc8166c595b91ec515f3427a004c1d2eef04fe60b1078c19a616a81b32b992754b4b7ddc90320cf8830fe31949dbfcc4b120239ab79a90e629ccaab793c903fbdbf310a6c39647e3c4ad6daf2a20ac312277c27425bb2ac3c9c112d7134419deada8ef33a92bf8e584383741e43a4ef7b866359b6b461f6b75bf0fa7a32b74b08ad496452b8d68d34782981d55aae5a804bd10b47049ed37b6f39ec01cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc28b5abe8a52dc1ba66a8b3bc2380a3572377d3ae6fda98bd312bd28fe31adf9b509fb71f3af8a7c7c7a261add165e1093e43d5eec5e5c4aee8af43ec8d66d5957af762f9f20f864368e2f4edb240912709790c584553d46717b50e53b69df9a7fc017be9d8726f09dcec7b048de33738af39afe5a477bfac629d082df951a5d8b926aee7c50e28ca68639f1d9411fe79dbd645e8e51533429d56df7fcddab3f8ace6c73d5c1a2a264caedcadbf3071e954b0d80f8ffbc608ad1c0f86389054aac0b965e5bfd263181349f0a4a50b61b4ae8922e4568859597996de7e0b3208125b0a34a17a532bf899e5b67177fe03a85cd30cd875e311fc6a799d83673b58a1592e4b0ec1f3ca11b690b25ae23bd791c36b72b00f2903eded160bcb2199eafd6609e6e605b460656b5a4da32323f88735343d33d5f5d77fff507335e228700ba66cfd7e78cc4219116b7a125fc6fdef071f0374ee7dfdc51358e4b77ca940a745dc55257fb28ca0e094a7d5210de9757db64f16c5dd48bad471b48a79d3b94b784d956db56bfe1cc178a1575cc02c9709e9edf0b827453c316550d1d13ba6d6605baee873a316334174bcca7e842c15412bc20c7ffb73df5b951d4e8cf195cb6a97712ed870bc71e51504c5961e36611a45b7f83176b99b160601e76de247b3b33682f6d37d1bc963c24cd092a6ac0ca654df9537fd29ab7da2f75e077b742ee9f5209aa2b21864875a65cebf20a5d99e8579b8363171f837ce2e6c11d0b6bdd5a5116dd5c707b62f4d3e147a427a89d01578c3d8c45e68eb4c52925ca476dd702a3da0fe7121a1d22ab84303566f6c66d877b8038cd757f2b231e58816fba69ac9462ea28724136a3f93204fe9774b127f147210c14b1040fec682fa9f1f9d6d7b86be91a49daa81ae4bf891e867ee660ed3555194b047402ba180edd5a87f7cb64ed02b74c59c4720fdefb2aa3b300bb196c6b9b6cb833f37b19d3ae117fc8e4418d0a3e675412ecbf91e37c794b757f229518830565fd784b4234697e2e753492b701439cf605b73884cc69a4a0759c359f948d92eb73ddef74db952e9fb94139e9ec6445a1a4392f24d9f1f7ce61fe0a74f7f1330eef02400129e2d471846058e53dec6430e33dd1c433d2ce3e6bc1bc3086197f032597ef3e58e779d85a3ca98299103faa74f97b939b00718961d93acf8e318f87a38f3ebddbff5265b62b1c8e2ab6dd802c881a446f0d13c7196512a6f5de37c048130a234ca273f96b2aea500998ce2d0892fcca9d69cd9b830660948f1918994cd03e3c22671373008af08422574dc64d26e24cbaa2b936920115bd1a0c475e3137d92619010e83bc00ea254f27fe652e47ed519805592283845547cf57e6bd4a3b96b0ec0e135ccff6ca1a9beeb35fb28442e21fdf37ff8f34dbed9faa65e9bfd834c5070c310c50b894ee005f5ab3f44ea261842d5d0030e92696bc9b4d9207fbfe18799da8cb522f277b44919b8f6e83e8bf2f263cf0c3c2e1d9ce67c9bdac5da8302c94eecf63bb8aa5ff0e79a8e327aa3db94fd358eaf2cefd1c06991b3ca1cdde94272e58edca2a1efd558ff0d28adf596464485e14a43c7d1740e41377fc4bee8e641c11404c1a29a5f12e883ce9e65ddf4dd03a9e8146f93d6a08d7c14e7ba2c5e6b80986e29f431491073ce83e9f5367d1df50501b2bf00d69ad368b42692e05e456e04a841e7b279d851254f5e282620fda89e284732a039c37a9619c206611563b0af7f2c4e6c083f311a3b0cdebceaa3a1d13a93452f7b45d98579cfb5cc4882dc43d09a01da3ab7329a264e4ee25382651b27c712fd8f9cfdbf94c70be42a38d9ded2dd773b40a282df249f8bfb14cf11c958445392bda1fc1088693d62441b2bb8ac631c1f542f607a851ba5c087b683df4b1bf238dbd2d816105397bd0523095916a51b1f69134c11547aa8556890e1d2e2acd956c342edadd40960864b0793c9db3c08cc02b4faab2b0007170613721426a5a26f6a388e9222ca0229af327aea5bef28823f586006c40731c5d22daa7bcb4f7cee241b097c66e9fbbfbce9310eb47b04d44e4cc77652e0cdabf58fbb46c52033c0f49a7ab751db50473c2e5d5df4bbb0bd8e1920cba674d68ccf4694f1c69cfe044e71abf5b3012bab1570818864d794c2ca9083566d7180b3daf4a867910b2830e2962249120d652c1395df965c51e025cd797ea9707ff97ea3131ef4f0fe89abcc4452fccc3ac902e2e8159747f865a048896139207203861bfa0e5cb3e7f305d8ff002f2cd725ac2a656477a9d315228d4e3ee09e89c8f6f36882f241bdafaff17bd9359c2cfe40902253041d90ca550be2bd0ef416f79dedf375073c6215777f33bcedbc704c3eecdccbaccdb03f1e8c8097e90ebfbbf2e7b41e907962b917892b7d62479c7caa402d7026a8dca0d695007d0370c7c7bdf80f39f59baf5761062f1aa496109305799e69b32cdd3c0e87bf032022382952959a3b5a1e2f1c53432db168915f233851d2f5a8949eb19694e38349fc2b4507558dc824d48a795461e8e36010649061f1793d6b7c01a5bfb95d79694ca69846d40dc1500736a331fe74294eae303744264e6ee0d3528b38f0a717aa64c08be18bfba250965d9bee386ae43ce4efb720c146640c0975383e0e5f421bc25b3c0e2f1d5253d6747b8ebc7b429a9b6abac520c033dbda076dcce46e649ef933fd1b8d53d89f9708f46716b668;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha8182be62945266e738ee5faa983148de787aac2649296683dbe96c546e87608d1b2fe5e34e72163176df1e7c438bce293ce2d5e6ac0ad806f67929dd5a5a68057f5c97e3c1284c4284f89c4fab5b692dca0942bbfa944d247f93af7c300dbeae2ff52c8a2e0cc069fe9bd0013f5f240937b29a632a7aea3d1ee1b078207a69b95c586118ab0ba75bc2986cebb484b4d717367cba4c6bf4506a2a22d4e1039fa837576ca709d2376a35cd2b0bd7c8d89243a91a3150324c1c0883a09e7f1a18cbde7221bfad6aa89fee5aa5e0441f4bba36b8781f916b48675256b3815da88d3c09dda6d957bde69ca06a37a5d140a6963674665f4653af55a2736ae7e3d5f063cd2aec0e6b933e281d75fe1dc57de578442da2dd7ad250ad892751e35fc0b85d536478d8d4741ca5c38d67a0df8275f6124f1f7019d6105ca4f1c09221340bf86edc7b36b6f7d9792cce8c2ae5e8cfc195ee4cbfc4110a05acb2bc6cfb5a9af3916fa8ed0e26c60b2a7bc9cb47bc6949634317edb9f02565ffdc8f219570c9419c9b2c97d4a0a842b09d2193d3087aecef862fb90dfa47677ee65d1824c2ce3925f4007cafd08b0187e87e62f8c35eb222474c0bbc2fb4e7882c88eb560602bb9c1628e685921ee499875a1956c8ff2cd96a0c55ffca42f5524fd77114619bd8ae6195fca7691f7c01b43843329f591f667a73c767461e984c4d2ba06a8b44ed7c20a4d92cbc239ee771d099fdbe3047b8eb11999cd81bb3fb75305533e52ce47a3022cb90707e4eecf28e5f7fc60b690adc0eda582777e390197097adbe845b81ceb3cc0163ab164ed193abc46362783949247736912d04a1378b394ccb9732ecf15b7288ce363fd9e5aad619965580bf3f84e0884ee100206d09b20554a2b2e094f9e5455e10cbd64baf9ccb9e6bc7cd6b12c2830706971f0230bf1f02de94033725e38ef7523dda442a4bffb2d977247256f4d922f872faadbeb50a0bf201132414437649f345411a788a4d5713ae17bce3d7a576a385e637d6ca691b7c90c77fd311245391bc21b61569382009cda6c643c8c5fc7c5e8436f6a709cf9d5acd0d99263a779775bb407af2233be9d17da4858d1c4e17ff9b5d27a5c08747afe93790355d64b9bddd7c6e9b78519fb0a31456d0081458279fa347ef67bf92abca3032d1293d75dd4b246085a3d0191f111c7dfe2cc1afd9fd897d6c03c6456eebf96710775080f29079463eead89a898394be8f9dce86dd285c4abe9e5c682f8818bd917708f97f83cde9e732ddb336b297dd15f027b77f36b80198e296c1f4a8d112d4559b7bd61663862a504646c45b488b2ad29c5f43bdfff1c28c69b2570a3eb1d2636468766feab2fe3073ba8840030e83dafcbe192d00eda6496ed616fb8b44e8ade8532dd757b4738c592aabd64c1291d4a680e1f706f411c262a122119b89f442364a644eadcd91a7932aca2c21b650db2f2d5ff8b30d5c56cfba287047f044c2fd37d6fa0ab28c75424be94ff4bc98b8cd04e2df9f81e2a5cace72913ca8faf1ac648024e553f2035ea56da773d75dabd6c556ccaa05c207749f1f10d8c1de0de3d654e0d2603a57f605956f507109c6a35e58cdcfdda8604d3c65fe2d90ae64703f8737d061c6c04baa7bfbe8f6740a55df0df8ee6b12fda630618d58fe075599065c893e45034cdeb12380ad21106e84c8160e864bff612601e25d126c36f7f4f0f66c2ca5e7e64cb9df21aa8ac08f6ca079e3929334d0f5fb9dcae2c2b479f048b5f710256982e7a5d00ed0ba62e11e10957fad09ec3e1574332aeded515514c43dac12e9da865228865de507523aba096056408866a5504f1ecc88fa8748807bb0d1f616a41fb0a63f567a08df53ab0e34b133aa6e29c9d8dda94221f7c41e4459d60ebf6e852969c1e8e41b2fd998b84f9870ea3cbf171f5d01a0cb6aaaba6a30de03f55ecdf03258eede1578dbe5c084c8f5cf181d0c1e89e6126d96b0a75ebd8c2b283f825eeb933b98d1113cf4ed3f43e6e053fcdbb6f2ecb1613f440ef426219a1bb88b6ca96d51a1c1e542535381a0104198af4010a718c6760ef870c30ac38a91afbbe0229d34766514a594a84c3ded3e525ca4f80b1d0336e588658f8c25261af38d00d31986dab3421520a0c8f0a1011941c3c9806b170524ef2309b40551c5e3694606b66b6ee2349454a2b73ca66b83468ca3d06cc583a4c22973c0f16a5569427fd00ae576af7725af985aa7331765925f1f6171f0c77338f0d9d7edf4283c14372ddd40d1fc13dff85b4846d60db5f977560e178a51e48ebf96a5438e2f50cdd75c188dc6abefa85b6a940fee9979cd214d8db316ab67d3d51d0f085741410fc9d5e77cada2bb2415aa7ad142a51c28eefb48f70a8712029d97519487d272090a6f53900a5e6e8bd14ab41f3bdd98d86dae0bc203bbb2755876006a899310e3498cb8037bc845a9a292b7dda56241d14eef85eb2d9ad0d28d0519eec88a80a50b3360d71941231571ae6e964ac30a7fb7f5872694e7d168c92901ec6c211b9e83066b9af5586505c4bd673983c4fcf89ac6962a6b6db605d560e7b5d818870d784210dcdd7f24732f33aac8c99b00478ae62128b17bc1d6c4a169ead32c32bc2e50e53832071951e24fdcae2df332fbd5b596c4e2f851897e2ccd0e755322be58c7222c14452aee200734ecdae5619e7ea42c960dc17f52814099be4c45eebfbf1e0cf699f04a415a985;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9e83c78229b5dbfe34bc2450314c12c48d90a1fb6791df6d25d9d45a4d522d38b36fd4cda49f3ed2698d8d3494d70e6421bad6337996d6961249df86da019495f0881601e2e84ff8c41e28d0f695f9626c18a43bc1dfaa44d5b0205e8ffac0353fee5c1fe08d8be76491448c5bd4a51201af7416a6d9c20948cfb80ba6a1314a027ce624d99de373f0676dc9f6bf5dfe890796855302bcc36a72d5e698ab9cd7f0664c6004e2eb94ae5cff6745cd6d211017fa1ac5554007eb02716b7f5c47d8492ef14f986ef590cbdba1da05614c2c11bd197c4212129adbb509678a295be9c1fa6a3efbb0b678f71f1783495ce72681cc469b42ccef1347f4200a9fcaf081c2668a713f81536df2b38ff960d5b0ee86a6564fa5b84b78d0147d6b049ff03c4a3446db0caefbcdcd2cf747ff347b8c0a3720c843711adff53f41934992356a0801094e29f26d50f5f8e94a12d6ceae2c22b3033ebc7fcade81b7f62e6a9586d065350e283b71173065fc8683efe3a1064a44f6f0ac12b503a59fa17add6675fb59825b08c88273571dbae4ad54469ec9461dcb7619f06b9d27c07b629551e89626bfd638055085b7488b15641fc2cb247bd8103e7ece66146d82faeb06af3cc3f051dbe20152fbf510bda08a8da3ed8b58e1116d2808d6b40057df9732c72f1d37f12c5105d03276c04ed04b7c5e27fdb781775af63086b494da44c8b95c71649ffc461d7b1b17ddbdcd3a6b377a384ff5d80c261d32b266e90d239462f57b26133033f5108fc29ad09fc88677bbff4b85e5abfb07bd7c395a9e84adb27e3bb0a36114a8ff6960301296843b3eb0e6747b39dd100d725b31ebf7af1dbeb998e3d19cdf23f7e0abf89e627b102da79f9124339b360b0fa1b9d853e59506f10c7bb42691ad6bffe73a0d3f996b7436b61f8b16868a9d31353ebcd9e0e0bd1cbb363680b0458facbd4c965bb3a8731e277b6cdb2c76bd115a66d02baaf74b7e2daebe5a155a370c8f0f585194c5a3c2909fc60c13987cd7d557199ad9ba188a2d79dd575fa5b870df5cbf215d270dd4a237e516417483fb2c290e4a7f2e807f135201ef9ddc7b37a640d1761cdbd8d67dd9df4f2b1fc84e2435b076ce59e2d2e0587ef5566160c10b50de34b2401b7d4e1472bdd7285dd8053e840318ba480b414f32f99aa55027de0233cb9ca503aa45ec5a41429b43745e4dbc4ff405710620ef51eeee8151715f547418b973d34c664ec41ee43b3c44ab864951cdffc60b5e4f25dd88b2e6adb2213b6d1cf974f3d4f50ae40a028120bd992fb37178188a331f183e89176364101a740a01e39a1be4d42b0aa548eb252dfc33554603bf7a2a16684aecae87686e4c4def26b76c89fa7e0b992966ae97504099f2b7c8b889831dbbc705844758aea11ab25bbdf7db9706836c28df3348b4615bf0b1daede4c363c2f73df9ff237580eba01bb0b96f3c6e743705bc8c1555f4d2e411ad44aba39eb65c56d7986795624e62a38d6731a4adc644a2e1dac1892a732e402642347e5e58009bef0b2d5aa0278670c6a624bb44a1e9af7aed84364d255103956dcd9255f1d18b7adf0249afb489be4fd319679a11ae1631857e042e6ed4eb0055fce3b2c02d5e6549fb6ec6d28b7bbfd63f8e321693b6e4d517ae37533b82a986a637fd0f424d736b40b469272408d9f6d5696e7b56c49fe4936734678757e07e761e9ac1f95dde64ce1c0917ee6e4e81bb813ea94da61f06c12d526ff2080555762d7ab9d40f69b362bfc9ce4ed21b298161016edbee456795ce6aea9355f4057a61284dca5ffbda6f1f2661469912f98d3d15b39bd1bf7abc208cdd012ae844d9ed6ec22c820c8f916db9c4bfffae4df25f645bf5decba3e967859bd617a5dc5dc4dcfee14a0f4688874af4ec62c9366cba7678b02e58fc345617a94e2915dcad88c31241f6e58f72b2b6f7bd131abf3ce2206aca7729676708e093370cb2ec0b42f3b32e4ba88e3719f1112b2757b11be62499e8d482ea67c630c51eb169fa8e3d69ca5151a8ba4a4e28f7402fff42f6c2c85697d4ad56d1ff3a968463b393f3135b3f048f79d48a90c720bd694a4892011bcbc6cdd0bb81270b5259fee1bf49f3a9429dfe689697c6b3420f8dab790045ffd1a79f4942d3ad27e146762af4b86243f83538a9e36bc26bd213889dd98ea0da2e9d26c4f9f61ef832c93714605eb5153089ca13fbedb37b52700d0db95448e99419d38236786ceeefb1cb8189a700f33858a605746c14de2aee88daf4dfce1779cc6a0798b9e1edf426673e97e4c93df0dff92ec36b565c0b99fdbc7f1288f2c07103df5371b97119412fa7d8564f5d6eed20c4d3202787a9c36baf39ae1e4a8ece5ea440022717259845f1642ba62b4999dbe964180304c4dfbcddd727a800f884ceb2b296b7823feeca302e66c13a56eb3f2f287adb7eb0fbbbbe89f5ac76bff561a247019e4daa08e6f3259eeb6b570e28431d9f35ba9c3c155c7932c40c560dca8246b6e5b25a6d152c559b7f3241ebe44c860a7b2e35c06cbfe227297e2536627c08cb8eca6e52c6c19e7cca9f106ec8030310f6aa9037c35b9c72e9910c8a2388456a878ab62e4cee288d65aa99b5384ebf99a54fbe76d3bace2ac877e5b8534aa0aac05f1dd324b9d9d2c3171c4b5975f0b2c48f46043ac311e0995de71695e6f5c00c47d6a278e58e9be5f0cff3f65c6cd259e4b8e105d196b72c1f4355c05cacc083;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2b03b70f3700e6f244a0c3a554c12317da90b05230a139a7fd28e18885e53309770069bf8eff1f9a2a42f704415650cf1aefddb402e9234395caf2246ee5e0b59d648116d1772e08d209aeca6d57c20b4e74e678c0338f0a2d7057c103979d0c04072e3d9a43a98acc9c07f3b87323c14a61a95ecfe5074e8f510e635e171d97019dfabd76ed3aba96357fcf3052e9b2764d227da89a39822287553a549595d16db258fc9288512a88788f3711c981ae4e3e37930a0543e15e73a118133cf313ecce2f6f4895df2ec5133432f65663a00e0f2182942d4d117b13072201e3f92a0fc68a73e4525e08ae2f89426987ca80f8bab7a8ffecf979a16735655d084afd15126863b83b7c412cf3159e97594cff81b0641ae11265bf030eddd71a72b4331c0b5f363f8ec993213abf1cb8951842feae58ce0cb66415939b8853bba05a1afb4316d12b69305417e8637a86a880549a5021500562e2d972457609f85bcb0bde52aaff12d6deec71d1d49cd5d62429b7aa51be8c543b2103ca7606abe80c2db213e3f363f69a1696b6e761bcf13ae0cdaedc4fae2ad4c19e64c23de407f69b10d615cea0d162e9be27ca77a7e97dab05f4db0d9b98ad68b237a1909270880597381944eb9d9c62e6023280d3fea37903a0b363a958cbeb9308bc1b9e8e974aaafed060b1d1dd503635c66453a054483f83620b1b04526ac9c14eb412d139e3e34e63874b96255676ab8078cd07c0fbda29cd69e3a4b56f3fafeddc58222ee6d2f2d5bc0616eb4f4cf44712410df397e6204fb348210df55686d701fdc6740b1cbe0bd8ca7807e604256b3d523ae4e45473a6fd33e723f7caf4aec7da65aeb5a98d63558f62813ab6f9858856e5754d11d72c043d10f67c0cd9983bc03c202e2df3a6a9d0e6f845b913e03bc16b61a313281bf99c7ccb3193d5fbe1473b49f9a1fa9460b9f07c54117d02bb79418e6f2b3407280fefcf313c32c9ad35ec5a161fc511b5903f0934279323068bd0ca43bca5f258b77e5401e3ffcea7ba8762a3f428c8f280511461a3c1122ae7034602c2fadc31321cafdc3ab54c8d40e84c9043500db09c7801964af7fbd850eb2a3215d24ff0741cbcae437572c7482359e1fc7342830d48f7bbe2bb00727e958a598c47ae5918ff0a470e834bf0aadcc9785bd911f02658065ad9cb438a8814be6d0a8163ab18c9e2a61e17b52c5278abcb8b6c4da94b8edd0120671ff0f167835d6633e62e760dfaa40c813422910e740199f7c0498f44bcab8b09b5aea19b42728d9cfd43fd01658f3f7a033ba94d9b7cb0e528280e733ab8a3e69d6835a5f24468c99d661fd094d7b44dd63c0c2b4af6564ee38d590af68231965f8f6e481857c23140621728be2327c6dad16a7cb2d7868c7328b067af555907f331c7b7a967e55bee7674912d942967163865dcbf6742bfb72ffb7014bac1a4da1c69b9f4595b2dd49ec5021e47c1c6bc8801d6c0c97c14aef3b9bc3c7fb2d2fb201e5c43b2ec9fae182a5ca0e6839ac7363103e0927c0e4b9a7bc2647ec6e6d23711dc436c599bde124b9b191185231f40674bca65a0a398be90bfef63e5191de9ee836133f0470b1ecf633680e2a72726cd37ed4eae1be0b242f27e2eff89f06bdc5c6cba6d073e076c41937e840acb41eb6b97bfe47e8ca83e6c4804a5e4fb133c15f1adce124796f571d948bb91611ac108e7d47bae22164e68895a6d55762491446acca5fc7c68f824bae687a1b13be5305ddb660f1e468a1cc841262a74d4d2e673ff2fe3bdfc015870bf773696a36e45fc9138c574b7124bfcb569efe7c48f14b84037bce9698d2a442f12c0ecd40b793b738cb068b358ac2b671f27a5e9be87b84a6daacce390005327d5606418d454114240be4df665a8c5a7ab087ec7f1c2bf5dbff736adbda27e66f588c9e8c8663e21f6768fcbfdb0e6be1ebad9c85c4aa6c51b60fa769d529bec8b59293e4b8b9b81c393faa2c77cb9561ec2452b7ccb1994d87a5a9406a2543f76e1e6a5f5e790932a930173ededfa3cd46239bbf1d6f0c0bc88024074a38c3aa007490d6b43b18e788b0a1cbc7de2589283eecd71caa376269f1b108b855cda1e3d2a9cd61190538b4e71da0f12266cc5b759bf6ef3b6ea09faf4ba041f6ee95e2d460579f8f687464bccda17a31f075267d0a1cd7eac4bd16a4af276c86246133f8a177050e1a03006158af3af185e6dfaa3edd15e879582e4dd77bbc5d63b1a2e982fd019fc8ec543138d7ff852c443f290d14254b8eb370eb1a83dd99f354bbd485d6952ac25e210a51f24979afc503f9c28714f7b8968c5e661250d66eafa0737a16274c5032e7add2e2fe4ff709704479f54120dfee160cf94697d9993eb20fade5b1534cf8c144e32aebc3aa2e24818e793bd2f4e9de6c2efe495e0ba355e1af24de5d24e9863efcbf045511ea25d56cd8dc0672cf20f54ad753cddf0b41afaa11afb0b29d7de95cd8c37a526f1d443360cc6f9a6f5e868f7746378e727b23fad6765d6f0c1bc2c794e87d53c6410dddca7c43001297a0144c6b2b84bccc65bd6d0fa9a0518507b4581b38b0ce9e7fac813e31d737ea9b28090e64df66b89a55fe309409d7827973c8ea998ce489bb66d60b5b1cc3b9eb163281eff0f9e1bef63487d45bc6c7e261124729ea7bd18b31e829b781b55d0ea051cf5c1b921369bbced28b39d47b1afa223943d307eeaca1bd9eae52cf7bbe6b0d882d562;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbc3da013dc2c92677109bd0a5a3f679c0cfe3bc8432b615ed60a7f2a1533c2ba04e499924bcbfb1a832048222db7ea5ce5b37217abf3a15594f3c9103b1b6f9905081b4142122ddd630f161e4e66b707439b1692bea841301c844750145c22e7f60d3035f657d6507a5cc9bbc62d761d41fec752743559a29dd0dc347ff0230600da2139c0d2a38846b85942b4f17c3c2fe9736227a9ddd7358a39e03b9feb85dbd4225188b4cafa8c504a2197452007c33785d7b7f9b593e5f2bd4c8e286ac74329ff1e7b05f5dcfb5d72fba774652d6c136bdbca287013fd0c86183826a5a72fcbf154c6b227327da3782fdf8ef9b8bc64624a322af483534cfc2f98540e25dfb2de289b887c0ebc8ddd0aea6495b7c84ccc4a9253316fa12c5c80ed5f380f82c55568307184fd3302d22b47131d833bc44d2a91c35ef2a7fa87165ad8c5b92e68eff4909991c4bfc2de706cd57ee88282b359eaf9896759fb436ba9d788177d7168ec9379ff6c28f237ec6972f0650ff9ced0a5675690f416bc4c1040912af97509af4209e36bc75bcd7f385ec1b40644a2b46684d55c30284114f6960ee37df85fee69c5e9ae59856ea9baa934680ba25669765bf5090b1043715fb2701847f338dc121fbfd869254c3dccf6acc0396e5d9e5f976ade5333dbde546a0a1a249c73d18f14df7b7a92ada686bedd8ef50cb54d1c5b85330e85280db01c8b8db457bd3de19de5d0c788ce0536f6000ca80ae6917c0ddfe3b4d5489efbe2369caf47f034f288c5e6520a4a8ceb5e95de6eaa77d34fb361a196c5195b074986492aaaa31f963b6d702acfe813c838a4bcb78740877f90e470d288747065a47ee248f274adbe6098733d07854ce2f4c4806b34e109fcb65cf4c5ffaeb9bf6675036b79ee8f6c609470ae8b4f7c24dcf6279336fc77aa0d91c37adf85c0738f544ea4c61b52982b093bc4948b6b3eb81b1c53e012182c141fc0bf1b18045fb17016b510c5ac79c4f28b806f76f848dabf34fd81a23e65881b7fe3a19c6247bd421cbc7cb7bca1e05c6b4e071f15cd8c47954d1d866b9c31586eebed2b714c32c3f281f721f7ade416f4669ed7f49106d1189fb894f57b9e3416f3251d74ba3d1ecf0f2df09eaca2a85a13add1efec29a48b2f3b1ba6238434da04d925667dc2289cfb4ac6dc0e8c5534aa77230bb907f946abc59eaf54dad745adbdbb20dc8f8cadc6abebc90661d21c37d5e91898b34f35c6f4f9affef30e76fa98d2f44efb5e1b91c92daf14f2b6797d57d341436b7a0f9ae5c630573ab751652339f89a3ddcece3834e83045ed7a686069f4a2ec35de9e56c4346e3ba3d575352955095953ae78bcb7f5ceeef852a4702b589190e2012077355742314df83743134e82179731b2089836d544c2cedc9cde09a47739fc0579b851dba32235fe5bb5f0d6d3caf3b337837e670054dcb89aa9f4bcec0493023a56f08473fe3515b2ca2143ecffdd00103d7d1690b45d00b60b54cb5a876a5eb7d28558c6be7de8bfa5eb323432f32a5362d06a826945cfd2e05ce62a624c829384629905c149f371f8e5617b502b589c590cc37461d9a70a7641bb36081cc07be243500e43fc5ab797b8159b98a367024fc94063d89b7a8682ad75d7c0594f0abd1bb5f6f4c9c91a4e9f0b3c5440cc1aabfad4764007330f7fa0ba3ff4a6c77f936b02e43138770ac93113d53498381a28da0f07143e07a44323d4d809c37599cbcf439cef90eeac5c1ee1c5103bcd609c941f1fbb26a3c8895e106a85d49ebbdf260c65f9ef1deb7b8d7a59b5713ef032de7e200a6fbfa9f1aca761b8c3cf8bb185585bb16061baf5f9eb09acce0dd1cdaeb7ffa13fede24dd31a6bdc2f97d5779a31731f9381d339865954c256c715a2434c7dc849bf9a61db980cd2096cc1acdb63412f5c8f8f74d05d3e411e585743d77e18d944845378c0c04c41d4ea5e7d974ce6fc8e3ed0d1db93b2087e5d701c1a663e06968e472d3c8839740fffa4fee2caa6cdbb6b8d128d7c02f8e8e05827db1af0b9cc8e0adf2a697fcd016ab151a0fc9b07c2543f4f8b9a74f69d92b0e75fc60496eb53aa6f860d8b9b7191f482ec3452a687d0410eb7671758b7c193afe3f2eaf503751ddbc3d52d70ff7fa604ff3da4ece537fe18753bc7e17f850fdaa511410df2341ff301e0e14358679bc22414a96d287f7dc15b32ce3ed0b601781068f7862d6cbd1a15b3229e89ecc92b43ce8a79fd661252ef56653503f4a4f5de1248fe248635c48a6b9be14257a89b6bb5f32ff49f2e736d10e4e91868883d540894e4fa7a3381df4c4e2e0119db153e5872f9e400692ac9967150a6390bac4f7a5b655d567a51c819b4f921f5a26b1eb26a51eea368d6bcfc8fdaaa0b54880b90d128f10c742267bfe5b63262cfa222328bf0120e7718e8b4846dad10e84569d49c2b9ac4c772eedaf0b4a2e5d1a59b84046ba7d4b781dbb80a116e8ae724efafebc875d90b023d3c006cb88a6ddbe37d5d7215c6227db430eb40833995f78965358b503ed450dc881f02cc3c965107f5084d6a4ab1f2b08db744d2c8d8f0df549b1c35a1d737d105a03e77cce94a73e55ec77c6af8d633823c6f677fd3ea92b74126ec948d88a9faeec3fd1a8493b1ee33f1c6f5990b31e93073a0bc4f0280d81d9159c0f93109daf161e2e79e166789ed5ce09d763b14e9f137522caeea8db71ba8961d48c47c4260eabf71277ca4d3499e88e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbf772925340adcebf2b0b17503c261eeb153dd0c730bc08edbea0ac16434c9beb267a7216bb7c8dcb425553f8734f3e41e82dd0997deeae185c3fd3a7949fd379a4472d6f67ca7d2c09243b852a9e37ca76d682aea979f9698d4e8d5d639210c8f33641834b5689130dbebeced5b5e278ad2b9b64b2d0492d7385a36971767a09c10da0e1e098e086f6f9e4ae55ae3697f48f197d52641ba718f22b7257dd4f591dc7a00b49f60ebf0137a8d102b3ca666b1df4d8cbcd8f420b79cdb8f49d100b301b08425073130b93fbdbabf927bfc5fb5934b724578963dbaa394f264ec2a6b1f5fe891691abac0514b6238c3e730310b3a528d272c49de7cc229ff6f352dbdcd6026fbd86ff29fb3cf11eb03a962ba7ead0a16627340f6bd9d63564dee553c1ba62ee5184172ae74a4b854334cd4d8b8b5139f98525c5704005d6f57362c53f04ee00e9b61239b6bf4ed0d1eec7fa8fb03432517ce58ec798abc50d1e6c5ec943db01b70071a9ec25b829873c754f336edf90be2a94375fb2cbfc61e9ad5b3b75fcb7eb1bc5e9dbcc90a4fb91a78d9c646bb3481a8da6ded49d184040329b16f51e704f5aeb81769b8b183d03d144a82e284700b11d3b10e2b70c4086e03725a487cdd6631767ceae4f6b51156f61fc2d6ac150a20cd8daaaeafd3a1401cf81016c1728888de091d794a0ead751706dbfbf98c1507e4986467b53e97e886e2fe1a293809de8c915b7de441204e8f2eb8d1cfa7aaa967d746af6afdb5b0c4bc3b9171f7376c986254f0593875dbc05d4590d2c1b56fae924fe2c5a0c7307910457d059c6fb15c9a2a02e4605810c9e731d7b3c0562ed1db4e684976329d5aa7b54b72969e26380108c068f00ca4da00a82402ba231df18fb49a63687c2e44445cf661a1292398259db81603d9d0ddebeec5f2293b979fc6ca4432e056d3137379a19a4677a45ab38ebc5697632a0885af74d3a8b9938529f6b5ddbc9d64eb70397372590ecabd67bf81e102baf8a12fd3e2b01310a6a732a6a26996c3af04f872ca994d6e582191858d81a129162a2d1cc4fdb353ffbc83944d6a61d36dcc8dd66df6ae8cf3f2a1411103f01353f31ab85f4869befed38f1f7bad9d7b57bc6c64b554f6ef2de32a732f585e8a0ae3cc2674495dc93c4a531795e3490efeff86adf9308d1ff92970f7c28cc0aefd3c759aefe27087f193c6bb429d020b1c8d461f2a3ea1c8ce15a5041de1cf72d06a28071d9850e9cab85a0379b660095357a819f3d521a5af0b2d2621cc9b6700826c5de7025eeb504b20cc5632ee1068e6d068cbf7a089dd7e40da0fe5d940897cfcaa02cf01b7b43e909dadfee7f87774a669b80f6d1e471443947f19498eb46a1e325d361227f87818c0f0594cdd5b576217ff196aef1930fcc77144f35cb5588be83d226d0dcd8bed586c6432acf56dcf1c001f63a918162034c307c360189d646b347c04dee8cee44442eb013c628156c45758319d54664241f599abaa4ee3ea199f7e69f722c2e1ace164bdc895897197a014a93c04af287269bf464168a37c8117410d568fb5405d062e5d8ec7b5d675ee042b29a5dfdeaf5f371b4089d3b181c38fa1a814c7a17174de36442cb5463d8f22c6ae3e7c6b9b6d1d076dff7451e94d2996f16a10a71b2d4cf1526ee97d09f4811e12039fa1f838b774c51027b99617c20686ff7532cb3c725542b0902cab58ed6e8f21d3e9649e100b2e49c63f1e396a65f5c7c8ba5069ac1a32db3eee8b330af4f991cf70fcb4fe9ded277078e4860059e666278b90c7b0a971adc4da1c53dc16a1da99d5604da037fc81b83ab88e748373e3ff344c623af5185885356cf237719bd6f3c8fd59c706b402e2ea6f39d43a818df77ab4e78134bde6568551143bc1e6ebd98d819d5df0378d434c1b0e6f4578aa7a565d582b0e841a2bbf3c91d125bbc6a994dab83c871925de412fc17fd847c6db39e2b38f114ed2c8be0c2b968b3df1264d331ac999382b88abd0f423271c1511fa0a234f962088dcc01fc99dd20660c89e439dfacf1f63484dcd142e1733156a6c442733aa58b74429850346291fe1ff86bb3072ffc12610d85fa23957f95d61d95938c56e9e3a4b0e517d9b5d3074ec5474971b7d741d03c90ed155a6e541b9dea63c3a5e9b37f09026ec68b3cc989ca06c4b29dc934b9fbd42bf98f6050c29cd327e53aa04a6971f79e930528dabc14a318287c2e3ce4c98af398b0f3d7f6ee02ab6970f21b07a451bd41dfc56652a5d340cd31d8774a9db296f732eda784428edc289cd2f9590ffdd1be33673ac501a674134061b21a0dfef808065bc8673834ae8960b23e6db01b4979fcb872dd0e3476532f4299db990869761f84e6cf46e4cdf5c5211537464b56d0505aa4e90839b512ca97c3196bcac3471d37aa6d286e8e707a3351a65755c8962fb6a3e74fc584880cc5ca958df05782a6183db8d4127a4ab0ae64a381e5cf9b63c18e68bda151e45fb4cd4afa7e143cf8afd3d170234523a638d312412e292550ba6e5ada425c946d9f63221f4a36dcb677af85cd46a5db97593502fe9d31b0118e464815d2d0e3272488a7202da71ed8af8d9c1a54c36d075d6ca913dfa8490049638cd68d78eb02fb02e45aca4b1c1078482224c5a3dba3ba3bff2bc949e1a09eeae7730efe205dac902f29e1c8a0289f6169cb4c9228a52de7a6d7b63f4439314f34e76f9460a9463cf1017ec0ee967a8dcb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he10135d64c9ca05dec937485e7b92235aa4af08847d805d929d3034fe318e65221493533db596f750ed0d20e474ff7ca7827e5078ecb435a014508e862c7c0e1775588cca427ff5ffdd0596fb2da3c28ff9abe7d62000a4ea96052b78c61d7e1d3a123387d8acc12e65450a2735f4219a4cd945a6cd4c7ca6e699da2162368ad8d15595b42c6e1bb827e8c86cac3db00fd1219cbf0970576fe3a7f2bd1ab959904e3b10e72676bb9badc938cf13727e7ec7c3a200dae0a265cac8acf313b3bcfc9b7abc7a5679ac05e6d9875c669473d088affe04026d25f50e97cd24d8a5477843534c6774467f96f9000152378da57e42b6f39404954281020c1adb946e262cb1442126ae2a4280b3fb8fa381185ec92bc37bcd5fa33c57fdb5ca6f5ead103dd50357b7b35b8ce1b632004b751023e9d89f98f8f9bb95da6df1bd9dcbf91fb35bcb4c1a88f7b99c74d2ecaba4fa80f4f6ab9ba36497c68ac68ffa5f7532fbc9991d9229c4a78029c812c8b72bffcde653b91fc106088ac7331e61281198f7087252d46e8d5fd1f2775459e9dd40db9890e6982e794db9759edb054a199a237d2f6f0102696af23188a819b09d33bf913d4152a0722e08bebfc3d94e9bde7c8bfcc086ef1e7af8373759a57f6a6bc55758685d27e3e4a1cb067281ce059b94eea860f184acef503534696e44f5ec9d69a58af40a0d6d6826d1cc6b99ce2cf2e8c94d8a5f69484149021bf1bc642c310642c6316d62d25008139e592c4fdbfbe1679e7af9a04bbd42acbffc7da38edda488e97b1639ba06519dd13a4aa58c6b9ededd832ceb561cf31975fb4fd22d9c9f60e4d5e6353630dd5d300d8de3bfa6710172b1c9be498820b22e0de55e54824a48d8276fa4f73f80b22a8cea2be8cc13416bb415d2e288e0ca5369528fca25dac355fd2e2ad9280fe1219da6c453a91729b8d3581c3bb3806cc60b452deb36e2eb552a55a9cedf29909dd56311378030dd01e37d3f22e2b1dabecc9be779eb833e0bc36abd9799cdd3aa7a26ebb16cb44069930c218d0047d46d7c677e4fe2227eab2dbfb04c7ab29be8a60da3123225fa007a59fc851f0f948fbd1ded853f2ff2d119504fc0e318e498aa184b52fab0c53b6c191a65439cdea8c8de143f5645030337cb6b3e53f6ec8447892be338984e920fdfd46de1abd0603389c30d61b345198b47636065a75dcff7547f1333a846cdf092429d9fb3443a7d745021cfa24e50a36f790984d872426f9235eb6ba4fb40dc531d033875a5bb0a196d1fafdcb57838c9e734e52909c8116ff7bfafba4a4105251753a89e48743ddadfc4f234dfe7d11e868d388117b15eeb5344380360795a43273168fce6a388de49445732caa80d74165898de3d23fe235fbb8f3828dafb90068d5f0752b9559485353c8e98603dec8deb5fa97449987edbfcc1d159cc8375e51f171da8699cfce8cb4618fd65696e014175c658806ee46e15583ac51bff53d72364c8726b08664b9e9ec60fccdee648c10b2c5c1c7c8a57453cd900578d9e90ab3dea4c34473b430ad190e62431a6dc3ccfda2c334957896ca825998622bd43ddda76e13cc8f6f7fd47b624e4daa6aba67ca302b5a876dc6d26197453f75497a6bbf1f12cf8569a5963df63f75a24bc20132ad129b601da8c53dc88fae25a964ea12c3a35083c5752e0389585d9c2e477d4c5a186855de0be87b0b8e72da3aa071a64ed6017143268ffd5fda7ff2f7ae719a632061d72635bb60ccbd908bf7a911452c67aed220a31ecf869aa1ccb7d66acd8844385434689fcbb7a8ee5a36b47e6a3f3ba5b5e1b042f348bcbe3bc9d343832de3a67d41de9264f9fdb3be1273625f596303778ccb0cac035d6bab54f2bd0e8e1b89701b58991966bb9ff9a4a2afc7a89d8fd9133577f78692e7c0a66aa10e74c3b6fd0eef8d7be3166713808568ea38f4788f9395bc0fd7fade7ed8afc5f16d7c44b7eb1fc15cd271abb6cf768422efab29c06fe468be99611033c6f9b52a260fa22dd697cd37597a91d0e96f5695ad3e45a497413e81521b75ced319c6dc8c49be4b08b145d1789bbd738620602400d0454d18047d414cfceeb16fca9625054155243145ec2c9e754e74768a5acd4d209b0ebfdde9d27b12c4271f32ba2abba1b3f7098fe44e24ad14bae8c71c9f05ef6e13fed5868f6424e3d3545113b8f4245d033245ee14264f0c8a2ce07f94d2b46fc7ff25ab004e016d44fc7044f4c698d5250ddd40473e8d6dfdca29ebc9c9cd849a19a3e92ab50818e362818b5379ecae628819938156ff1bfc864649c0f8ea20f29881ac409908719d9be9e512c3d03f2b15027f3e376cb53040c63a785ede63d8167728f96db6c1c8e2765b81762edcc7b1d7f87b3812872535b8de6acb9ab4bf5897f2a6c891faed561ea8c08799cba6f2e1b58190950e22aecb0d7b478369747d3dd39474b14ed140a8bff181da2e1d5ec4d8da1dfd235fd8abf9cd30ae255a7bced372765d22fdfddb6cb5fe9f5ed88747918c06ac69abceb1285463829f7d5e8972964e50c273400c71e29697f6c2caa72b235a5a8a556b6a6be97977d5c42c1956ebf403c77d5fb655648e49ee8d73eb39bedf5ec3eb9689ff118ddb37306f97484c6d256c2bc935c213d3f1146d04dc7a170a86993457c39022785ead4a099b9ea7c5c9f66fe397c290ad4d55f57d38637edfc0bdbacfd00ecd434bb5113c4580258024b8792f091d3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he76d5676c21606c7a85ace78e9b7fc24a26c712cc6a861be4a45b24b1fbe7c1160f10c70893971558c4300a7290b53bc4f788656d353e1b42858d1c997be3e1c126a24de4aeeb08cc9d9105eb99bb435cfc599b7e99df59ff2f5e9b695ed5af378632082149a146aa057895d4b364c84dfde6a3e26bccf45cbf92302a41e6966ef001de6c73b6ad18b047b4f57b466a8e9325b4d6f685cc5aba537f1aa3603aa0ef073ad9d0062be7d1b702baa54c042cbcaa7237b95d2a5c624c2ddc6ff1f2dab7760aa6e32a7b5980b805e11c492e92127b1b1bed4129d77a9375fe6ad995d3a1c87537fbf235baaf1e8456cc47f50ddb35a46ee578a345abd76d178a1fcf5b13879b59328501dc8d11bcca404681a642379aa395637174268117cb82a76778b5e1d43df9e1b39938a478b9c94e886b667767fbde387952d0d20c0dea52db4316ab1b9a273ecacda367e89713a57ab9e408764b3008dcaf9eb91d7a58ce0a15e22ebdf02cb4072cb841fce87dc2d350c8b99e60ad00abe04cdc6e0e22905d299a6cebc723220ee6b57022d6db798dbac238daadf95d3d632eaa249401d287e86975950a31f93e441c005dc463b87aa3dcc61812bb827f536dec42af2bd8d4815040c6b84cc6434b361c6e80d3ba6617e227b5f13b2beb6809d3f6e69fefd42019aa87f36aef640a3de65b0f8c2cc5e4b8a74d94b8983c73f2ffe04162ae45b4a9c549c94d2bd598f4f470c91cd697966ad80d4ad1f94ae260af380706b4d00202dc0f021a3f2884d2daa12d60e671e8171318a3bdef450cae4fac5488d238f59ce2666f7aa7864bf40305dad122ecd1816038b0a465ff72b2f61bfe0c6a7806470bc2a3f59d51f23f556e4e82d7e4612a4aaed07ce8bf6d04003ad57e32d1b651fc2e5f96054cf5928ee941f62eaaf82db872d096b051c8a8b7a54bd4e3e7af7fcefb3cc337c46095c89a4793faace5516350fd381a1b9d256d36736f1d0b3f8636ad71212e636f1935f7e2e70d44468b48a9a7e850bc19145ca8bbc5a0c751e9d30a794d87a726217d5624c1255f998b296510fc3b0ecf81f1d6491c1327737e260dcb66d6be354a0742f58ceb8d1f8d50ad52c735f5456e67bf9101eed971db6bd83979a8ed429175b41d1b7ad160e4203eef9819e62156c99f2194f046d29bff187a7cb73b8739d70c375e1c5c07d49be7811f53f647cafafd1cdf986b467671d9f5a7af0e458b8c316febf9cde5967b615b51bb4161745d3e5c7e5302da3cf6b92a4fcd6a9949859ca1efbf18adf5285318aba013c50a9f73eeebfefee538a09aa87e5fb4d23537e85c733b25a16901b3577aaec8c003659b9460bba263e900c42d53e1a0a40091cf8ee64384bbbc3e6d25ae322792626af8edc675f66182639e5814f76b918f5f18ee96c0e352a3f1eb850009fe3338fd567e32e300d18786255efee3451f60fe58ce1a62712866719900bfc4432c4c7b526bd1459747bb3f903e48475b5a06b54982f5b48bf1d49b0db5afcd07f7141dcaf3e0e8e64698205ec72862e10457e239a63b66ed3ed7b6b4f83664152e855104d0c1ee6c8acb1daec477531a0b57f0c8e0f4aa22ccfe8fa3429074252e04e2358328c4e8832225641b8a7180d65b433e11647bfc7f6c5e716bd7951d2e40bfc652c80adc29d5afff8c742ad3f9d6e8a3b73b57356cbcde4ba23bcf4d6ade15a44ccb028eaa937088549b970cb4390457a5176eed550dfd7da3e30cb6d64998bb3d5e1b7abc8f2c48ae9cd67b5763ffedbe18011649eb91a7d67d97c9f9ef9ddaf4ce050635be8eec68fd18fdce7bedf26566ce58ab072cd941dd9fd5c48eaa0bcb8d0063cfa2079cdce1ebbf1c278bc00d938a0cb2e59a339a6dde41d8d445ad83484da68a65e43e00f573635d6535efa3454cd376819e9787de872aefcf5919d17617a8b9e5f91feeef9c611789f198a8f9351c252962511453ba5c3e54e13ff62153f2cdb369ce9ad849c8063d98e4ebe54a57509657f1bc3cef02bfdfebdf6da490d5c0631a2eea7af33187b34ff2385717605fa401f0cfb2790a1ebb439afe14d7ba52d28d0f94f1657221d60d8413dce2d9bc1d23328cf01078836d57aee4cd710d105e50952a623c91787ec1288b34157164487d6d2b50f25ae0658ea092619a6759e5c83a743f67a5f6600401f7d77729949f9e417fd00ee352af818c7cfde820d0e8ff0a0f43c9d3ccdfb83d280c31943723a50ffaebfb8257f7f3d86370d26b72edecc5c5062a25e4835e35a2f819597d8473e0c5af804f313c619ecd81a89eefedacbd2f3c1beb09dc4e7202522cb1186137f9aef685f388a7a19ce0323799cdbf323983c0cd481214ff66214e7c594ea80363479fc985d6cf95584bb338d5b6b17c030b5cac97451d229d1a2fa43e1c2359746cd2aaee010af4e8b2150d4f87f9a50fba1397f736eb6675944cadc116f0ee64daad31305ba8c1b45a1309867ca2b9457a16d27b54a67b664b9b17185f657d73942d3ced9a8389d1909f4b0a5254aaa3865f1723509bb69fcbdb37ce752b096f59eee98d8c7c27ff4b2d7b27194142c909682de0394678f06beefc85f8a2618dfc50370ae4cdaa94bf2a48c69e0268e68b96857a97882a1bca14c34be36498679956f3df469962e18a2f9f786d7b96d8b0e13d880037b967386b8488b610a57a2cbb26d556e5c806afdf288092c08f1e7577ee40ce1e53a0cc5788de013caa53bfc8a8ac8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3b6a63b1b80129bc185bd4b77cb39bbee83eb8e00bb974b2132cf576470a89efab31fb91005c8b5e597c852951d8fde84cfc2eabbced85622468c14ec2c30fc99dccab21b72f1d3f69913fed1337deb9a108648cb81f54496e43e62ef86ee1b4b8903469807fc3e050cc57b42561b0f3c902dc6ea2449c32ce0a50786cbaf86c833290e440106830070978b9be520e63f84b3b3b2db017f699fe8491b187cd299f9a092c9d7aa8677613d0cb0896930c2b1453f2ba414778fae5673e542fcd200d5451e3de71df0bfb3d18f7bf1bb3cebd5d3f20438718e97216f00809d3503854f1a021b3b1dc7524869985cdeabf49e8a1957ba8b68b03c37431e5d830a3ab85e3afba0f34fdf1f42fe420bd8d03b19faf4336a59764a28f5d9bbcc73a76591f5b099aeda3b78194af58728b85e0181fea55af05e1c3a3a65f091b4f6ddcbc26465f3a950308ce798ecca4b01416e5f013e3a32dc27b88dcbca933933e8f5993c7a0b9ec1ecc73047c1525b1c8311a190c5d093af056f01b398480b0426ca4d337590a49ecf2d2956e77436fce4681007728c4c40781f694e8c88236668ab58698bfdc6ed782307dcd5635e5e1825017af7a75b06ab7f2f641fb2dcbab571823d5fa5bdb2a3c038481971fc8a02a277cc1c32ccc62b01ad8ef8ca9fa225a69dec4caea7298e924fb192057f852a176d48cb6fe3e1c3ff94807c05ee5cc5b7003bef549dee9b644b5bb94f51f7515e10f80a0a7bc5188d46e81328b90410702ec715b1bed32634964dc3a090b47ad7e9e59d88b08099b94ae0976abdd06121543413a4ec0f9b2ae7c429cf7accc4520c113aa6c22b9ec4fd57c66e2ad6e943625e2147cc0826b3d9003f8eff9dac75e27883338f40afc9014bcb2692c1a04d8619eaec32b1f14ae2f5ca927e47b0aa5ea35b090e14efd722a23a8250a161721bf08f2d8b0f24ee4cc4133d88e71852264fd8b93329fa398a26492492a5205983490abe333be75e1e8b009960f5cd484c598f6e92f2440e5e4326de96d118324e6d74c2eb0d35f2f44260122e24b12d44c87f7bf27f6da8b3d66578c90e819512b443f4e8ebd46c616767578d97a1394b55db60670393e95837ce58cbfe11373c43e06b24be70d013e4271c18f32f9720f1ddf7cfd7d0e15b45300e6fae02755a944dd7ad96164e9fadb49063fa6085077db7afb6bec8237c0c7838f3a16a81443da1f2ac87b85a4e4ce1462984391cb02babc93b8fb26e12f1b27ffee9e62a3cec84b6f6ed34a4c6d7cef546554add42a21aca482b95dabb8d94b952e09259431c3e984d0840c08be6c5443403ca3ba22169907e02adb3dbd51cce460e363fdd57aff51d225ecaae7a25d8c9be54cf0e6b5f5a49678feecf5d75d52fe57476fd440d9194a397dcb20087ce8b7e8b324e220ba5b86bb12c81b792c5dd725e28220c05457bce02ce9b196e4013d145c6eb1f18333ae7a5daa83927672ab78d2a3376433b80e2bbe6c62e75f3e0d136387de2c8374c5b2cd53e4054118af90317a30f01b79ccf33f1e82179c71394a641b387a6ca193697dac1fd5c12176cba5060b7b5140bfae1de1f80dc75d5b69f8f929f66ebf92a5e35ae0ac55d45f76810c88757a5f69dc0bce95167a6a6f979cdd1718e702cd060d97fa1d0ca4bf748a02a2d41e2ac5a66405b0b0ff7d6d56ad034eebce7a7b78f0faa8d298f174cdef292395c09b5e1afc96010465611e1b6c718ae4b8dd9d62d48a0c38d0b210e147efe36e5afddc6fb30b61b29c2e5fe4ef4a43ba7de7b0f0637f57086b0793bbbd04e510226615d8e234d4401f746cd487c7b0fbc7f0e67c0d7b171b64239db3609bceea4be5a7df986afaa550e63056f1f102d5040a8acdda08d86a3895a8e93f0716dcd2ef2c486c5691fc8bb907106d94963089e4e05f1f34b7a2d1928f267eea6e16870d6d84010f525f9660f0f089ef851931617070cac7203fea5cbf5116ea32d7dd257374fbca70d6ff6b84c70afb58c6d8f9c267497e1bcab10cbaa98d08d9670c2eb260d2624e42da4e5a8cbb9d038f856b5e4febffe11eaf83222e38d70947fe245485c8818488ae67334ca81a869a9b632910f1e7df712de4962fc54b74ef5b1042019c9a16a1cf64293552dd1b05e5ccae834df86e3dac8da059208d9ae6890eea0d522a4faa3819ab50091e478005cd5b3a238f8d92914948ab2f5555d7962e471d2a013249ce5381c35c1cb2f33512d8a1aab144e78870a9d61424d4c7040de749702d2748062453c761f43d5e7492257e3a1b7477673ef64d32a4127589f7c5af8b338985986dd7d231924cd541db2271464b983c44d7e193e9ff842b5648fef0ed8701f2cf8efa13e496dfb902fa8630d1b4716beef5b345ee90d179e7688da3ae5dbe5add8b606d6dec2962e1faa52a7c75d8294bda50531d665009857a75b6b042d50baaa98e5648f0dac550b52fb0207764417c03625ed28e321932b42c1ba00b2fe3621a701c72db6ca815d0ceee6d0a464fba6b8543f80a9c3c8562a63069143d66c8c43ac9640e22f0ec43b241f70dd72f8b0ae36d24a2cef1776873dd86ea829ba12440e1b08b069bf98d2eb0ebd27fec2832e4fbec014292d362ed246ce14e154786cd509c60e172ad1e7b08eaf51871c738d3b19cd850bb6f4dab839c01b8c0947754582b1f52a842895ab33a5fccb1c4ae7fa84f477ffcf720896ccc93f356e64997b2782897c196e851ed71c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb96eeb1f431357f0f0984ebf752afffe2f0686a96d927140369dbae955793cf19092d562503ece4e07546476fdc84cbe8a73dc3816b2666b0a6337d2e86298ed103b7f274dbfb6461cb7c5a17711bb401eff1465a29ddf984c4914c714e9c6fa18c48effe46fab53d88239c75b80814b658acb31e0c7237e0d94f955e7a3b3573c7c39e0b7aa75f3d5d09de9b160698b7636876834f7355a29d1393674c205394b691396dfbe225e6c46ada779d8d2f163a3ec63e4b2235259a39366d02bf4687c7cc5d8926ae572613c6f8c39da7f79d43b41f1d55473c8020f063aed52bbe6295e637eb488f75878467d89c67235a02fe40f93da2c3c7a29f8036e0b18a3f70ddc84d9e60467043de73b7a4d65e015d7f2fbe60d0a8fbb7dd8038b627dadbb52727f3a016539890f9adf43410044da92e4f35307bbb626c8495b63e6e62e0edecb4a50ac97f533d1de4859d66135711ca65052997f1ab8b0374f5c19eca1fac1540620268ed2b460581ac466391c0a85e41069edabdc91227bbbef2aaa3958e6f72a30bd1c41045b9619c3cc7d6043f6596b1358df7ed2eb167c47064a0ad34a74de1e12ed014e979500acba5e6f183795050b623fbe92b18ab45a4181dcf25f51b1b331d24aa5bed08a7620353b6467ad57b43f2e71f0c63746d96562546f54f823f0555f593b3dec7b2460918ed9cbdb01ae880a334aec6496cf9c5196af4cec985a10f40135f59310ffe5876fe2433b78b1553dcbe05ac070604b4ede8a9f043ca29b5d02fbb1f7dcc8273bc494b6aabb5a4bf114214e1a49bfc5b7ada426ab5b56781ad396c7def5d29b93c54725ab41194ab0bd7a4c32ccc59e32541aaab124d8db871c9b85c8633f0a3a0bea3b6d839d3795c34f01e700e46ebe16975a556256de07936f4f533b0837b416261a75a174ea825211702cf598cfbdde8a291b096363bec141481d4f4d03c5dc5e237513a2c9994dcbe3b0bcb31a193d928235b7c98dda61ddd309cebabe31b45eff62fd24bc5fc585506cebde42855992e96ef8be1b22e6c61549e4b419c3aab533e1c56fd9adbae36d954921911d82e2e1e2c39fb2e92fb7da5e8257198bedba42b147ad5b1c99fe0ef552c5df5904047fb2c466457f4dda4f6159cf1745025b2758901776026db3a6fe9939d91c09f1b2512b9887a23eea22e8c2ad377a678f501f5f0f888c75b868708ca4293b84607fda4a06093e406229b853233dcacb1422a5f4ea95327fad95343e8d04c5925aa4c8995bdca3d29ebd6d5f4d43174442660953f4c624ca461b4a7a713492cfcb9ac1e5df579b647cd877581841d284b47056231ced2b9393d97f8313d0cfdaca47fe98082e778f00f7f96cb4b54119fb5d79fab962faf8cce14eaa439f451de6c6cb178d2376052bbe1b9e2949053d943e722aa0483070937ac6894e57af27f6f1c82dedc70c13e5298e3647ab11e37f38775368bac036493f0db4cf86515b27424792a902628ffb55604bd7056042b785259cb699f530df5512c6aa2636df017aa4bd08e3038efc111ec55c4d74e2de27c7155479689c059b34d361c22a46f3d3c5931e440b2e91a9e319f66a06f9ee3949cb955c5b80f5cd3f5516b1eb44b1bb5cb1ab452a0e335a8a2916936ef5ebd2d64c8519d7ec57c833819f2fb5f223fd6baecff8901de93726ed5beeb0435f857668dc8a5329e9aa77319bc688348e81c13f9782fffd91606158a72906d004e57650162db0c0e3451b4bcb1144207489ed8f332924d34464af0661f40f22582a4b05799e8e7fb4610c928e1fddecf111f43c4478f082150e7e77af4e938fd39c4c7d04091991c51566429f2e1da00aa8b08bdb89b2f9360188e78198b57b20ef9dfac3b2dd22cc8031218e55eddbd1807db73b84a820c197d3bcd243cc3599e3cdb8c0d72b47b44f018f0f88f139ca9aba98a604e9e3ef8e0f2098b344d8a59f9ceb6ac503ed64f0c43ed059c756072935f85653df62a3775d385bf9db472e6432bb770f8e193227feffddf86011d8e90bb73231ccf2ef4cf1f7aaf9655fd8eeee9106a26b3b5507831c974ff56cdb2f12fc22defdbbec8dda9bacd4fbab8d2b0dded6b63095cf01d2e94f64b053be2abe1a40e18459dec292c953a0d19ae175daa6d93e880bb89d5da1af8c7f3b72c1e9d43b4d26774c6ddec42939cdb1764045c74991b8c4136e659bb07e1df3c75e0d0120985b52ee0538c4ef9f39081dcf920e8bf38f1b3951a8f5b73e2c40c677e46f3dfa366b45568b0fd480cc5aad08d653dfaf3883170b95e9ae64358d35b7fa4544004c04bd7182e126043b53b30929142cac6ac6ce1b600dada3c8b04b6daab49082a19b5e37395550facf19f2b114678f36473fb64bbc2b8c7929139d83245f6de42b6ef5fe38eb82a47718728fd5c89bdf5b8eebb944debad0f536817ffd949d954622232a4d737456c87cfac6bcef537e9ddc4255d1a4452e5d34059777d8a2531c92df48dc4d06533dcdf7dbe9629cc9b19a4720c4fc7be9d3441a40faafecf90403fe1f56f8a62033cdd72d4a78509a1492b57fa9853b2bc93709eeb8275768cb893aa708e603e252edc8d9dbc13cb10074a7a0e32b951c07a1632a6e421a64c92d6226c7f26179491c70f386afb8b0a2a904e1fd849cd6459df9a6276ed7bf3826dfcf0f8979e77705f961d57cde10b729f2f9dd70c76634caae7faac2dccf210128932df5a921d7ac8794f9eb7b50250c44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9c68acd1f75d7263604ba2ece261505ea7edd591416db24b95ed96c259fc206cee1b1bbe4f9c6e3286e92e32f9702939bf9da493331caf500ea3ad91bd4a04faac88d4fe1c7f9a7e44e59ee94f1dcc2f2cf100d4e69b14352805c0b5ae29b094854da548a22ad026013c3b6165683a9912266130d3f517f05a325b0672bec12e2923f92100e3f982b1aab856378e30e93a7c7e34e6184b1f3e7bacc68a6ab728fecdbb7224bbe531cfb97d9e1bb5f40bf2125ee11c3bf95301992b9223daa8da31b727c4099b5928b18e83e44f55df0b799fcfa988327e13038a7f327cb302257049bd2ccf763ba19484c605a56ec1321ef081e6065126d13ba485f1b26cd7d760a92603955d9e7197621a56077289b7cc706f787d9c5a0c52cffc11d0c566c37dabb806e26fc80117705a437aab1c549ecec644be878b83ff3000ad2f30bedcbc8c93d5aa7b5daa98ebd43bede3165a45e2464be67c53f9af41bbfdc10833580eb3c2e6fb5b885bd34fbd4b362b91e1a0c0f81f50aec245ee82410613779dbc15739a54290858459cf0c6f00717fbb8cede9353de30305886114daa5db41548705149c8745566f0784e38193c37263386ab91475d9685724c305bf4fd61774793baab0ebbceafec8d6e0f7e5365dcf1c37dab528ed677e4cc7c50779f24421f3569d83fa85b4c30bccae73c188df9cfb2ab2aef127eaee5d68fe8cc937769f4f3c9e0091aa6eef2ffe1f0f8fc8fe03e957ba4bf0a04461edd78c8bcb24cd0cb1eff67b9aff1d857ba5b9f6912c30925996375b4876af5958a02b4d26e742a29bbb79b5c24343caaa4702ca69c2eda7b334c57636304badfdfd5514fabe70c83e996cf9f5490cfae91b9a71d85bd22371a5039d4d725a4f2daa24578095e1e847797581896f7bfc8f56993e2a01dd5abbcd7282873602c650d41889a2786bc2a11d25db12ce5a26f0fa64e3031cb03f40f68ee4b39a3149e61de3bf9964f4e998ed7cb2c844a7d8865169a19b9879a810fa5c50d6cd94d3eaa23fb040bfa598f46fd626fe9844dc4510d397d2318684f4596619013daf810ba61c0382fa055130049c11650d1934dcb61e564a38b170e4cc309e92fb9ae5bc147e065999ef28f66511674b923d42ee53106da2ecdc30e169040024b6ba5188f565aa160a46b9632dee62c22d9c058e5a434e1992109291f92d214800ae4714a79dfab7b9def3ac01d6389f4a2bbb0e7a552d10c45c538858deb3f6370a3df57b0f1e2370880262ca1cd75a5648036493759e251fde361ea155447e40a6a69064e110e709d82c122c441a7529075ef3fb627fdb8d974eec2fdea44eaacc9762460f3f6057a65f48404c5bc3650d46f05d65c7506ca17cd4d4a40ca68d1c72e0ad628fc7faceca78d1e2c5d06af64fd0d6f916d11106587cc6203e9db221987645d0dd02329d746a3d64fffe609d9cb3ba3b3b454a9e52fb4af8efbcc6ef45230582864db54813773b51bd67bb2d9d6b36d9f2e7da894f837d93a5d325ac263f16d2b1ffe25950250eda45ba90441c88c6e33d6b0d37bdbc0bf72999a76e97516a90f81772c46a49f5372842c90416eaf092d19cd9997f991e81d859feae3d3ee01d6c42d82da941a8f1ddd6aebcac0ee993926c871c833e741c0f8c35b7d06b340128ab8669e0b10c021d41f010678a18312fe45f33d17cf2e6099e232f3c45680cb3d8a268247ffd8ee8c530160b36e1a3bc154c61402549694b6767ef62521f4b1e46335a02e15af91296e4d456397c91202a943ba451694a14619bde799bb46eb8257053946a3ce8c28f54deec51cabf52b65a5e970e99b3aaa420b35658c0df937837ad56aef376be4affc69f7b45cdedb8aab592cd77ff6e0765eec1c061080149fb919d57f6142ba436144e293c0b8fc0eef58c33a2989cedea24088cfa5ce4acdfa3f8c72cb689e583ed4920805370d6fff1591f80d1560918b71eb4c2493b36b3311c94b8d40a99d79e17614ea7958ffc080124f22866a9800e5787580467c8f1346c022578c7207b4157612a31ab667e6bcf10f141d0fbb3644722aceebc0631977a44b197009a4d7fd852ea13b81bbfb3705f24c6b3894ee1339e436a78076646ab9a2c36084a4951b7838e22e73241e2699db3f03f2ab48971d2da9eb51d7f8f3b175249dfab146a58e77a6ac9f95c5469ddf15fe10b884b941f57cc4d6735fd965142b34fb530da9e0d0b495b78a6f05fc64f5930662fe378a4f71cd98732330ec4e3437db6d8c2e535eaf64c93e9702e33cb1b8142fd9a20bdd29b4658bde01e03266580818f92c0c75ffba5572bc1b161ed5559c0fa8e309ac69793b59c7586f4f2ccbf53ff5d5fbd0af7f7cf60d22de0c19b7ddac6191dae161fe46c186e61147235a44d1efc0663e4bfba9e2db3aba9bb097243d44105bcb27b2506777d3cb3ec606e93d3c81b57598918853ea55c2cdb6629957202474dfe2999e30fe60157ab7bd1babe236c1a9d61be9fd92e357597fbb7090b1564ba4dc4f87f08f82cb682d043883bb39589b4f13b80086b0bdc96d4faeb67fc2b840275aa38450ebedbc46b36e3cab3d92f04de3fba5ce192c25cae22449264bb59ef1c98dd303898dde35972e222e42af0310f257350ca552f1598a8ad521a156b1fe32a3c88519b125d2f5a04f304d32940c46f4eda418d946e79c75011b3afffb6ff6985337cd699772f3aaf4365a21cc4400648c69f1939806bf59f9944e2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h82deb3fff014c464a6308d5b9853a202550764f97c6ae6dc4dfea209ec20c3d230643b347d9412639a6afb5e936c1a5b2bdedd49b9ae9e0a4982276fc3c1779f8e68bb35628478fbc77efcec2804b965b7ad3da60fa76af34f5a1ddafa449039683c5e0ba164cb63bd85127f73ce52a7e59cf41918df799a7924225fe2c5de19941d23ad016d75c97eac35f3b07dad1509b458078a38fba2217d58de37e31633462567923f72b9a26192b13f5560fc6f2cc35ba76c2eda88c58fbf23e293764c070dfdecfbbe45b25a4a107238f50832f7cf98fbe5e1257f9cf4faa0e511ccd04c4aecc51db8663300f660083ab76b4322d53e396b77b4702b4e735f316c7a7089871bdc52c5da90e9d4ea027ea5cdb5f91c7d09c78efc3e8e878d37e571a64b4867337b018ef79143f1f49f199f717030c4962f65287454d182569bda7bc7b79814820a9a74252f436a83d808830cba6aadceea82fe0b3c7d553df248e015399e7bb5018655e7e131ba27476502b875e64b913e2ef9904b8b1ea65e230445ed96833510389c8e35646ff1eb355b51b57192be2d2de61f86798c296226baa65c5356ac681b9ddb17486197e67bd03c5f3c867499017d3487875540d8e27cdff7a645f00979ea80d63b62467ec07f1e8c25b35856bfe344ed026fa5c6cba1da0e9ca59e6b3dd6d63495ef2e43bbc0c8783817b0f89c41a2ad85c9a77a393e00b58a5e039d3b2ab62e3858cca9bde09954abd5798132d1a692fd07ec15ed25c96b0c6881042fe28b997ba080b0606ade08279c4f43e0b96b855017d57492c932c5ba423a873c92a729f5c281bea94dcc17656ae4c43aa21634932fde0e8c9a5fe97826e2b232cdab8f23d03a110f1fede74e5315593c17512178354ac6076b716bfe4c26c6881b38e9daa14a9ba1b2869c884afd57350ef1cb7cf2949d1a6ee83a40c1b4675ca0352e1f364238d48ca4a787788314fd3a44c0001a113b67a33b0c6fecf9bc5597039db75d097b88c718b90265dcd66c06077b9b5b0a98387ad4312fb1680a683d20a21a137dbe48173743461c085369242ff4644fdead7d33c786bea808aef4f4ba66c274fa8a33fd70952b0ecd9444e6eda7d3e9e150fda10229b8482816ec7b731d4103cbac4551c23955bf88410a41e9b371f32725f767bc2840d4148d30d90d4b96a48b13ed9bb43de4fb7ceefd8684601aeef917c741f3233fa8e69a90dde916eb9f29193accfa4d8e8424897b050ab71736c60d973505cf7bea28e2fbb1f1679e395cdd9b4ecfb43f704c906546d29b08edbe4fc7c810875dd59af2f75d90a3f1f975755c17b6c691673dfd6b3c9fc364635975671a984a296d9cc8690b7978120f357b4b939131df13204579ebc0d5954e295a8f50fcd5c8b94e2b18692a434bc58f962aab51fc13f0b94f25008ff919d4eb7c070b65b00c6fcaa701caeff6ac5672f30dc15c6022a97e4def44e97bf206f9f307655a7a44d4a09f9fdb525fdb1da9ac16f447b409b85a5e0669159ffc363c2643805138481249632b7d2bbbe70518741ee0835f1408b8556b13623f6efd3fb844054b997906456b09d440c5473704d7318cf24bb576297d64003ca2c120aeb20eb9cb22a5c858edf95154cbbdfbd2469f9381db7dc9caf48456d84b70179c7402cbd41f601f1addbe9e7def6b7207a423a74d2bafc278ea2953e96c91cb1228af5da4df1c6a0f9b00a1d08fed84a0d84f318ed9a765dbd0fd649086b4f3fc0482376302582aa18c157e2cae3bcd7cc3a69592ea94977132a0d0ae8335a4661c33bafe6af6d19e807fc1201654725958d21aa5c246d0b920e31878b3fb52c28c3302ec1add4b4d671cb4253efadff1a487496172d1b0bdf40c9caa20e41dda47c4921e88ccfad0f5a827c27dd7d7d886c32f2ac7b2d9609b7df5b46727781986d5868561713ab956d94db8b9bd02744d7962863e20525441c667b8c196c504cdef1f2b55fd2e366c988cb7459efee802348ed4c0066eb672e941f1ab820930d2eff7da5bcb065a12f0b0a6fa3eca50ce4f38d1c3eca17287688b9841a163d150545c99be3fccd2b001d2b30cb592fc60db79659f73ab906fea74cbb5aae6554caf035e85a16f048ce6392a76096dc8296a461e1c3af4676086c17e77cbb5fc638845c7f7f55bb5edae7bdb4db79873d745ca6cadc0f8776383803b4458a7972a0594c099726866563fc314f0440ca55b6b1346e892cbd210df9e00c63a78a66947a00b70728bdd5622a681724f954c5444c26fbcf423f11baf2488f746cce575e628e587504df05ab6dbaac039ebe9bf96463a48e836f708431813273e739c02369c4ebb6c813ab8a87330ad8ead7cae1c387f30c58eb169929299afbcbfee98a5425f4fcfb8b5ba6cb5ef925ea04bbb8f70ef32fa5dedf3d96dc5d36d5f06bae1ffab74bdb625be12778e50fe1783455bdcf86f281e3f0244d1056c7e157ab526cf16bd84abc7fb8cdf837a8426a9b492cd62de70085725a685bb661b296356b2c88cb467bbabc5a5c86c5ce0bd6f0b69225b35771fa5087c0725361f2e627f630a2185a053533493196eef5bf7af0ca7716d4d8661460de50356611788aa367b400fe9e68c33b86ff98f7994c1ea98929b24ed33ac18510aef7c04aca66cbd4aa1ca41430747b6251fdf6c3866b4570dc521fb2a02481ab669629b32e5548d2045e7e812caa1425db709e71dacc988675c0f4cfe2cf8b759360332;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h36f32c54590db89c622bf916aa68e08317dc66f8c63490458c2a02e6de8a2ae964ba7417c4b1c4a79ef525d968e4b952e5717b6c2a93dd309e90da113ae6f257e286ab81ee7f36f0a3d12a3d9b179a39c193afb9834ff6f11eb0e73f87324c531ddc3fc436353242fd249b8af9a6e60b1a43f50f4ebc55ce19a663d0f9fd3df0b7413335b7627dc2ecfa1a7c99833787af59e7692e2e6ec7776f91eee96ac0c6daea458cd773a20dd5f49f321d03f96a049d7a4f0682d38e7dd763c1f938ed34ea6a3b635b7ac8ec32681124bc508d4b5a66b8990af164ea5cd27169485c0e3c67c5010d081531e9db157e38dea301183e5f9c2e4b4607037e6c15fc9ef0ff833113b71973fd2e261dd97fd62c21661047d16be567c3cf6238783fb16044ef0159caa5e0a6550cfb288d8ce539b7eac37915ef9dbe7ba5e1b493ce5e6def219c7581340f9891cdc18410a3ccc94f71cba025e15883b236c3b4474be11d61a8d64a7ca5f9bf8cba96d1362ca28d8811fe26dfa4d5ae982896e6a0d96b75c289bec0deb25e439c8123ffef3f0688c4508d66869ffadcb35629b31466a4f2f93c3a3416ed7e740332eb9e225350d3d4d7bfd363a9323e3b70353c7a87910447f5c4adbef4c156d3161a3bd37df548120d7e8b0995fd02d0b511e4807eeb941f03e1489a937456a96a202ed3efcc8caea74b406a8e700cd6174a205bf5e989aef9d9121af825c585f3cb93e4dc8cba1e7492c1bcd62af352ba05db2527c76f449fdf7f164aadaef4092841c88b9741c927f52913e6f54857eaa608c33f69ade3499678a20cd779db21e14fb5d5dd8190ac375c371f1a4814f34422f96c11c05a10984ab6a30139cea6386ea1993e4bde1c6bc0b4190a24224da9236df7363d6f716710e8472e0002a47aa90c13bc92be73be14738147d3cb660a4ac9d61bb7ce477d27b6ec85b5d855c70a91e5107cc5adc990c5cfc0bfb43ca2dcf68900866b6be76f29ae90cafb19d3468a5c3ad34772adc2463f43d49b2c06062646028d8cf36b527f12a8006b49a90f5d24880e306b372daa2db2c2d5f91dd4cecf08e4eae9423e8f8a451248e174658f812afb41e7a2a908720be202e5e0a68ff0ad317a62708cd89bd3ff12a30ae5f26e2e7ebc1bdf96bb9841b320df1f992eadf006e83582bbca0cbc68b1ba18eb0842140bc71705aadd78013eed3285f8890bb358fd59a32d804f0fa7febd42d5330f345b4013f03e124feb698063d71ecca8e3a2b3f155a44eb66800f26a772a57dd7e5f35a7e3504cc2bca94a45ab203670d43fa4b3fd95106599a71241994fb3b85c6d4659a3d243b45d9c509fde81ecb47b9794a9d3a775d707ed03ff9e02c706b16fdc2f03b7a36b504c8fc491beb5b908518cccd1f34899aba8da700022a40467a272bc8c96445ba08f3a15d4fce18c2249522a605db10f49805d483e6850668bc55cc859557355c5cadc6c4fb84bc37e6fbdb6b53c50361fe86806b8b295ab02ea7d094a5d9be282026311812c4d9d3474536cd281d035ae62b1e3bf197944ba214414920ed89cdbff28062039926f184757c63f004e31dbdc38df0cfc07ffcfd6907fdacc13378502d7ddca8007b004ecaa6bb14a6589cd60d89004033a361181a14c7e38956d7455d3f922e3a8c504747a3551731e824d0e880ea8c8e48cd8fd94a2ab412cc8db7a89e3b9278c5e2037c42ac16e0aac3d7cf03fd92884183627f4dd638a4a92eef7b59e13446c157cc56fb39e31758dc928cba86b9fb318e3169a78855899f11f296cdbdd9e5bcd30aee12335df66f4c5f2f11f45203bf13a8a7f27f5ca1528fb5fce0602130ff65ef0198ac60f0461428ea4f0becc72c717197bfce5bf5afd205906532c4c9864c64e4a45f8941dbc2b9bd85d749e5a09ca90e964d6346e799018dd170c1c0f351ba9b78f4bc15ccaeeffd7bbb30146880ec3b5ed285758a9d7ba8c4ae12b58653ed7470908ab3c7f65e0a4fbef7a66203a1c28cbfccb47d7a695106a44716447082ae919ae647f348cfd79924c5b37136626dc08ac34dc33594b6f54a47e6fa6e64068d7c0c1bfbd28e4e4b7a38acfc9110b6ca0782c1d39c888e22a05bcf30132ab93fdaa7ef351e59837315fc10dd58b5db80e84db112e001ce23732b37509d7ce1191e003fe6d716c4dcdcfd50c7d204684321103d59dab663b72cd9012743ddcd10b2b90411e3deb7fa492974ac8d8ae29cae235d19456b5c21e11be6236aa495f20e2e64128f09face8032781a39a017a5a0e22e26b6d6cef36f2a376c2c6a3577d857e219d7aacf3244de24f6590ebad750f24677390e8ff2a42cf9c42febb4aac0953cb15696dd18b63003041d0e73af93bedd13e120299ceef28cd5b11f7ce45760e37ebaee3b14042e9802a98e3e274714129b0f7d4603d7a24375432f543daa0b6b44f77af01691ea38b44daaafb1e7c33da867e870a15d22e9d4be089ecbeee2678a40c7d793238c211069837c424cd04d984b8a9d33a92154ae10a653a8fdc2176c8d791c417092a814a0a3da465f2e1fd2adf59a5b33cd51f10663ef8e14fab606999da3df2d2d480c7201c038cf5eac8821a67cb9bc0a8fab12c028a9224ffcd62e4e628cf304c0b819f372d70ba9dbcc3044c0fecbae0c1da8b9dee006df09415b41a2c56e926ef5a7a4b2b7f2e53ac773d6c6e148d7268e3a59b350e12bbc97c3acfd5f5e7190af6c18a39e384ec3e9ea6c87a00ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8c7a9713bee1ccb347d0c019f1e23261f83146a89bc677eb35bf64a360137db5a82f693e8a9728fd4be8d15145bb558b9d13b0bb9c1651eaf046797db79e1057ad147ca86b98471e14c1d32bee1c465426de1bb8c08689643fb6338b90f0f0ca2b9d77b6ca9e62f1fb23770c150928cee9d8ab82a3db48bd5b65480d531f87a0d1f3a3cf33b1eb3280259d998ea45a849072b11ed28b2f689179b74359abdf20703fb0be6f0768bf204793bb7897a3c8ea54c8087b1031aade95dd763b1d89c7567d5ca44a6a5dcb4bfcbd4ed0806ad36b6563fdebc2dea1e255db2b563fc6cdc0796d70dfce2e0ee83d27c648a05efff6757d8c37d9f6d3e5811aaa08d31c77a28024f1943b367b2b7b1db546b009de41aae5032a6bc7cb50ebc5493d4149711f309dd4bf8d60ceea4251ff9d66223cfac6bb805a536d34ce27d3692baa7d12c16de7bdc4791c3fc9fe3dbaf39848d743395a0fa9539bc25f2c521dad9d5ea84002905f6622a43440639b86ea5d949d1a09b51090aa9f9c26c4bb73e85d6afa45e65345a0e5931801e695e8f13e22af8840f97746fdff884a15b9b91f9a81323f5229ac78ae6ec9e4adb250bd850f70f1e49a021e52e646b7152443460f35d75bc28d53cb2688813f2262d0898e99a99e4b32c131e4a56238e9af7b8ffcdf726b9d79cb7b3cf60a71dfa85c5006f29088007d2b7310b62170f286a61c5f3c123052b59f79e3ab69c578f4143ac82e767f320d426f2171360faa6c384ac729d450a1f20122134dc3b036dcc550c0601be81ec036bfff570295ba9dd3c880e8c9881f0c8adca83f7ac07fa4460a2d47cfe902fcf0a0b34164f6892cec9d400dfbed2daf786da144491485d67972a0cab650e264c345d803b72a327e0cb5f6206c396819b32437994d61c1bffe645ea4deaf8120be4213594308a2b63f0e3904015160a8701c926d4502ec3ce4f9f1676c737f4e9c92773127a7e3616b1cf496fd6254aaa7f2eefa6532d8427222b1fa7aa2ccf80a1e372d8a53eb6d7be40d1e4c836eed8c0389daee96a7987bff6bf6a3f6ce3fb08efd00e47f156b056d96c9e0b25801ca71e9906d01719fb9cbb57c8836d9832a67d576ccc377d99746551a5d67625b9419b3be46011bf223d5bcd51c1ea7b35026b3ef5785f303c1e7dec5c49009d070e37ff4d7c532e0d47b38af0aed0591c4d36abc8aa41d43af62cb73c7a8fdf0c24dd5c64aa9ce409d11535d8a1f552d71349bfd62b2f8532b6d09942826254f70c9704630da4aadc3394e3376bf79b411101191c9f412fff87711d2e3c143d44f62c64dde90d88f58137bdf1fe919210e727c0f00f5d916c88baa124516473905cebe098074223bdb59f508407131bbc0d5d754c44da2f9c4f0da28d275ca6ceee0e87fad66a48d22f2c0bd2b7818634c29a6893f8a7696359881f519dc3c64288c8e8510602b6105d911aff914d436e00a5b78681e4e68d54cc68f9d430ff0de6e4a5d931396ce009c1a08fbcfa178c2a3afad271531e7b2deb5e2c403a26c1b3bce0c24bb6bddfbf68b30eabc55463aacecb83b564f2696c7aaa12dea6e54b7c5633cdaa5d1dc636c70263c59aa7882c2b79ec03399fb3f2c87f7a97d4066468322f68aec5533e9dfdb75570490536ee5b90b835b0ea60bff7fcbf96c7395efb38261c1b3a385440ee17bec9f00996dbbe6d11cf7c41103560a392755afca588b1560fbcfbf3db1d25503bfbfaf83fb21fa0a525ca2c85fdb5e8e97cc4012dba88c2e3d06e0da310581774fbac27fcd044d5dcff883eb557cee967670a89deaae072c0da8b367a6a1e43e5c1c38e846d5794848f5058081a5bde4068a738791d4f06cc01af784cd29bd5c1c160776d0c8d3f263e76e934eb36f5d52b0b93769648ed7d5983a696ff1dfe4f62687f9ca76b310226fda6c040ec780f905152f238aa1ccd6cdedbfb8aaa801bbf23e8e7ea42f5e90893aaaa3da7516e9177d9ed87fbc89c00557e8002d1add7ffc96abd38c7a9a071b3f1d85dd621f9d4155bfd78ee8eff8a47c0abb0f1371e7cec6ff464f0d167cb00b58c1d168fbde4832ee75aa574cdb87ab5bc6e92db095b89fbd3131be899eb1ef781d256fa938078ea1f476a1cc3ba8ee3f0055f677ac40f55e3973fbfbce19d4303e0a1ef53e9b84c9ef60287cfa37b12c0eb2f7431f01163f5e3f1bf34d4b7738f5e0ae723a39e34d7b32b65b9fb29556bcb046b37acff331e8303aad8d4f919946a4d23687d2039b3fa4755b5e5fc9085e7a375a074329ef04d394e02a643db0af8be6ef213188f01476164f27d9dfa9ee16531e0b67303cf41b6c68a791b35379c97d62538d3bc0cb9ffccee891fc2ef369219b865c9823009f11912b9653c4b61573f2b06b3470bc1d5f8217756ced69c0d296be6dafed343a214c767924429e50f9f6ae6ff3063f3dc45b346ae2c57bd752540d70342b769c81813ffc0b6a037e8006275f9132037615cd50ef51f3b170a74649dd801e1e14d2fbd4d582ca607e0e6b3fcb79c3be272c224c2f0c9b61da988049d0d1c52ab074b400b02aff6b44703c58ec6275fd3503725f9a5c4b52ac240db640d4d89c505bfe06a6e77da6c4df352f6e12e5533d8b7c324addd54271dec327ec4ed2247118450010dbde86b1d4a5d2a1f217190921951f43a9977365f7f169d7a7faaeb72ca4480a0395f2e486e317709978f84c7659ab9507e26811fe225b06f18269407391f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h925c4bf9a5f139b1e0d6c2bad4ea237ed9ee35363abb6c8ae82ef5150942b9f3d5d56a5db96596309e6d1a7b32188360c4b4f6b60deed78c7dc8bcaf87f9155e4738cf95baf3cdcce4ef80077a7c91cdb8b069586248c5186f76d02b54b6f80f319077fadd83952cd2732b8a524f943a6b03080aff0bc003a2e50e61f603d494230286637e287f0043d02c23fe8f93a91b7c699194bf383c2899a7a1168100cf70859246f430a0b7c1a1761d164057f8f35876ba4e4d979f6cbf5cd1ebc1ba2098fe971b91a73567dc2c41805af642e61c962a687eed2a94c3827cdab415a74afd54c53eeb38101a49e6d0341af03a5a791563dfac759328645cd473587720a6a88f7933c9e4e4b175cd5b8393a31d1dece3f799c4215f416bbf946d629b67480b53f12461493fcb4db999e50b2b0a1fb89cdf282a917f690cf5ea9141b9819ba5d4c4087053c92c8a7c2aca13159101389f7031538f47f85b1ac663481213c129b393d157159ff87185c1ad43fe341897e7e3c92ced562a1b0a591f3ddcae95e63c14fec90fdd6800108ef82c91a6251ca7b85d00e1024d919761f7e217aa21055228615def214bf6c2abb76d5d75c5073b4069a0be07ca3873b8c0883b7e12feb5361e372a7efb3bdd9acd7a8d4221522db47af14e41c356129664820b65761f247474b73b1a2dc23393109486a94f8e98bd3c92d55a57fef65702e0277931916b022a5ab730ba40beb4d73335161845fb88adc190c859931a9dcd789314ed5eeeb0570fac0f4ec968b9d0eea935e6da0dbc6cf2bdfef91a2511ad63c5869293cddad4c3d2421876c2becc8e9c41d0b356f97cdf4ea043d13772a7d8ce383096eb52c881a8839e5a43539f6e54953e22250886369f06f2ce859d9e4d7e6ca2ed6e3fecd6416a4415faddb7ec5fc0166b72fc4b843996e2811923360408eb11423f859cde65e2c60072572312de0ed7694978daf1b4aa48d60472c32a8561eda045e9ef6338778d6716e362eef27e61f856f4cc4e850578f0ffb12eff46c8977af15c9a03377b60a83c5724e4a118a863846fe65dd2359429c8795cd6dc80460a71091500d935164459a01ef914715dfd057107ed1fdea9ab3944964876aad662fa0468609d6560c5d183ea2a874a7ecf4ff2ec0656a9a02e649067a5a835b12bca3f6d77eb07a8c2488bdcfaee841c6f211d1f7a2e14fc58be9358f4cebe98f01ab00158c46b67ec50a8bf38e7014e852502483fa5e51f7fab4bade7ac3380bd6a2a30e98e37824588c8594784b477a8e4b7de00c60a3893246bac60feb2637097c806add4a0271ce00085ee0a6297a40bc4690d58721d2361215d8c33012bacc194c4d0c6472fab632fadfab9ea94596a9353ffd3025b507bf7bc23ec31c8494d404fce32e097d43ab14df2be420e54a499ae00e4c15a19681a1d15580e869b247a4622a798d8dadc159f1573fc9e76bdc7f6825626e068e470bb4b5ed60bf077202a5e0cae00586c31b367dd40c1e39931624cb97164da5b536162b195cc7181c87509be6e5d33deee1d8ae53dfe4ca13cf62bb3dd807e57d30c0b1251993f3ffebab3f44728756b6381e7cb17b3ed3759b994120c36e8db526affa98644ab35314184e86e148dfd4bd3ecaabc6156db363f6bacc6088fefdacd1c4a4a9d295017a3f0d5d82bdbf7ec3202a8c539a4d8c0cfce0445c632ca59a076d4fdeea816d783fb08d5f2d27f38b83c424b7ac979390f1e79411cc9ba62248b981c6c2300c7594f9c8db7912f42752943901ab89f763935cf1c6c787a399002816b4eb6f57e4bf866195ac78de7b101b1d13472d15ffd575cbab99b9d2838daf8321008d4909cecea6e7c41a283c927479609095aa73762faa6cfefff6615f0ab39f86854aa3dae7b7fdecbdce7cc2ab2e59a85933029f47ac7805398b9617af21ea7418c6ca954996de38d910ec903ae1a0640aaaf71873968d3f2b7a787a8336a48eac6d644e3010e0585bcfb7bee5958a635e77d5e6fd4f3930c0f002028ef7678033895ddf86a2fc63e2c2f20af1a868dc3517327feca7a688095804a6916de2a72f93739a2a91c16d6ce671f0fc9796d40d095fd50f058a8c19e7430f4d54f227125de633c9cfb331e825847ccb2c49f5530f50a565aed1ecc55a862a90aefdfbd59b814ad64b7e0c3ea236fabeeb9fb34a36a15c299d3a2d11e588dd56763f20009e7914849ec8c607540a230d96055f8e2acff85948168e710c49d74bbd9cf92cea94edc9bea168dc117b7cb28f93a695e3374580049326609d827e3df9b656c21f93e59f93b4d70b9656b8ad12d9cd8517d85625a049815e385807a6d5eaf01ffb137a4d0c7bdbea196fbf9a6b0c8900c01651a45224ada2725abf9b03ef0a342727cd40df50630cc423d82e89db677ea1d0a055283780d961637aab54cd8e5cafc6274f2f9f40fc926333383bb8c715716b4aaaec083e53fdef0bdce76ba5d3ed38d442c61bb3cd6025d78b8d5b87acbcfd5f44514b0b46a59551788fd84b2d58482aafde52207f631d056469b87dc684399b6c8dc5d6abe7a28fc745e14c64fbe3e1f855a22b7ebffdaf837300d979f06875d90e0c15ed227b7f6e14a0b543aa7aad28aff4da5eb6dde51483bafbd72ebc74aca05ae749f534b8052fa24f8baf2782839d857524f6f94032280e577c8a20e5b400a1c48cff76f7905b437580c6484ce4c714c74c566f1f4f2b6e244f45935b0ed27ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h509883820e0bc70b91c1e6508089c986b4facd66e50ebdd3b6f027a117550f7942d48215d505111130b34d7c1e9564e120a4e01f36b6e8c1c5f3c314bd8628cb310c3380b0ec385c863e681dc672a86df8f0ff3f1de69160b5ed7621fab1b35a8b2efbea1c1d2cc164fb54386c5e7ea74b73db83cf1d2d8e4484c0e2a15b97df03e1686999245ba27669ef07b295c1f68dab5e5a7c72b0f4cd8555b5ccf693266fb724c9e5e9882bdd6398bb3f2b395f899e69e411bfa043d685b9c7525a85c3712d9aa54e990daa7049a6b0d77555148edc5bbc5a292563ed10349465a5a9072162baa71824317d8dc19f15efa3532a9b733598784f83f803ae9d441a294a708b413ae0124e792b3e020e9af369eb8b410d6a25d6b905327db4a52cc5e744f3aa762702e6bfb35113053d00ea57966c1ce0bf5f9f58d2e9e2dd9798696edf4dc92cd51347475aad6c5802d45deb452469cbda5af881f7040307d9cae2647800503353b407759f872b38d439d540249c74f3662d54df163680c3ed9fe65e80844945613bae4ca01a1aff7932c4fe06c44ed78665451c3098c3b362595fb47fa7a3f86a1d0288e9d0e01a7ba278d2195d97b96ee7f4abbdd00fcbe74b20b14d9a25225de52cd2c9faf72da574bd4bb7b9d5e12f84f6fa635a7d33471b74c0719dd2552ab8eea3a7204abccdf7fe3b363f174f7df83dbd2774ee86b67eb40f3f80af01c0bc80a257903cbc86d7ccf7f537e154f906625b7e1cfc8082f3d021268d57d86a2e177f3f0d238a91c51b03d1896e4566539d42536ec9bd9576538f8b36ec075277325325478a7d3260a5fcfb42fbf844ac000ab261ad4f1fea30215fd34706d0f51aa11049da1320ce84711afe8d8d4bbd0b1c46928468934fb6b9775fe57a36bc9d680a3202a26ac0df791d2cac8321a5678fc088234fd0ba2022fec8be0be5dccff901717b8d0f838be2bab6a1f9e21a768753b5173b1080f9eb84e5d17115b363f754d989c46fdf3e1a018c9cda49a5df58ef76dd445368e665796b7177872c2e7f719c363953cd8dda2f27a49cbc030ebcbaccd58a3fa312cb9f106b6bef514583f69781fd863937656e4df31123a54a9e1cf8539682ee8f1b383d6f0d6c642534d1233145e9d4ce7c62c429e71b89dad33e532a648d888847e6ffa3aba015546c9e0b878dc258b53367732b424122a78fa890a999a1b6bab21ea65a54b135998c22332364baa119352bf95be17d339dfc7692b91b6052d53d51f77203f26340894abd701e55625f7eaa8d2761170a6db8294283498a193a28e72cc12d40701ee3cf37c45219003bce9fc921452c7700e8989db00196f67700022bfe8df5071d1fbb9379aceb49203205bfbcbac2fa8adea862f212eae05724a044ee3e5d7c5fd0b67169b1f524c4eb32c9308d2846f6940c874c4c3e2a9a804c3d448f78d56e0417fabe39c1ce7b950d741e73e518d59d81a5e370c8bfe62fd5ffbf0e37309bdf33021638947a87d883ade73fcfffd8ac38128d70b72e2a2b30252ad131b420dbf3d1f097521ab493d6101c2e38d8df15db3227824ca0bac0d9b1b2783607e83a9080915847c98070576758d726986852ebbcdea8e9ad433560635096d7f0fcb3d4e6b9d02e2b4f5ce5451643b74b95b7d8b86cdf79c98447d628b7bab161bb4671a6f7ca879c6ee19c61c28423f60642347659ebee10b51d038b2890c7e0dbe873e7495e0b1d32d28c2f4f72338b81a7edf743d86d9afcd6db94a31c2918de8ca0021ce07a54cdd1fbb0b18739c23992d0ceb348df1c4cc27f123bb9fde2735a8f8bc386c9dc9e71436e86c8bb128b35c697007c7e2e683801ab22f86104fb28b9fdedeb3eaa2c103e54b8a96e1e8d369f1310fae5caccb45ae0e7a96e079b3e5b277786fd47790e33a9c0b02ae66d5f2440b43957bc156f8d6dd9e870ef9643976dedc5f37da62bcd694ed3ae0d61454bd4fdd76fecf7379c8a650b0f237c0952558d2d66a6bf7ab230ad7195acfcb2cd009f4600c0a3ab0c7b175fc2f81dcf80d230cc554fc5a254b3b7e1f8fa2aa5da7b5ebdebcc7a6a8137f122fac025004c5511141237f8a207ed19964f1ca63e92ddbf1c8fd376593ef7595a2965d9bda3f835a6ebe561af3599388e76d5bb5970832743d41e73df70e48e0fc42e6b6819940a6f3f6d9abd7a7615e00ad6f48aabedba712267c8f110056d531d9562617bb1dd2c856640cbc52fb7dcf3a9bcfe44c5608c6f9102c4ee746fd3d621ea361766e055bd4f1c70d036b088ee675f8ee4d2f059efb92dd51920f36209370a8014de8546add451605b52279c10854e8bb248f4368df030fc48ffd079834afbbc73c8fece8fc6d59654b365b050f111a4a3bf33c701c0c304055010cabc5c21149d7235253592fd90cd9e0006b70674c7fee9584da81aba2013d704b6844c027c45c4e6ead999060f8799418ce31801f9e91ad5d0be3429e96ae5d41475b80bb7d961b232ada43ba8c2707e2d91f909120d7f3a9a0bc30cdbf92ee8650647a0535a183b1f31d7ef7c2e3c530133b1b7687c2aee01a0b7042a37a8af314f8dfbeda88e2ed56cadd33a90f62815a09d799436276655302012b2e767c1287eeef79c45b3c02fb32bd06f172a586cd5c5e5896f3a2cbf318542539ce343e61321d4d88660e234aa8ef66515028a6cc102107e72941e2bd8b029c62583e9e9bbda272922161e5c1bd6e8dfe4c8eaf039411d7c4880;
        #1
        $finish();
    end
endmodule
