module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [16:0] src18;
    reg [15:0] src19;
    reg [14:0] src20;
    reg [13:0] src21;
    reg [12:0] src22;
    reg [11:0] src23;
    reg [10:0] src24;
    reg [9:0] src25;
    reg [8:0] src26;
    reg [7:0] src27;
    reg [6:0] src28;
    reg [5:0] src29;
    reg [4:0] src30;
    reg [3:0] src31;
    reg [2:0] src32;
    reg [1:0] src33;
    reg [0:0] src34;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3])<<31) + ((src32[0] + src32[1] + src32[2])<<32) + ((src33[0] + src33[1])<<33) + ((src34[0])<<34);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4700e1a880f0c2a929e544a36e3813c035da4ea49858e98983b425b55619555fdb4de4a2ab914d0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb980d24553ef483d83b94beeeae0672096568bb6cd227e376e70ffdf6fdb91bdcf7a25fcc74c30949;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha27b1261556307a7f5dec2bf64c3a26206d121735bcc44ec7049b521bb179da5a921d5c5badcdbbe2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2b7a2230de237820aa4e17f8cb4d18e16d45e38ea56b3b5c9bbdb2dc5d4dfbd659e063948f571930;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f536b373658b1da47a96a768b29f841735a23659287938692eefd8e44245285112496980b8d48f1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9581ecef0b89da6b972475a8fbdbeb7d166a2dc5a5a321627d26f15ca86b125a85b8119e2010e68b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77a27f95897e09ef7618301cd3cfef1cc31ec42d0576540cb34dc4e574bce86cd066e92e67c0af138;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cb1c4b83914eb10c8bd9faa3af9753ddeea6868a5815b50edc00037fca533c8732605ec12a094413;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h595c71cfe9862235e5da22ebc202b5e350112bd167faba0d53ed9e0de0bd281354a6a5a205c614093;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1a7ebfded680cacaeec8186f413d37863818442cf66d73b519646bdba4221b20a221f291da1b168e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e9894be5779c743b746fa58853789dfee81036844325f9ea49e5aa8f53272e5598e5de3df17cdcd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a7d6309e73bfe4ea3b75949648badf2477d9e08a6fdbaaf4f4b38a60d91eed5982fe93cfbc11a41a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha77d96ee92396925f9d67486a66c1bd4b7b5989d5882e906a43eda64b807be7cc58158791849bbe42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e12c0d9d7c3a1f32e7cd662ae86c649b9311957085ef1d191f06f459c32ef186f4504cd15672522;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c7b4faf21a60e89e4947b117ed5119d102ef55e69a45e0008215f69f61877bc335df7c0d5a50ca2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c5040fa45efad9f99a3528787c2acab2c725c5afe6a5b203cd3e6f9f2fefc3bc9729b98106c1c6cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12cae6dbbc4777506e01582e9d800aed3ad9de5b4f6ac661a982a17c76925a79731df58ffbd7a1e63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6817d57d6dc3a773e28cac37cfacbe735b689ed5678c098754f3bb0b143e210d36f1e38c92eec9454;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fc855bb4f9a0cdb441879acd6f954593aac84119e4764ecd8ef2a1f31b03686dd88798d208bf6270;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h427433efec78ce0a1506fc15428e3bc88c6922092a56a8e5a94316267df837ce903ac7f0f0c134ccd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d124a2a29a075866adf9c049771d5f4b13643c231bf82ddf97705ff306367cdfbc9dfb81671e8e9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h195a4dd0cdd0ecfdf0f71545edfba6292c6dd28609b3fc4ed2aba0400d1d622b49ab9db7c7a234b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54be35872ff4a6dacb3083b4badf4a8583c218f2c8ff43063e3329d4f94bfa288a9a16dabad4f04cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3f6855001f123ebc3cf334f75a2e5608223ad5e2dac1ac16cfe31e04c51c3e228110f64bc351d6e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0004c3a2b8f052f6820a9d9a50e020cff01400cfe0cf79034f974ae8bc715c41578efc79340d5b22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dd59fd90682e12d03e31209b04f1968f7902f0467d54775c944e792208b9862333c7477e874be8fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf76de075b1be235768dc7c090ec858df4e283694444dd8df61fa2538e306b4ec8167593d28f069493;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59be60a1fc018e0b8589229525da37387d5b563825a4ab350839af0c10b72d159bc022c0994a9503c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bf68d6506ecd2c5d8485b546d31b4ea250b77cffc8d84e1f2e02563063107322c71bd4de7e40278c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48310535d39cc271bdf2b965d8e87544308aa78f1d454f8461a1f12106ab59284f3ec58bb16f8913f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf517239f33a023294820197741c17328e61d3806f73a134d83959e334c92490262ecf3f039984bde8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7dda8d16d7f1f87cba36854f179f81af947a0ead242ff5699be061d7725a40a98f2cdf34e9e40047;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e30f76e4438a165168df062e3cf9ea9b3f7ba4e9b71278cd1ba056ebd68a804e20fa61c7018caf9f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e40a49a7b078282b6e4fb03fe7a824bac03b657d39296fb3d72a03b4642fd74b1772e639a2bc9bf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b5c31c5d660267ec7db3fe013200c91b203aba3a36f99014ef629f6d12141e39dfd45e7e771f5393;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfb34af51418d8f2dfbab7dd669883928c7fe8f897041755ea882efd4f0b01963d47108a0faa6abef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3872c3710884d5d62592771b12406b02e19603a0ba93d3495e1461b3e7ea7f4e03f8a99bfe203824a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23e28101d29f0a4d4f5339aff7ef58fd194bd6571a9ff48bd42d8b4cd76b019c1d59ec79e4b42eb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba8eed78f647a25319233c93b5c678549a80ef44cdd3d079272e69c593bcf92dffb5b411e9221630d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fe4ec8ac5581a8ab68848b0e075dd86db4aa15eb9fb8179cbec26408a6968ba42def6da8d866080f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3b5959441603c56eb1c55bff839e8d764d9542da48a8c211fc1719fcb5079904dd29b06994785c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h330cb49535831a77f15c46534d683a0cfa97c1903728d0c61c269b3f4bfa758ed0ba98ae7d5bd8445;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1f8fda6959189a0b37665b6d5f659737e0a96ce3fe93d3d6c6fe1e188c30c85d70209d3bc2f46dd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h241d9f61e168a212b90307334f20a28bfc207e6d84ab8c9b6563a1a8064055532171c329205bec461;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b08817602495bd5b490edad7976f281b5e504409257a10dd5ab2b1e6a651873ee7f1a16a55bec8f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dbef161f577bc342624658cb3d7111337bd7cf450770356fa857eadd151d41a0232aa5095a48bf9e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5259085ac8f3d35dbf373c0876ee2a67513db157356f352ecd9f1cae33eeb41cd98e45f713bbfd6fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ff4ccdead0fbbcfa1775fb932a65e9a0eaad953e36686292a6731a66233da0eab9f49ef637c122c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8fd83c78ad9bde33b8f60d09133ea3fccaa29a791568b0cba7c93f2b45552e79e5a8628edd3b4d37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66a38a3b731b635622a864bf0000b90981f747b868481628c0e1e294f932941f69b35dc1b7142076f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49a35618e735d3a3dcc5a0f4fe46a061ea8f047e1d2f88d45578fb7bed2d6c2edb5e0829c76268910;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h273053b7e72298df4f165372a0146db6b0ad23c99d35e659d47eb5f2aa9ff9ed7faafc6d7b6faf35b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd08d9d2165a340eb5b84a5094c40b2b1b78ddeaac2d955c84265290e5cfef61e70bd978dad3ffe15c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a79a5566090f8cd385aade6b368016cda1ba18978b31babc3bf656d2fb8b36d959d104d5fe4b32fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfec25d6af885a10b72d7a325f94e729038111f43fbf381c1219402b30fcf95c925030fdba1ac957ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52c00090406ddce735c90d639ca18d83d947bf129c7a171d1073e0e9a76b43e049593b2f469f8fd43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h402f609496e5eea571762f7503a7ec1a82e4503611c81cb778004cdbae49db4feee31547df698c4d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdae8fc0356b2746b6812ee7afae6c925e0eebaee55e073e77884d4c586a731be160084ae7adcea386;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2afc68676063467a554e5b9338fe97d3e74e22078d5db5ff0474775e1816462e7beaf0ae93efb7fea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15cab1267db685ec1d44573fe03fa15521537f918b06e4eb4d176c92e54fb653062be81117e9de150;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d7076ce0ed96822f7dc841c731163b7021be01663d74d75bdcc0f634be37998896aa4cb7de798f64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9abc3cad540847ba26cd560c2aea89263e2b5fccd7da9fbe9bda3fa1e4697595718b0094855ee627a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha155578166177e7ed6962116e145ff18e6ae2b968d634e4c45a5fc15a34e72b5a33bd2a90bbe2da96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d8ce4e90e7e20ff8132ee8f6d4bc968967741569564fadd0bcdb6860f4d435cc457a3b1d221ff768;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c83c090ecd5eb44db86f4ec6ecb42d2f50d6e43debb72f06b1cb517f281c5ccfe9b42ab848ba221a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb17aa181b336954b9d90c7ed93a08474fb470ea7357587d8059bf926ae3b8523c7d4c5d8883496ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80e3ecfefc9a7ffd6dec06a455c1e104cfe685cb713b89ccf3302e9744d703d66c6cbfeeb00d123a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaa8b6088ab07037d4e866c6dad9ad8f71e41b27a78730475ad73a8ea3dfce14351fdf6293cac94e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5472024f2b30c56a0035081c792319322b525b7c464f522df6068fc4829ef2726b58b068b3f82bbe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf077b7b765952a2a28419461c2ad148a0089cf0812217b38ead5c982c1be0fabe9aa3dbd2f1b7ba55;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h568d04cacaea292ec3eb472767becbfd4553f87a021237e02032e9048d5bab8748f7eeca7d448a721;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb74c14485580da2f5f037ae73537a274d9f2b50bdb6cf3aabdf0e9aab37ce350968cebe94cf7234f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd18733ac080aef2952e579068432b3d3a7a0385824288333c45a2b4f80ddefa7f3c051ba3ef72188a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3702f5233ca097ff3c7a6e0b50acf624e7c985be480f0f66fb0e74e3e34d3ba88485e4ccfe7aa10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he533936ab8d4a3593158004c98cd63127bfc19da3e567345c71ba965d9ec6a6059c5da020159a5f90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76bebf781f174ffe01fb5225fb243935b1f57e71ef7cdcc4c3326a1becb2eb2c487fe948ce510cd06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h893fda4d6f6d992e7c3f8b8eb4b63aa1a60728a6ff566740d79079f7814c0708c5ab9627e58f4c006;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a75d485fa9a389954be0f9ac4d9ec1568cabb8f37143910822700dc6039a34bcf015a269f84e0338;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1625d203d880294a486bf3b1dc743effe1d13dc8267a40d2ecbdc2c9ef09ebd86759149d465acf732;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1fbe1fca8f9a9974ff645fc51263cbeb78bdcc6b5f85e61d5efc364f16625d89201040b2254d93d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfebbfbad611085243184d78c487511838293dddbae68b162d177ec99b843cd7dfda3f85db33788977;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd284cbce3bf9a1732ca5aa0328b0fd29035136f529df4b0c0d52771d3b1dbb8be001c9117f74b82da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h814e0be2b04445557215b4d9a76ae50d46e47bfda8c7991e70a73a0836d4b99c9b2a39228f3a60eb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f1a3350766c6a5b00b0030f00e98f73620a8f04ae7025062f177d4f1ab3e1df2d72ee15f75c33e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c65dc7b09a13adc81e22b693299315c293283f7402e5b92dfeb9f57b50a195644e0b772f234d03c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h681e0ec1daf12f3db3e0fa192fef5f8b6554e75e7d8efa047c873bda3d0eb116ae2204ecf677566c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f7876f56831efa06af621f75b6f7ec276343b913785e04e492944ddab17627cd37ff3a661c91d620;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c6e85c7434dfe9daa39f0b12dc05f4c575adc8aa59d6b95e485e39b04553de0406f8a7e0ab1da03e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had5066b375928801e57b64764dc9c5dde750e895acea58dedd6867657420c11bf3c98b9d1768bda8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3e25c5c67a640da7ca08c1162e05afb9d3cc124891c68f5a9dd37a6bf83ac3fffc0e2b3306087f44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hededba4dfae3b97ec1be68c3dec055a6b9ae92e0f84a4205a11d4887eb7744945e6033df04426eaf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfd37596c607eca18f035d1694394bca16ccf90d635b177e52f77df4beb3622ba0d2958b9c8dada44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8642a3efb7b0d2cacac8e57351b4ca1431dcc47e43990b8f20573b655f173466ffa85cfde07d81c7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h712b18b4fcd65d0c9d6a7523f3b4475691a2ffb049f2e553b7dd73b1ca68b868de61f620b8745cb10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae5d8125de12de9d4f8e558f3cfdc1b439c53888c768406f20757c263b4cb84e9b582078324a8e494;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he31e24d849c99df7393bf48cc156ae4b1cf2034130a99c604de6ce9fb3acbc402f4a26b5a031598be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cedb2445dcdc621250c73c206878301cb32f4c3726e27d369acf27bf88ed5e6ad78d870ac4ac4ab5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h221168519ccf5b73e02b6f21375bc1ead328e12c8b35cdd78ece69ebd717e07e5449600a6f4543e14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ab181e8d1ff78442f7b65b66784cc211019b0b43d13f5e8079f4c692ff62b861cbe6a43761e32d86;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2698eb4c3591c788e10dc854a716262fcdb69f3d93401c6d50abb4e5e6b82878fa39adeead28f342d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9d2241c55cbcaa69e151c338f750fed31ee611e6033b69a9341ef446ac3366c766b57136243539c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66eb9a53357bd5a43bbc7f49de935fb514e153f7432c0d09583cfe8f7fed5c534b9e71ba48f6eebaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b888e0ab31c14096dc0a4e5c5029d6db0cc7774daff79de28a2cf898b02c982939680e1ffe9556da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6643423c0b52728882ab5c6c433cc7605da35a32d16cc1a331f99eb6e518f3980041bb4288f6a769;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdf54e179495537d2ac199da14ae94ce8a3f6269be4ad7de363ffc99ac5a9e43e9f754d93e8be51cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ec8af59f488ec525e3204fe183322acd203cda3cb549b9d16ff7df2284c5bd00e37cbf5bb754ad72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d3c6cc0037f80d536d5bb64a520ff0494dae6bae0935c9f520bf5f29a4af019eb8205b73c4b4e7ed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa4d2af0424cacfc5e237a022839f023dd805c62a3929fa6aec5f3f09578096f51d00582bbc9dd2bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d990b051b0af924a47a3f5f22cb0ddcbc9018fe758e86cf3a91e93e6bce83e84358f3d275af0b07d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62f182228ac5ed7de6afeb3b319574e91fdd29ffa9761439bebe9d2ad61c49a43faf1daacc24b20ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac2caae96d81fe9503e278a90f214e6a2b98324a309e1fffb644a7bdf0bc1bf501fb4b0921e5915f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53b1b75a9199e8011e6da84444f16744874bcc8d3e2d4c3a2e11d39d3fdf0384fc40450d9c5fbddca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec7e352a4575adb27d42c2f1932f5f6410ca9e01e4d10bc2276c2d79e53fd6cd7d330dd44fd33be2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28145c6c057cb4710ee33114e1add923ac2e9404523a492f54332e968115044ad1723e17f3b8563cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a5d690765ac3718f7afaa46db500f28e4c4807c76ccb6de5860a0442c709e91f096e0e12f50b2084;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeeafca13d8642d89ff1d30e84092f4e887ed6001aaee0af8d2f63c1c710cbccae2c2a5afbb3c538d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84ecbc00afcdba382ccac459e588849efa4935ae30f966792519cb8280329cba918b1db3b94265a24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81faaa818b43313e544af2da44e0ab3e5c51ee61c9795f0b9ffd5fdd5980fc8c637fa05fd90f3bda5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20b02b46532316a1dbad132b5225c4e27ae114a46427b8843cf54827e5478cbb11ea14c8622c7e7fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h812b194fb36515f2cb3f200d8eaf85dc5178952525c1e77142d84eef5fbd8c127160c6a24bec8e84a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90d5299b9880e59989ea16a3d75a2fecd0dfd8f2683dfa415d7bee78f3c424c1786fc9be05d288319;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd57f352551a79f089e0ac9fa26ca44c7cbb00b29d7d14bee03bf0bfcd115e8a0369d8cae180396c4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cdb86c73705b66762d1fbc45d79234aa129984ff63a302d430d433f05abde2f2cdc5f1f352421351;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1da816775ab97f4bbd863fb2ea6d065373fa23b3fd8dec5ff90dd77076bac4aae51b031521cde57a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91cfdb42d5ed3f731b4d779ab3651663a64f35d715cc33e17c763ef7b8b3cddf58e99d3db5475f7da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h639aa569a3edadb07cd1835dfaf798dd61dcc8523934960db70611d2699dd04f797648b07edaccca5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9b30be06735a7845ec14b24992c5530007624a3a7111b78608d3f77a298f3417e42e99a1b8c7a16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3bc69ab3a177347e5d1f30251c4df04b0f8d1c82618de19308ed11586d748f516329f28629d46c78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h277a677528b0221ef29fd84f4c8af59cb27a4a0a40f893a3343154fd0a4ef172d7f833204e3e67bc8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb65706d2c8a80e2f91c01e7dd4feeffb883e729f91f48237b4605053d7521e169eef7e8b69d92b40a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25a456bfed83c4c87cf102b080c2c1973081942635938dbc05b77a9d0f9b4e9ab797b8e2da1007391;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h193f13b1a587bcca29c74f44e9ca64c6fda7466c7bea69b1ffd4f7c675535b18ddf2ae8e24177987a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a7ced9edc2c7900c43b11d7cf98e96f300932617bc601f8adb5d6f9f843deee0b342f2adabb3f394;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h439a0c985b513439056c78905a67963da84ec2c9f496bae23ed35cdad89a79195559a2b5e84fe6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cb86b4a621ccf94de95a5e50c5f6665543d71a718d70a287442017d2921f6fc40a336c128e6f7e64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9dcb3b640073b6164b13cc78726ea13bbe5dd363e40a22efeabdeb0b41f81175358dc11adaf8b69d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44af0c88e8d078a875a30a166c79cb986e1f409904bdd10f616615b20f78066cfa759e56abd4a5546;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffdca1874b136961951faf0648e381b5725a612af968ea35a841e9ddcb03388cf40947a9fbea1c3dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h751f23e18cc80925f540306b13aaee8f7e4bbdc64d743f0197932e291bd8a0af48d9e6cd6f0fe8c44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8681c2b9e923b883906d75fa301e5603411e9bfa7111a11fd00864c6b32800f7f8e8b028065bdd9c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd675c4ce7c6f7c75fe3bcfea292471f9aef06e653741fe1a6e29092f7701e4417180373a8e7bc2a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b05fc243b46ad111a060a50d6cc5ffbcedac143abb92d5b7a13af9a10644847aecd9660d1dc3d3a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb8106ce970bdc373cc407f79fb4d14f26f57930c3edc1a6fcfc6eb1620ec19af7ccb93896210bcd1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc619e33883b4ed014ef9e7978d11e56e3bae40447e1871e744b21338332fc02386f4eb3f23e2158e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26b3e3c55f40e1ce573b4eec9cee1150389c6c2843b8213eb9747d012845d6b0fb970ca960ebb13e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3a8dae3730ef5068ddf221d2dce2af0d82e7f2e6b7c21cbc2552a1258e7e9540ca0d64461202a955;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf950e2e685c5025ae2a11cbf8ba1e7190b18e641aaea5146af381586aa2f17301f7e634f207aff3f7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4ae777f1491f0a3b2ba39868e36842dec3fa28563e36561a8c36fa7a6832fbbe809ad13e7a6cccb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a7eeeb0227ee646a688535b8e73eafe764c9a627f5024a2ff37ef14c5ebac96c61da67d1be6fd829;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbeff4fefb020a505c4395876778064d3df6fd1dc0c8cc67d7a51ff88593fe1a09055425784f92269;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45e1d114eb59db91406863b401f71b627911a55b90259645b78672f5fdf6f763003e4dcf0c2bc23b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc191f26028a0c0321035574e7809863bcb2ba86404b2f1701bb2bcd455144877378100a935c8afed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4022aacc65586e19c4b4f3774bcd9a4384815dc2e7c3b97c57497af9231a7d3535fbfd56e94c9aa08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c9a835f5bc77ce7efa0a4c7980ca4362a4b347f6f9613bf5fd3242a715352ae8323e7f1cd4af003a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd220aa96f02e82290d7df37e212fae77114bfa58d9e72d9c170c359778653dedc86848f4bc9a465b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc1fd1be9bc71b561050ec5a8334ceed0f077b24e61ef8fb7e0677f48eb51411286684dcd6f548e6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a4825219c8e02cd26e1b8474c5e28ca80c63c0f79f6f8aa72fdd2797f84940e6320c92701e1ba01c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7759a78f89825f07e4489e4f4b8337cbc25db90b55d8b014f8176b002395bf11f113010a344b4964;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38f306f7c360adffb4c5921ab5688f01c965c71751d79ddfeed07014a6e423a77821cebadcf2afe5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5bafff00066a8ce036b0c2846261b760df1f97b2f6af1f359bd9b8c38d56d0c1f1d0ee1f4221f64c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aca2bfa24c125dc2fc74df381f6e9bbc69834ec55a23d4320329cddd97898b609db82feba2bfc6f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef061ed5818e627e55fb46227538e0d01e024f5dc63de4969a990f9ff572de2b5625142408ecd0a38;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44a39389d2732fcde2370c50b243b53c20c370f0990a53ae98578d5930164bf283deec78944a952c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14092a2938a882ce66cac8cca625625e7dc02f592586ba6ea0ac95818e5dc1e2dfbb04848a08675d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b9a4401e7ae57dee29f4843f09d19a88f6e15f25d5a6eeb672ae74965dc939379ba4fdcad323a65a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a620ca4a105234dd3314f4a4bd03a7c0c6219f0753a04efd6873259c5192fc94dbfad4defc0e55fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24750fbf6bab5b3388d8d6b29def28a890db35ae79f4cae75b73839eb53216c8c2dd741b94352531d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h124198f48b6c839a63b40b702deb7f316cdac564974847fc412b8fb194876d8b11b33dde5f4fabc06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb463cd754177c6e55b54ac845359ebd0c27d92d2fd072f0d17a3c567046d7a37c35bc3924ab892220;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e38f513ae87fa74a2ac40a4a12793421d579c36605d7e83ea9ce20fd728b8ae39bf2770f1649db2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h183479dd7dcb3ebd2e93ab652a0f946b92fafa1af6775866e70119f03743f2be44fc1a38141914ece;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he10e0eb48a9fc69e21e72abf78a762e13723dbbd3bd0f33e18cd98c08526ff8b3a4ef3f4d63253171;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2490648367864cf57ba1cf9b3af729a8b645ec74dddc8a0bf8c68a783dfc7682e00e337e5d034167;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h702d343143cea81184eb6c11e9cd411a78c988530dde52d8ed18638d4a3354108e7960c558bee96e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49e538dc95c302f1605bc8a2dd8645c3b4a50d496d1ac25b4180f8e84f8e6e5d1012d0d55e47975ff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaf97b86d598e4a7c0483ed60f7426c87d06f7c03198e9b07ed28a3059d56cd2044a87f886bdfc07;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha60f253ffd30a6c4b51cb25eb2b0d1c5c7676649b97909bc164f3810fc891de6520c33484f7c6c238;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed9c48a89337436f40cf00919ef90fcb0588b7e2ac65529b10d7afc32bb088704c7c07fcc55eaa856;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f21b8b4096e4155fcb26e3b156e187a33905dad37889a0e6a22822438455dbc8cfaece132dab48fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15f9b0cb691dcbbb8335db62fa623eadf8de3691dd911217882349e4cbd5be94f3339e27a3b3d72df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7348b8b69a258d4d6a37367f84d0aad23b82790a5bb618ff994a93a387386efceb142e672c11fa75b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9649be1e8f638745c2dac8805ff854a60c5ae1efe0be1224e4038d8e7106696b601afa4a42a185426;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13194f190341dec85aff2be15e2dbe03b620c9827aac8be8016d446d6a2e21b20cdad53ca869b3f1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7af323305308136068c65d8462f857ebc0dcc0babe9618d55a225d79ff26b22bc56d9fdf88868b816;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecb9d58133dd596f57b76a85fa4a582ab5a2376dd81f3159c5dc7d2ab96bc34485ae225d26039415b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13a33729a971a7dbd265f44aab6b09f6fe2fd10076813c457beda6a88c26431bfaec9af8ccaceca8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17a5f16a5d553ac72b19ed2ece8e5be1f37a2554b21c690efc417da00fe9d35678ca815429dd38312;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12714c2e2965b99347874602ff26ffcc8654da597c410c3be4ef050e3d2e3ee72884bee50eecdf4eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43f98b6fcc2029b43520715719e3ce9883820a9a4e3d7ba347e5afa473274e51b33ce988b6ae8418b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd11b6b152552394a81ed23db6dd62bcb0fef9f4b36e79c99b4b9ada67a7ac7909e389fa068a047ceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda36f97c274580d36f5365e7f0d7d188ef8b465f2ffb1e09c141abae5d3f7ce0cc8c124c2cd29f0ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf961a29a9a1e60cdcf9efc7a9f39fee945b7ee6940b2331d339781c51497a507f4f02a757cacf95d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hede2d4378969f30c31fbee8b7c2a5bce2d889610300fc9c68820967968e2397eef97524149a3cde4c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd47adfdaf070d9fc8c96d96827315b2f8bed9588803217c40d7ade0ff9201e22351e54c66c841ec7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2567309c41361df464898e1750525d7398c41a64fa5f23e6dceafd12951d487679f12311d9e83ff0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8db82cca85245e723dba6a154186fe928f257f6fb037fe0ba8e0c25fcc002abc096425759541a8a39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h380bfc2c07fadd996821ed62151737b7429ce2c896b4a4001e71945fee1bceebacea0c9b79ce2cdbf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aca52cd16124e17f1a975efc925fcc74346e7112f33a6b74f1a0fec3a31ff9a3c17682b209c03d1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c2c96a2a68a6ee0a6cd0b9a2030e9287051f967635cd47aafb335600e7ea0b5f5c495eda343a1689;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he910e7875337c3a0a47ad6c914b4f84fec96346556cfda33a27c81c35645445973c53eaf2d438ecbc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d77ba7968a36fe38b89a8bc1197695f5bc2b2072979247e5e3e3f64497312aacfab3372ae74ef27a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bf56ee49af68446d387bbff2fc080ce255f7f31c1a0245ae8aac94fd53cef19374ac7b7f8ea76947;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1219c547624dc77f87f0d3d8d5a2632797ac528299c400ed0f2bdb202bdd700989f13b43b5f7b3751;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h209b196953aeb2cce08d88104efb5ab8e36b447cb1776d3667844e075f8d735ede16e5dfbc7a60c3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcd7b8efdb6e51fff686df13e5211208d9bf04f8584c103e3714ee6c5c2c6684e1da1ff3423016983;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6955c333e35d1a60e21e3a7a3c1cb6a1d33f4913835aeeae59d31e556ab77a8384e972edf021db436;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1acbeacafab127a90e3d079e41de10f0e8bb2ad4b4b3d7f9109e63e7a11a6f82448807b408e46819e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf75376723bebaf479c45d7fc0969e6896ab07af9d49484367ece883466ae32f9be1ffc6d950e63c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61fe99e66a300a0b7161252b829ade68fc2550609cdf47bd43351b3d5961cc47feed3e25bf9e6ec93;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df30705813e383bf343c9940398b17f17e2c65112762512d758f8e8b2a70fbc148eb9061cf753308;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4bbaa8dd09055219495d35885e0ed13475104cfcc576f7b171375c3874e9c44fd9ce19bc480f6bb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4458333a5ff9702fcf989fe80df9a0493131a9530f6a6130f85ba1b174edccdc75e2aa6d1d1c5a06a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae91a4af14c9e3fa972aba609acc9e2fbabdb05f6e9335cd8a69278d584752a4974849cf9a0d7d8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac5439a32088d5430e9a350627900f6b7440ca1502934ae7824e023d5c6d83a8f268932e81dc67817;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h653bf2d866fbbb9e5d0cd8862893c0b8e442a6a914c64df19fcc62995dd34fcac430c3831e2a0926e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fc24989326b34e4ee4cdf10297218013ab3bedec6d2c19b3c6683b3855b6c624efa5134629db0172;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ed474c7fcd21f79d6c481bc45f8884b96e3099a725f73908ece17c3646c403bd82d98dc91fefcc41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa6027cee375fee309036b2c1acb59708ebee392c33968e3b4f2dc688fa6b44210e04294b911c563e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a9c52c41c8079c765e0f46cec64b35bbc893193c833d7a6718b56d9485ee567d4192e6a50c487b53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h300b5a2f7c7090495133258ff86455fd6dbb1670a474da704a8801d16e22fba036c3e8e479399734a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef712810f492b1ba94b55f02b73399b1a97a8e2fcb968aeb6b0fb8be416f151cab9876b41ff527f6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h596948d9ad12b91cc5d6a5c00ef124530b7a458ced06c00c2a1dccb477618b9d5aaadff872305586b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65b8c970d7dd972c64b6cd099fc015256061adab02ed68dbaccc1912b37b833396c45b1bec05f5fb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdc0fe7b28e6993a3529c6b987510c988e344ebdfc7ed50ab2b1fe1a612eae4046719f5a76d438415;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5a0ccb24272c101dd22f4d48b4a59f12e38c65536881975005b45c134a161824af3c00da39e68247;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2edd03de341dac4efe5bc6daa7d93fe761b855694404ea160ec35d79f3fc364b3488336626e0085be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaffc1fe72c4f05cb6a102cb52f327901ea58a3aa3bc8b95278b8889c3f4e9d0561e6bf3cf8a33625;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4900c6dc772a196c3834fb7891f27cc9e8c3fcf58d0f2a591d1aa1e06e8dd559b67ca148aa15a222d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2aa1b57227e9c5fe4624c9d9334899ca3ab3646e0cf69ed89e15a4eebe04cb839de3664f1c3961dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3aeaab9d86e22cc17008614b68137b011da889e66327aa5c20819da1db48e78ddb65c43cd29a60d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha455db3b13888bf1c14c283fa26d91b38b0644da699a09584f1c274c61c8d18ffee5b82f2d7a0e9be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h289813970544ae9cb6088285bc178f9c5d40ba4acad87970b610dc75d16f43a446848545609c473a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5730d2d239408024c6e1052754b310f328424052c43705c462364bb2e08e264c1b251a8597369347;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5e7de9a6ea6855bf2cc7f5713c23054c657cf04b715ae83f7384ec7214ccca254e45f9956fcd602;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89b1616f625f5986dd4f5b31f9cdfbf3b9703ad3a113c3284cca0808adcd8732e2896eddf00ed7b62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3e0308cf56b5cb55efe6f7a4dbb356680f7bafe8d29efd652e00122121c513cf0a536fd4b22d61cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8a3dac61534b7391db4b1f2f1ae367d33a2448ce2609ee0d83df924f51385f6db5024e0fff9f7c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6125bdd5de675cf51c492b0e2f987356861345dae08701d6539116ec41eb30757880b26e344984bce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h283853c75d5b4c13119cce2c5c5a2386dc031e6d44c7066585b39a15e89755ff55daaba583b4a8cb4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dca10d9b389996b823c5191f4bb36cd91b73aa99410afb52c2b5f53055853a3b0f988e356bde0594;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7359d8a0a86439ffa9192f1cf0e5506b58f2cbd2bc9f32c0e0ff23f9d93ae2335cb9c2a0a79b7cb8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d09fe01a6b7401cc8f403dd779835a6686736bb354ddc1c3d075604e13fbbdd3f7afce092307961b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7e188fa2e0cc36334600ff710c439342804a2ceebed30b220fada805b2a1a9132402a2bad7ced1ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf88474b93a8bf2b63d941ca2eb8c62c5f3aa159aa0b4bafc17aa21b0862f4269f00b15c9893452e82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc54977780c1c1065b954e140b945ab7db0f3ade312e11765ec9bfc3feea12f78565eb7bdf55bf337a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8ff5402bc5d23dd783e95832b0548b823799dc66c4ac70d6d89a3fdef65f47546d10e368f0b089ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7eef7a46d6dc59b5795f8a751623378cb8297879145e4e461527465310f98291884bc727c0197386;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc557573c5ce8d453466e6f539872511c6dc4ef4a33db94a30a7edaa8fcf81d1d27955eaada7062ac3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47b370e322702cab91151cc2577ef8dc512796e1850f62e2e3b47776196bbf3748526cca2550af596;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h342aa52a7bb9fd3f067414635fdb367ff47332663dbc183632032789691df8cb949dfcf43a804e487;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ccd53113891e6df073f3264c64a25de60373958344b1872e6c5c4cac778bb68dbff073995177a36;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f76e440b74e1c4ba059c299a1a31bd01a46b99b3067293bf778cec4a030e790acc480b900eca1126;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefa73be6779525e7b925c2de2c1522bf1684a3cd602551fea06b6e1815891ad48a9f395a441f5b5aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e8b0f69986adcb4948c9861c480bdfc9fa0353d16d38a43183b74ab866e8db5bc80555d4632abb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dec556c58c26a021ea13efc1f0cae5f164f85fdcccb4c351a90fa8a52e28c88053ff55e4b5532308;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a89e1fe73666b4a3479aba7401e36c37a1550e32069d63dd783a3961d732515ed79b3d11772486cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3a6b5c6f350b6978f7df4e73ba57a20739e4675a926cff70709e59960eaae17990f1f47df7dfb74b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f6867f6881fb5e28ef8794f43ffe4fd8a9da2b17c44c433ff0e4122a78b561f050cfabc630924265;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc0e0bacce88c4d7a3b0f8a54fd7caa163f2aad0d49b9750718ca185d2ce621713baa58767cbf81ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1418d613fe0739a8cc4546843672dad4cf6b5b9816208121d86a9ff09fdca9daf17869ac4ac9b3ef4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95683e18ee67711f3f0fe2d1fc3607be92dd03d4076f8ece8c63d0323412827b6a5613b3377c388d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8940dd0dbf69ee596851db25923165995fe9d96a02138b8478e4277a8234c94ce092ebb6faae6248;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8af9c79a8da36659654690b2de23083674f940f58ffdfaddaae088dc753229c8808985d495a7bc3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfe37b3114adf58cb0f82367edb6adf306fcf34087a0ce05cd6ee8d18d5c889a6065f5f16f9db1718;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85c117127df62a98591376d5a6cc53863e885ef061a18ddef546f6574ff5ea98e3c740fa297350d9a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9322bde320a87e23aed36d00e5855b9dbb42043257916ac8453b56d8013fec79cb9cc3a8704f89e7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee4cb76966c8da7958bc22261c04747b602bb61c5a01331ea95d932db9e9ef1043f1dd1fe9aa33272;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h501c4cf9e146c1292b81eaeee8ab39ca8568253fae87a6a4a6cd84854ef25a6013caa9253cf39d7d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h309d0a222cd76acd8994cfb087f1c7ac67b6c5290f8bc1e2fa14805593cd05664453990160cef42a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfec59ef1e82a6a7f9740bdf8533d6d87b11f1a964db7ae529f00477d602d6886e0c0e0c60908c39e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fbecd83ca719d196bb81b1fdf0a52d26d470ef0ade9cfa19d7ff33722067d95ca13ea646d8be825b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h590d83eba0fe857149f816ad4c47eab138794fdee9aa95cba3399c9e32d4bf9cedc32c90227681c56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d44817b942f6b427dc9fd0cbde368992bdfb6bc7f5c979040d335cfffb854623928c9b55b0553523;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc17233883bffc759b26297ce2246f000c54441facbedb864bf72e86ca19073e4b0035997718d86bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6670948c47bdbdc1f5a77d6b6247a6c7765ffeb4d91cbb8e629b0f2d15d7f346364b5519053b6c28;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73361efa5ab3fd02dea9112a2024a90c0c6839dd617353a387607b51c5991dcf9220b5e1491e628d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h677751b1fb5095fbea51c99a17fc146bd3056ccba71bc40758752311df04d305e8b4515620e7d6624;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce9b2009430ca2c6f69ef268d7837c3babfecd487f6fa9dfcd04c07131500620df837d105fcad9fd9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd09bc04765346563731a8b74a92cf0ed9355306d071670541d757ec11434b6d9453d90f25641934ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c76c9512af9f6cc33eac0f34868c2e351ca02fd534ff3aac5a8c625c7c93ec7a415800dd0ee464d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f51fac4c79057d988bd2a6a825be17659d250403f7b539f4abc8ac745d2e226cabab3c782fd1979f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba4c388d41c23454fac7b362baafb7737efe3cb49adb849dbc269a19c88d57542824291b939e5930c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54a2e5ae716dc19dbe41466f0bd8ce83fcbdbfbf5b08704e480bb24a61a65f1f4898d46b85ec086cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fdfecad5f5509313bb2cd5012ef05075cc06b2297397f7d1553966d037057e70edffbee335beeae5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba9e1985fd48f0edcce171322b63dbd54e81d836cd1d45694bb07af6e05640aba73ad76b7e0a6c98e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b94eec6422fbd7a3df472cadef6758ade493c4ef3e8b60c709b921aa209fce657919668a05a6d0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha78a47540367ddc74c7bc5066dd7956b35b14ef6f6b356ede2d7b7807082605f1d985e54b43d6a657;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ac7de5ee5831bc2a158f7fd1974832865223c94fd623fde633db66f85f33bf53bbababf2d108f5ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he92ffc33b6a41213103d69b39cfedaef9597c6d31fcec0d572ea087ef43060fd4dcc509cdaecb4ce8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96626ca76013ef577367ac4c216d8fc8afbf76a61bb3eac0e602f1a0c132037107f40d6efc4c9b42d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2fd6976e8b6203bf22bcc46db60d4245c8a64325d6fa952895cfa92fe2a378277535715758b3c9f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae6670045de35a5f0ef753dc74e0f7543025f8b3a42113479dd7dfa12c65c7f651e6b5c71e03e835f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61f42fe0a2021435faba31b034bfc3ec6e187443da941d66e154bf00ef1fa1f13f2b85cfd990cc268;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e47eff77d3696499bd1398707a959519a13514e7a0cb76e9b4bf91cc096f8ae7c3ada2f873401f42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd697eb10f7c4297e457183caae89cb02f6c0d35bf43117b3c6f0494806b4a491398de79c4f787158;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f9fc6aaa1a11bd1e5996647bd3c5c8ba9ee0eff0b4ef4e0be03940b8b16d101214ab10312e0f0caa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f00982fc8835759510c072352965d939eea7d4f95223762fd4d3c098ae0ba70d84f310258872dd16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae1ce52c6c954514c647493a1f3fe1967b84d570826149ec2a878fa62f3dc17adfd648a155e2ad4bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3baeab854dea4707fe3735ee584be15ee6822bd1d1695a887daacf7dc1b6d87ef7fb2aeacdb8774af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4daca8ccb63c4f72b8c6871c6495ccc5f59b809820070609e1c1e76ff899cb78c6652c0b79353ed38;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h560f99769e4be3a1f379cef68565e504d7f8d2938db1e020a479fb1500e1e1fb333c1653aa25805c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe26450a73ba0f8cf7a78aee8d330c27dbd9491d13650c00120b4bac6de526e79948f3acc60d195dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2c8f070d3f2085148abbda181250af21642d9344c529fa31c74b74fe7b347b6afb2521a64bcc6a1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a5d51b3b19fe60d6c92e52725e07ef69efeb2680f12d91de9d1e3d6bdf222179d1ec452fd02850a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0d080a51e2de0c84ee4313610b811089224a791e18b3571dcf5b48753ac7e7365593d51518442b11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h451226d06caaf16f04b6342efe4566b9d09be4bb7d192ca790a4295895db89585d22806163b352e32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91d20ee1b94d65ca3d7fd3e90ef6cb0949b9ea58bfc18cc2d37244599fe42ff820144a09c093575a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4a17c1671229332f047413983205504dfeb54426f5b136dde604383350c43591a95c80e741a89b7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d70392bf497a36be94b6ee141c60174df11fb9229cb2ada493a59048377efbd2624c0f998b01ffa8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h118fc70cea3957ad9aa00f5dca39155d998809b7fa0622aca53177ac6e8c1821a5feca9663e467e16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6aecb6ce02e5b898aa59617322a1bc53ce783343171c8723a5a29a5ba1bf9eda6df5193bb1277870;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df49bef7408ef676000c03408cd8a7b3e65b43fdaaec6f3686a49cba7a729589793fa86f09bba228;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h127b99387b43cd5a2e730efa4b84ef45b7ad14c1bf3175ab9fbf29a40ff1473be463a990f6e1324c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h912274124f4885a0e480b2796bdccca5c3cbac58436227143205404a6f4a1d4f2450f07707c3ab6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f16bf4fa43a6be03258cc5edf94f95e1051bac07ebe30b9d2b89d2dedd4c2a80d8a1ef85410a782c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haef6994142870cb6e91cdf8b69579d0ab440d87640faec8f2e7fb0718c8ba56e728391390c40f5949;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5573bb180411e7240863aeaea35745c766cc1ec2fa8ddbb2525682099f4f8b3d04e6b3ae22d0c9f12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d0e34f4be1c3dce308d35640b75dbe9c0ce62bbfc5344d1c7b97c07211e1f1ae1d2db970ab14f8d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd9df86d3814cbe49978ae5d37dbf80ed27dce27b12a5f5625b84af79f3c2e079c25b1d79c77a1abc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3047a43adb267f7850a49f61244335d6081c1cad856e5c5ecafddfa769a5e34320ef7f43b9dedc65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4725ba23908f0e5ff2f67514fbf62069cb534d84c4d2171b9a7cbc69de8361d165f153ee844b1394;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63766a92843a49871ec2034993d85066465e0abb32c0a36e047be0eddcaff848b0c1010628fee20d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h153bdfd4a00222e5ddfb5253317dd6d2a07a36982a9d0443f07c1f9696ff0c06ab0c76e4b0c9217f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc71d4d6b064ad4c78b901845bfea9a24dc3f34641461db07a4ca96625ded1e878e881bcb9c34afed0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c7c586f3650a97e2d667f096e37d085db00d2add5ac97b58a558ea4e438972f91a2d7a328735847d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30bcdb64ecc8c7ef7f3820a831f74c13849a1c3b65fc580ab7be841d70cae3ea9919f69f976dbb9bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h637e37bff93dcc1a5aacc7dfce5900c072c3f29ccb6f03a1b5592e5652d50bb4a8651f8f1a4973091;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd94182abeb295a1e4c321988389677595ce583c067e41fd0fe9f930a64f1c65a5f548ac33350e12a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7e8bff01bbb6bc0a504016080e8986cdbebb6cc7eb6d8b840561e83b2216ed02851904c483d8b38d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a057563a0e49d7e9906fd3ffcd297e32a1f921ec556f5f73cc6797abd64cc6bde49cf83a55f9f576;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce9a99b933d9e70bf4ccc51869fdea49ec320bb606f9393e4d5447799d091c2187fd3609df9cdb00e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0909745610f60a959cf97193da05373366ebc366e186f2f2a8993e3273bc2a092827f7201ad130e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc239c88c536e45607a0615836fb86acae2375b8ee9a550174c32e48d8fc0a2e720a68fdae3c4fe857;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1965c5db472301d0118499f936af0ebddc4d9a472166041d01e41f7074f0365f87a86db9857dde43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d460ccdaf32445f91d328f9828d19b24d841adf07275e9859ef9a4638d5a5883961e7907875b6ec7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6f7dc9f9311fc90a2227e423fe24a865c4cd9ea395dd0ceaca6f8c2af2bee9ed71c5a8f389cf042c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha933f52754abd506e017d5cf1f8856ee2aea3942711330cffbdb9d960bea8337169bd52884cae42e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca916a2c49d6d63f4c2f3c2369ab313bbbd0ce3c613b7f95afec00a1e0e4f0143829f62bd3ed322b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34c27521e4242e9f3750beac967b25be94aa2cc3814ab9427ef7ee8f7339928700d09dc2e33e5e07f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he67834bc053a8871d18ef0da4bc573873e31cb49d1881577b814a5ed3bc943a8cf10aec0a913d2ba2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f0489b9a1bdfc3c430598a3aa07413365aa554e9afad59af523cfadcc75ffd4df086655f63ddb0a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf77d124a674c12455c3f4ddbbc4c62396b9e2235a74fb39e6630447b00c203fd00d42b7373f4da004;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d008f1e7aa998f9c6602528ee4dc04496889f36086ecf16d500d3994c237447dc171768e3f362643;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef2d9dba54d9d70df5bbacd88e2469dbe04497341313bf3eef7c9a23b144144814b42898c0498132e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b9a2d31196842c1835fda17633abf3ce7654b10a69c5c242a7e072ce5e966e96b8f12505e6fd9457;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26a189118520a07038201ff4bccc2690104bb7c9f60f4293c3d936e4e74bbd88548cb7f01cd669226;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a1e327b3df2830da94c35c4e7f04135a64015507b82d2f021210b958f5f6e6685eea5192d557a14f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d55bc230d3a66924828d771005aaed50df63e0da6a68c86d6a17381b3a01d2ce54c2077231bfcffd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h736f28007457fa098c4eb8539982580a2c1472c9d917a21f8e4263d386172090571efb1ccac865eea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2d293f2ffa7689c4014f66fd2b421d63983ebabe4dcf741cf290ac5d796d92294d133f4be52bce95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79ce26daa48cf02682592a8d3eef4cb1fb086780888c6a8284fd6810d1555c80e5a5c20a70c15289a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd81199657ee4e88b820e79fc26eb8d804903d337ec1231c8f34a725578864d091e69d43bb76ed71b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99055da7acc5f7693cbbe331a8f1edae401d626fef5ec0d00de9b9b710e111c72e6ea8cc90f7adc9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde861a68b6162ebf021fbf051e5e28bbca42b04c47525c4bd6ea9dd80e0802796c6d0dbf661ee0d8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31623ec45bbddada44aadb435feab084098b8daa8e13625692829660f8973a24efd5305a5f063acd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6530cf26e976d23d63fd34129e3c00726880de7d5711560948ddb7ffa300ceef3fe572182876d0be6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68b5b8782b3caa9958f4db005b1f298228c4f5288892a5aaab8e6cf58a72a65b290d26f720d6ce667;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h169f75ba3aea85007b600ad0bb116278392972939d14960a89345ab175138b7ae170301e1513c5f22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40f5b575ec05662ec114b261a0f3dee4a64e32b7dd3a44360afae6c0c6b235fc65e6a0531c45ca98b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73a71a9f6ee229d34bbfe85028cf01f52d6eef73f62921a27c512d1c2718c63a59416ced597f3b9fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd05b7be1c0b7009db5dbbd5cc9069a906278197af8a59c372f749ad93096e1007dbae2952b49803d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcea9512a026a0ef1fd74e3b013c91d0431abcca5b3a6ce971c0f486d63fe07675047491110a04c881;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71c4ee22900e47416b88692edf26f78e03a8de98a5e7d28b983a3e665030f0a0ac510bc6c0cf59599;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92727b3a32e9a307efeaeffc4552115dfb20c1c5b434f624f23b16d6800d321dbb5f798d28602b0e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b9cae49c222f15bb0451d027b9abe2220173ff65884feb9a0f27a86f13f7591d0db7a2d022df9065;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d109cda6cf1ee1c0c993afb8193773c7021a0f54e02d501529a1a48cc30ced64174682ac2fb7a78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb0a3f4f90dede7ad175f89050a20bfd488b0b187632a8cad19a95f210a5cf7d2aef95034947d7bff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdedb1c27cc149de99eb8f095f34a212839634b5d2d08eb8fbfe94621d9aa25d5473bc1df0fb83da7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2ca698ec9c2c366fc237a84577973ef1f5cd096e179afe5ff5fc776c6ee985e66a45d94110b91a9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h500d338f9c425644bb72b4ca14f521eb888b8ec969110a0b7c446d600f40c058b386234eb8d9a60a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b01c9fdfdac532f73b501ee50e8409d19fcd378906f9c5c657834bd3d27e538b14a872737b80eec0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h142aea4b7789f6bbbb18f40e55f0bf5c84e917962ab87740afa9fdcdacceee8c15b47a7160a8e0a78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha504ba66ad7d9fd8a94330b299f67b52b5227b7db381354a24a731cff88068af778b752cc6038e55e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddc7b7930cbe80a2dc6c39149f81160d6bc7b6a883c9157aa2628ddd2d13c225f92fd486e3d77c92e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha25622fa22123536accb54fecabe2d05b6e70d9629590fd515102581683fe3ee7259004c7cb865f62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d1fe6bcbeb59be9f1546d056cf773d0101bd52f35e958c32df379ef71c41357dd347e033d9f3ea82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h133b8d345e0cf8f51d7f93b1eade8595595da483563072fef977264e7db6e0bf038a39f0d43cd896a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6138f03f3a584b3658b30ac723230ad265143534936a75765e321e7b440f26bfad77a762dd7b69b58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8c3967eb8417551285f991e36cd115345606e68c38a0bc89d102fd3da6f8ed8087bbdb9e7cc2f8bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha541391a83d33c2b2fb2bb3b0a2c30477c2bcd55151ab2ae25e7915813e4dbed757cbb6be95b414a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9f91e5a29263dade43a3ae89d2934136a2a39604e414bed56b323b013c9cef7ec18b9d8a9d8d111c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c1ee3a1e2664a0efbc4ab33714a6f33bcaaa9882883c7b90edd084505f3fe40abfdb61be9509a3a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc91db81ec3e7bb9000e0979749850805d03caa0940f4bc456e52274c377e103d96d51cde22853ea91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he29b874026014abe3ab65daa99ec076fc637ffe060dbf1a2777c9257aa42e02506cce928333cab64b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h353fb8976a102aafde7e7270de65f274140f6f96bc9355b3691d1c33c18db51d44b4e317c29882901;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8b39e8639ead0eebbd7aa5f4977f522bb1321846b67e6b15702853eb449eff5b1f500b455c464fce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcbd57a83403ceb3a2b3a7272e66a2f1e03ded220fa803980f26360d891805effc0f162123b178274;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46bddc7eff2fd9c7e4be724d060e6989c301234a261770018a604edee998a9c3582299d8c70de6269;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0a235ab09a6252041bc054d6fd0c54325e611acf8a459dab7dbd7603fcfcab0543f16b24d9a2a98f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2748337e0d754fba7290d810931f7a6bba5b57c82a4cf7e24b64b771fbaf23e58b13ae96f20ed4491;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he185f33b23fff4de48ba443df1cb526a48c5e51906f9055dbc6a9945e10552d603be65ec0f7db7890;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6465d1ccee15d54f2b5f8e10c70f12422874878be35973c7635488b522003ae1de9b53d36170e5e8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f8edb2179472152fa1bbf011944acdeac54cc084a63d785d57b995b10ca89bccbbd3f0509853932;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d472074e2014eeb6a3f4c03fe25a6d42d4a3abca23e9beae2e5536381e89ace01e5befd7cdd2aca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7eb5cf65b86c097b2664f2bcf7d2f50b1baa15a28e708bc60a38a69ade7fe92f975bc615f8e0ec1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9953c5056c285d80e6f45de7dcc61c0d144b2ef688f123b5eba16d1d5cfa3dea87164c682b1e27da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2aab2e2affe70829ae88e8893fa34e31f36d42cee2ad7f40ce66996aec3cbdf029142ba02ffd8efd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8a7be19ccc5c1a61700875b67b6c727e71805f73d1a30af9dd3e39bc2f8f5f7a65ba6bf101cbe27c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa1e8c35bc33e187115ba9ad5ab915809bd0a4d7b60e384d465c67d2a9b3fcfe79356e07519196266;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82446d90b0a6d77831c5f4749df664dfe4ba6a4f7ba24d47bba939977d643e917a8df9b124b6a9004;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e7e7c1930a2f9a6cf341b47943a73efc7386e5427ecae2a8943548183b50745cafc498a48d1555c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7409931abbb49c33e35c55436b7ed802e7a7231014ab8334485aa946bf5170c376acf98d0834e6664;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33bd51782062a25abd92d73a6ea2580e459e4b17f796c19a1638199dce7835e0d6a0de3cd1dac8010;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbf513550e3ae87425ad60172a4af30e4fdcafcf2a8b51aaca1835ab4cbf667d1407f600514e99d2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88a66462fafb3729b3463f77ece5a336711478b97d01919e1f04050f6c7a708933d8998c9e8d6f093;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c87e7d9e5bb5eca63997d9fa7fc0a4d56dee613813de21d02f1f641aebd459b2eaea63d4e7270a3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95a72230cd0ff5e5eadc78ed518db730c2dbd3f9ade34f9632b0a77bb3fc4bbd1bd9ad45aff4ffceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1582352327678a5c537f12c9e6ac65887dffae62cc9144397a9216506cda4212e591272b78100d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f0bec8c0d5d1951a4d62f7e0b2bf9db6581dd43f7ed2bee3a79727f3de39758a9560f4d31d16ad4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed79aaa4582cb1e2b0185024f7fc2dd3ca8b47ebce2c0e3a2dd4255a7e9f731ff09e4186d74317edf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b7c567c51129b4719ff1cb504c863dedfd4fd58b345bdf7b2fa278023b1f646213a350875e31a162;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he68a63aa307ba9efac0b63830d5fd4d7b60f101417a26604f8de3d6fa76247fb32abafbbf7da95191;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc211e5b49a4df3419479f25551ae2a292e8c6f4eacfc56eb9aa04dadbf678afb64dcb03cf023cda6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9e548fba6116bc34ed80b705bfaaf24dda370bac0b43969b5304f6cdec8aa854a1ecdf511b9638e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfdd2dc641c49e0e415b5e2ac141d9e3c5b82e3c6a8868e9333ee3882d9870179f199413004531760;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16ffefab4b8d78852464b70fe9bc33b732fe47c2c2fcf06f5724d11275517cfbd5a7d8c334b1a88ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e2a12f7a983231774228d1de383a08ece25f20369203cf34f54170a11cfcff563554a85ba0416e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8954565a5d5efc48e040733a15718550e1acf75646bd0b3838f651cc0620b46255777361034152794;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67617e44b8e1c165c0a86d02e9957f1dbe7ebde86694125bf1424d9221fb61de4b2520a3522258104;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15f8b30d7649aafe7e6ce85e8e5043423793f6106dfa6f35854874dc8d90db1bedb2aebaf29f75e0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9d5197629d33f37c6d24948768367d00723e8b46907f88521c72cc0b14bca9314afbaf1dc5db157c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddfb7198563290c16aaffe37de41faf61bf861bed5ab9a0fbfe4c8f3ffc87eba62b6251b04602fcda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h849758227826550edeb5b99a311cce71e56723a0a8b2baf381e53eacfc8aa1467d915c8a3b24e2abf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0ccede9c80f22bce4e3976dd62bb3e73264bf3a00b2f8c3f7bfd2a67be84821ace0be9c2e980ae23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7ec7ab3b810008c062a14ed661f6c05557eec34e1f2a3b27e35046e03d46d0190ab92e604b557d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c9a1821981f5f573a992488046d8a31adb08e529817e7040ecf6916d23d4e6338bc5abd64f7364d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c9aef77de935b96e64c7e62c6361be1f3ef380360d831803780ae8de1b9542cdb780657702cbbdf9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9266b7671ee038a27efceb36e2891875158d7a3c4a4a7e4d79e71415ed1f4fbc12785ea09ae1208f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11d825496a51f5a534121a0cd5c99ae130a27aff32d31b922b6ccd9293d0e7b7a88b71f91e3c47637;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he33e5484f11f16b6fb82cf0ce759aa7d86e19cb7a7618fc40fd2a6f6ac490177757489ea623112904;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ff04820fe1dd8436bd5e249a24e3999803659e1e545bcf25123d0a1cad32086eaac582ce7467d9c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47935147d68f21ac65fa41c1d4c130b667db17f14294a8753f399ee3da87b93c003fb10408c5d333e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bbb8c20cb41d6fda8cb7e00eb36dafa4b2007a9dfb3a6b198e3d9f010caf02d944e48e2e945728ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3965e2308d1bccd7bc2780c032dbb5a7b60f0832f4e9d2fbe72034a2e8575a6abf34de5863e4ed25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h502104f144336a47b26d2b5885232d3658ab3925f6dd7266e37c3c0c6552264daa9bf0a688fb5d1ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6452599400c2ed9bd43a8799b644a64ec9ba9c9ff6cf0e695af204db74e37790a1d3015036ba8555f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17ac1bb49b674b7bb738804111db52a3b82e5eeb788803b29ffeb281bbf615966ba1240bfab370544;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3b8972dba3ed4bd6a32174a927464afa66a051bf6893edcc13b6d31346b164a0d0c3e3544add4b26;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4721b0e344acc6dd53aa43e1cf2c2a4a8fb4165099b11787aaf6958f11cb06e2fb7d35f4f726dae18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc38c51ae653ba7e73ffbd8a2568f6dfc463eaa2de11dcfd79fa5bed4d61642eb1734c4dd69727287;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2629daf1cc26c8f37d807350dda2d42e8346be57c1b4ed5f469ac1b9472572330537c1e25fe66f946;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb160803ca3608d312c3566253583ffc9bf61f9fe7d92597c18f1beddcca98b1b829d600e9eedf48d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78ab64a4357cb924126059eb00ae879e7e3b428ec734d0b5e5971faa24a4facda16c0bff81dbc7b95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc0eb7010631e5696212df856a75a9803ae135909b2df75173147fcb3fc4124b77732f91a4058ddaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa27b5658fc821122876be0e35af5bdc159edf1f1f849ab304dbea54ca5cac8fd9f0583177c53f279;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0e70b697a83406200d9b0fa0c5e517eabc4e6aba9e8df630404bbb48b119c46490aa8d0135de7f9a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h263464c0c1c7c03b7054f3f9a1f5ae99f2bdeaf6b3de67fac4fab37e6b7beceb8deb54240eda4e563;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd19978a6fb3e30755b59f79a79d1b7e53024c386a9c05284d412c59d1dd345274ed40c7657253939d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d167bf6dcf63beaea82988fe102458f0241143cbaa1d11d5e0968285f14147f64e323e55c92358a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6f04d34b3fb5c3e4495f0bd7bdf9fffc7424a3b4b25aa60e7c0274c1ea6be5ae74f0b8eb68052e78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heaa905598bc56b4ec0af2ad653cb8cbc5958392b8904e92346a9c53f2d0e8e672025bb3fe6ddbc851;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ddca424b3aff39f803f0652dff410bfc5f7c3748c6d0d76e18f797c4d25d490ed9b42bac6f0501cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haecb6984728241493ad60774c4234f28b58f0e8c0499e902b493913b560e68dd380ddbe9527c7736;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38748be7facdd6674d74eccd404000123c377d780f0c4feb34d27d7f6dc5452a4a06b9f12bb803b2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd28962969561e40538aed2f12606edd40f2f4cda17dac1ad98696019846e3bece6c562a784c5718d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd82004e599fe47e5794282d775eeb7674cf3b87d13de1298d13018158db1541cd9723727f993fd0cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5035509ac39c98523f7dde354de3bccbc848083728e89d196b5743be9b10ce4815428e1bcb02c51d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he45a026f8789add009a1f0fe3a56fd3544c6b37d3f30fe3a910c76e18aab2f825118a553df61ce764;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefa203029601543e8c53af2341bd4ba2240d641045537ecfc564a6ef85b687c81efecd8084108293e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda1978ed244dc444b4df52fa881831574f49ac597be3fcac925b7b3634eeccf447e3da6d46a875649;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b722bb6117c6f7c8a5524e44b606c579bd2d08229d1edd273a3c4cdbdd00cb0fbfc0183b245f7cb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd372403afa4747382ef06f9516495741afd03aaedd75a8d9cac4e25499de938ccfdf4b2e34c1bd6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda71a65a3fab2ad631e534af18968d458d381571cb124cd5220be406c831b850d0265a6c905890fe1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71938493bf9243c07077cdf383076598f2ff5baa9ae4e0ad85ba781843fa1c32914187445a651a076;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he980deefd6e5667086c46cb7f0835509b6ae23da336136660623cfbabf1472f26df9c2fe08bb71b2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bf7593050c8ed76a8bd1f1e6858c1511ab719bb6abcf8d029c023449868d5b82f8f8126dadeab63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2704d54750183f372ba9a1825c5485bc0b438eb1e95875dbd4c33c1b7c30e04c504b125fab2f6158;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7be172c2e9ae99453a9234a67982ea19e7a577963bd4c343da8328455a522e7bf10826f2856edecf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b19718ef641ecbce3d4d01e6060e6e579629f87df294d5d79d1a810696ff4d9d31191f4106de26be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5200c28bc6d5429c29a706968d1b2cb384356a0e61eaa01776f3a3f4ed6ee8043d15b10ccfe26c855;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c17a93077eca6d89ebc9a41c63deb8d59fa4d132d653515df424204c8e492e68f075395fa997067c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2fae06a4972efbce3fd172cf849d82a2f6a88595b6e3b4b1e45ff4d068bb3a7125dce079c3696b7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc94fb077f1033fcf3107ab5d9a649d6e81cde268fe1bb28f4b6380b96b16e08400512d3b0affe91e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf81d5beb4e47834b57ecf25569b9ebdb561ba284df0b783c0547a48be5cfd8d2d30529a193e512415;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10b28de870ded78ee8ada24733a7d0d74bd1387ebb454740fc612cd0b69f44c174eb2765068139696;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ca783bb047e010d41480c13a712d8642b7949362a1e05114230513414fcab718f41c8e801f9fe469;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde7776bb1c9a4657c4b6d663dc8bacae7c960e3478660d3e61e69ea974668001c2f3ef685a98b334;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0182be29e8ffa32e859a7acf71b6fb88b364ff346ce2cdcce70fcc048652605801a10a6ebdb40b92;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h121b7e1f2ef74c631188f9e0932211209b157836672f708e47e43f07db13f018e2c43ab73b3f1ee0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40c0f8eb55470a3bc9ea9f0539815c60fbcdd58ede95aea7e53750ade3a78e654ef0098b38f9918b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b10145a8185fa5b8bdeff3b9087f5ace02856bcd6d74a529073d080dfae57bcd13883179c931493c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59ec6b40c7ec9b1f9809607024c7404f4e5cf0f3b7c22fdd85194b1fd93ba52b35d1c2b98d3a237e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bcc29943e770edadbde7ffbb94326e24d004ae54faf0fdbb9839f20c1b09e6f9946007fa63c10f47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha856d3e6dcefc9d33408e737ddcf32a89985a1cb51ed3a2c913aa6ce4ec91737f39ce80f66690b33b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7564056d8b2f29f36733537abba3635001b1a73f664df589fc92a53afd38d086258ad1324b5313c83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd28afafae3d2ac16444eabc77197a1c3685b99aaccc728734b2e7b8e725c97f6a5b23890c8c7edc72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h448b7aa81d9520940958bf501165d9417f7ee50bfdaac3c1b9dfbb2f635a8b5219e24e923ea67cf7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79d489d31e8d1f536539767856915da6831b604baaa3dbdbbb2a0951db44fa402b6c78293320f6e34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dae86f433ccdcb14294fc97b6d5627a43ceee2f02eafb3a238d0ec21a3a06aaa3ee9adeef8d80dd8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24693b6896d1f2658dcd82a33b40cd9d20ba090ff8e2d533844b86fdff5c7cc9b3c53a1c1b4adea24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b35cef8550b3abe6612c66c47aa4a6aa90c8a8fdbc59997a5eab3a367e2fa6aa53bd3b10e4431ac4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6544ddcd1b4acc31eb7dfb78ec45b98148b51ce5d17abc13c600abe73fded3a1a4c4cd1a59b0785a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cddaeb00fb101c33c12826148cc1a84989eb94c4c28d3543d021151da5a02715af629d63cf644243;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ac748cd959cfcbfb1dd9927eda2dc92e64d16081cf0a941eb0b3727b4326f2ce913c3b9129b72f11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca5f904ae2b7e0ebb0c5efc7bbea742fe9e4845545166c057f61fb1cc8fe3ef51f400b3dd306d859d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23eafc2d8c17be79bbe2f4a349855c422e9bcac4bfa1d0a572ab74c8604658ea738f0c5d76f2b34a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h116d6ab2ac3048399534548ce0f8283f80c499c9d9e70fd4352bf4471ff8d72167e3878f4aa33cad5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dc197e3dc266cbee6c22cd430ba191a9b15a79a24a2f2ee921dc15ebc62e12bacd934365a2a1ea0e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80892f00fa05b6cbc13dbe31dde331728027f19f94411c6b89daf574104222a473ee6b9140984b70;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcef288057ac2201d953b63563f9e2a0509057bcf629da966b1634cbc3852f8f47aa660d0d5c69ca2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81fa8fe529926ae0769480a2d05af489dd3e7d1095c295320adef5198fdcb91fa1157e92ef4367fb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fcd32b0b5d2c58f9eef4bcf397d13cd8ef1f109f27cb6959455fc4a6e53f9c5cccc3bcb32f890f26;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c5233dee2ae1c17e26d8d9b432b5076bf4239ff9b09616b49f55249ef86701695f4bcc9918dced4c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f57fa6a04ac6f4b61cb5466ba01731cd2e70fdea217928f6294a16c3eced822200ce3120dad21d9f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc051b05bd6d5f9e3e0a60c52d56195c777b25705ff79bd72314709b53a94bfb8b937bd6b41e26451f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h269d6bc2937479b0f6bfcd67726a9eefe31c3f4d2a5060c43ec82694391ecd7a29a0457eab476e2cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1927bfcb52a702f4d16f43ea383b4e9fbb4864de6c118a8fdd162adb9c30bb0d1a556c059a58d98db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1e6abd9ca1abc5f41d32d7fa16837981f08f07d164524fdbfa7c7cf1550748032070393edb261564;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc90bf8e814551003a0eee82a9f1709130879fb0cae00eef9aff84197b09dbbc7005b3638e1834d34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86e5c2ec9342c0cfcde0a3a1d3a1f4062d7f8eb0b698ca085d4301468e96ebaac18d789ce92438dca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha287269a55446506b100e29c981a7e513c2bfe0ec604c2eb32bd80c44a45138bfb54c119b28b40e4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89d167e90ea09b08dbb067f0b28a2bbf9f80347a2683087ae81a9025db248caeacac25eaf5849082d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he174fc4dfb406ea673914d4b16f4b0ce34d9c4ed2464962b6e94115c85f2413a2330a9806f5d1c6fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7557b4bf868f0924c420d86d31185914193d90fedc0d9bc0fab73467435b53e5dbfbc7567d355576;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf791db806f1951b287e9e0a8435eedf221652fde0989eb7bfd0a0b28d4e8944f861d5104501ff5b45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87e28f1120f120eb261f0e52c483b75c85c41ad064f52cd11ae6e9757eb1a162821dcd740f0ed0506;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he91b0ed4c5b03865af4d34677144bfc644d99706a29bf3e61226e92fa370c8e7fd8c531363e8801a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce54cd53cecfde3e750027fea3f76cd967803adc68e0347852a40b82d6e9fbd5d1d2b7cab7f66d1b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f6915f6ec260e6f4e3a8e6296a0c8c0cc6811331103f1b2fe8c033cf186057639b050086ddcb0370;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h519c9879300e3ee93418f24541d70f87fb60c05edc3ecb64fd4df7a52a86bf77e312b83378ed991ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee72b1e19aaf382252c1b10cc86d33ffb3e414c085972356218b112c61b8f1096a3208dc8dbb2f010;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6abd8c34c2daf8e17c22e09b0a918d59c39394622f4d67266fcc1e423e98c4d94237dfacdefd36405;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7b79690ac37cb2f80284d148db25595c26e9f724ccb75374dc03bfc8a38420986f1fbdf2425d9aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96480328e6ed9994b8794e311b8e0b609c9f7d7fce1f2010c9b9da6e0f5bb2c675aa7e6332a04bc84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ddd0314027ad139328b5ca05a4ba508dd381f54aa6bb4abf311606f304c2c678f2bd3dede73c0afe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98a154b850465bf556473ef44d5f7e18ebc731c88f8033ba1892f6c114948eb68ebb617d10ef80cc8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5cf99535a1ade2dfadd5d927c540ff816684a5b8bf6a097baff03129b040a885891382321a77a231;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc663efc05f3fe4462f343f2953ed9dde9fe630f463bbc506729e0e531bab366ea775dedce499276e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36f86ae2c27aba3023577c5ffe92cf693d6dd713fd68b049b2b5c3a4da354a246ca842aa754d577e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fdc58bf0c1f98bffbcb84cb7a1912994bfff63c684aa9d22309cbf762c2f1d4ca43247770cc41b95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d6acb9a4c31e09d4ca6381b33d2b117c04a01e744ef447e24a35dd6923d5da2741f1aad9c52d8694;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a4f8d651c42285c3ba75d8f7a022d78d526b22d5637023a45a26554c0be9e8f721f36a47d7278323;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dc3d7ec1cb13bb3e617c565e646ca0840b5b8bc7b0eea96694b539d7353ea405c676fc8fa299bec4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h431ad000ca8be116421b82cef800ec36da69a2fe6e23ab304701d1c3bf0b9f90590e7848a24272ab5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a0a5d388c796fa0ff51d862ade4afe5e670d01ae44de86b848a8763e6a6bbf309467eb3a19ff442d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he02ce70d9f6d71c3871b4b37c9d9d774d3934139ec5bace0ac28b1ae9c37685d89c5e26338dc81938;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78b59e5d046d3b9b38ca9b819255eaf444619e64aa9d6a75c366425dfcad4f42390def8c9e537110f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h185b364cab5b11a34962e9f8d10481a8bb7f6ee0ee76ac83c9d78eadeb4dad238795837f45875fe82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42001e6f5237c6f146efd8155ad5d160385eb057cd21748fcb353ebf1913d13f8ebcb56852632b1b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha069250b11df00b1d269ef520c837870113c304a061d259c231939c7919743d27af6d0bb67e608269;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd6d9b8f2faf22d2c12b40b53988383b4730a5ee153642416b7660bdc9bb465f5a4a262a3a6d082fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda9a82f99fe9f13d6e73bb97a98346f1d590d6b9119f3eaa0521988b6eafec267d4565603b2c2a4ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43c9c75f2329e66b3bf6bb299e6db7800c73f479ce8cf7ca53a291a34721086d37fb61f7a0cbe95f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h281d5b33197d956a52d215a9be428ed1b38b24a92d924573b66a6c40eb214a5e4fff8a079e5a47af8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec451e501b1376b9927807437d6624d6bcc3b3e79f28f65794e6016e4972fd751e99abc245e503f44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fc02289803def68d3fd7dcfe3a8740952003c6cd11cc730a4e48cab4e15ef435716801bcd3095737;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62e329872d1cec9989299ccf2deccfa7d13f5eb860e966b725b354ffbcc83cc8dd5e8bb6f9c7f70c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49bdeaa786024a8df3c48091470026e5296434862b2412d67d87ad1d3f0d8970d18232d8cf8dd98ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba40ac87aaa1a5c08417a65dc8b5da07fe09442e9c0deb25d489c3b6351c18b8d6478a66c8f5f4791;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a43eb51d0a27c951d15850689319f42646793558e441bfe2b3ad29127cd205998058a8cd51b8f9d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ce0716a2c0f753762e8f53513125f270f4df8f7b47e43f1bce0ab3738cbb71f9b69d6c3f72df7d37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha193e13fa4db4a98a580418b47f160b783ec60ab02808c8e5a75693e6e41b5690d122918fd5e89b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8426904ed7f8c49803a4d86d29e1bf958dbc335bd2210efb0273265f037ad8ff921c447da3071bc0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24f709a737acaba58f842cee80047346844231e4ed17037fd61e28dbbd15aedfdf8246e6267c940a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f69ea2e0246a5b430a819271de842a7e3a8e3ad7fcd590065b09741fb02eb4ad0b6221d0a3a8523a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ab324ee94f7006ae3ad0c6d007f36c7831c46d93c91de47dd25e0cfebdfad992f99697c5bd14ed4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c084f5aaab06b449885274cd3e562e4fa548c38ca95db1ad779c71fd36cddd77ddd2cffc3890addb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2938545805324c67cf9ac2f21c7f849f58d8c127739815cfac61d9d82ad265c385730a6ca2d967946;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h181ab2102fed7f0aa515205c739da2ae8042146fd868c2f7ff3055c1f19c9f3a4959487bcd862a7be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b5b9ebeff29ea924eb3acff7034b5ce20518d3c3e69f0707f2c7a01649f36483cf00b478002dd729;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4561c5f12ba2607028e1260739a480fba349f44fc8fc50b5b6e06636f0e6e0c6d4146b837b141fb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca48a4d2ded9d5aa0c73596c7f2e2ededa117fad8ec07b015c2a75d35ed771dee1d9f6a6cc6d6d73b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cbde7c995134bceffec569b78e36681dd3809d5834a01825526ef980198757aa12352fff71fcdd20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2c080d0cb3178366901ddee88e59da967cff358e8cab57b44fe344a99d2c058081e1f8bf209aecfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ee2498ed8e5b9c45b10e5b36eda99e12aab024f37fa6b5cf4adb6ff76bfac984c17371c2824bbd1c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h278e249d2820ee4a11eac31d07524c6da0bbe6854093f54d9dc6d9402c61a8ccc20e5b32d932c7803;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0054f1a90b7f4ed74d753d1c2a6ec15704b25a7a922187963c6be7c2275aaff8576f32f3339058a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc1af58986af5192699edef600ae0238803caf6314ae1adc54d8178558bbb38665a56fb19a8c5a445;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb99d1fb37625a694c2d64e5f36b77db1ac28f9be6e0345a698b1d3bafce2dc2672cd522d3fea66cd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h102ab7d9a4aaf7e5ef3996b6c03b49a582640f064ed6aadc9a40317a7ea7e07caac16bd0635f86a71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3c4434a73aad61c7b916e545f11ffe5b64f8a00270de052d0d750f9701c79d6cd52c96b9a29f015e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94fc0037273dee5a42da85e47e5d94c9780e3c9c962dc4ce09e019909e035da7f082f96f5084c5712;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h669155b810621432f78aaf54edbeea3fd9caff761c78c3f2b3c827330f1ae3f5c15a3baefd9f69dc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he87184ee8b3bf21bf4f72e3fc958cff645bf3bc2ae1ef2114d9811bc31442dc4075ce1d79e8914e1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fc4c39e44d47a96beb9e3c86fd2b3c5705453e04e4f109ef5acb149e7dc9aba2a2b97d0e8e33787b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f895ef91e4cf01d8ea3c2305ff5ce89b60ac25cedfbff5c0913dc3b0704c4904598e56041b6c89d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39bf609b4704cb13c130586f5554224496f88e37c0179db9273c02c17ca50dbc131b71bcf375d2874;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51052d1edf618d1dc9d9b793b81ff4d4eabd2b338b9abd678edd409f3dd62b1e6cc1bf702597c5dbf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a7cf349ab1fb8680ee7f88ef982233fcdc22e75cdeef2c9486c98b643dc868c9b3c284df1433fbb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44f03eb0e578232df346d2d8a792f37e6de71f881a9a3abf7b9e61db6403533dcfaca5310d902ca2d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h544b17b00409c4ff4712e6854dd8c5332ff80e2be7144bc5605a0f3e99ad6a11383ab0084855651f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd299e40293b9f359760ffa352af9e3a2fdc491dfc1197706b5ccf4d3c60b76589feb2c0a452823bc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53a5f169443be3991df99aa2c8a53e75118a47c4c6142b32089da458b9803309111b15c9472bfd67b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6e708ed2172d8eff90b30ec967996b816aa77c1e267a14e5bf3ce7788479ff6bac9fe8327472da47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd3b778f6ef02ea9bc6d75c423f9673ef38ca956bee9ebf5ac8726a661912c1ab37e11786af4f3fba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h115511431c421e21329a47f8bab433bc68b8635db3178d596e5c6b3fe6a80d00674baccc571848b8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe7aab48c0c0372e7932706b1070e8cc4f8cb4c832ee68d65734668dda88dbbb94b2069e0bd10f831;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha393ea8218390edeea28ced8ba90b648698c2b28fee0a69f061c113c19d7d23384ced5996244a3ddf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf836832104313d47ebb10031b95da599a3b133639e97ce3e27a4c09fbde65935a536692d793cdd206;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd07fa88caf9e37b55a81579718e4135baf23baf562f8d2930287aeb6635f192698ad64b3f4faab9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1362bb649345eadd81e58e328edb4277da88f40308e40828bfca246ecd28bdd53d40a7b32a1d56d98;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h295b015c4839ab72fb0c623c0d8aea84b99409e9038dc176a8e06bf884d76bada1153c81e023d3b40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a0d5bf23d46f139748e17b56493395345b30e6b0f76991cc27f0badee8d79d244576ecafe60c31c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29b4c47b391f279b461e6aa80e2de6103db9b104bf80ce7edc3a89a47346693061060e6867d617506;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11632b154d5087ed231986a4af5f5bf0b655bef038125a78ec6c566abd6e5d565b2ec3e0c92fc80eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6b22d2a2122c7e448ee269725f1f26affb83430571315e43402f42a29dc918b313b01986503c0eec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1012c30064cd6fa2c28fd2ce1373b481dae66bf58c7b11184e4b5b7781f1e18d8c129f122df0844d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f0ce92eef11fcbd95d07e8879ab0c92d736f8a734f30e1adbe6c26a864caa9b4cd691ebdbd5f29b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11ba2b57e04cfdb388ada7192837cca34c4c495ec2e8afcc5ecbe8ccddb64211087ab1c6d67bc464;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf75d36e191d6f346c64d6845493fe1ea9a1fe82c895742ac971142031ae4433c5267baf9ca008341e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8942d2e9ab2c6e66ae8c1f527b071a3a8e97e367b1ff3b2685990903ee6ab40ba4584d51fd3323477;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h995aeff2ff03b42304bbbf9eea7211924b77655cdabd9ed41b3ee90d680a0fc03a2e95c8baac8e164;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2bbec61234d0f1581473b389b5b1102eac9ffa2f2f6f073ecee2a5340bcd685c0f1dbe6cac04ac48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ed6c02a697510ac936b0eccc0c63e1ad5679cc66951309ecef7a96f135298d0ac0095e975f105f42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c87954ef0d5d186746ac38db88c4ff316f9424d3df9beaf5e12f7813327f4eb01175ec56d5cd9431;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9e8f18f772c75baf035d65a1b1fed044cea42f1cb21adc0f095f5c81f7826c0abc8f8f39966c93d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d9ac969b2f5c1c8022728ba75c1dc7e88a5b0627b3d508f5db7eb8a95a584020c8363e08ed8829ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h242755039f022856f8a977704dc3718221b9742d62ea10d1dd5acf962387d7a26ddca0923ecfd3c94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e753fe221502cfb1aadada7dc4f4b6e659310c360f5cba7c3818bd58b171826f59322f34f6d8e3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h393de041ee32756a8642ca8ea994a9fa310cc02462acaab3c7d3fb57966c8e70858d0b9ae870defab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a35809d53b96d26a3666edd804aeba9b88f7bf5337af68b5d918fa71ce95bc939f050a151002c6e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93e921b67b320b70829be261883fd00f5d02f9b6bf7cfdadf9faa3bae87c8a7dbfce0b6d2b628685b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dd48495253912b667095fbd7e0c3fb7803580c5240f9e82870a1c9eb24046d1c3ae829dde0d3965c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed3962d66dcf1c81556ea991a34214659d96cbdd3d653f01351905cf41e9155495c1d936fcca57682;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had4ffc2299a2984235638aa72217dc4a070e40b9a4cb8c606e23e92ce188a3e11c0f61faa8ccd618b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3973d98b234695a7ce2ded10c1d5e1d00a98e861462ce4992f1d70d7659e7a57d8cec1600fd5bf913;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24037daa1910784f903a3fa724b214e561a0e46f6afd6989e6526464c8f4ca78d8a28ff00501c3117;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5d2f2c81af60784e6c4dff57437b2e665e9be11ab3c3e8aa96c7a0298ac8f9699c91d4411414da3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cfd517e2a942608b22c42a9f3569a38e724f738e527b841798a49caee13553be56d667a8bce73a5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2045e4f45ac2b937faf1c7f7d298c74a1088ee41884f3222811bd8f09bccae3548579b856955f677;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce09af003c9b9c61e5e9edb313643e03e84afcbb21a550ae51070118587f46530e510d4b95c7fcb61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37be2548c9428bb05bdf9850d5f42e6dc3b2e657fb0b303ef1718cf139f800a32bdc420c95c7e47f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc172594087f2d01ef904c52b13a47451fb187003c97f96b41e5daca03db4d897fabe7befd95d450d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d4482cfefde4e64f34978db2420c7f85d9379088920d532e787d39324a33dc9cf5872ec4d6148f61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82b5bc274558c8c79337b7fdb0ad9b710c0f0ab26e8c7120efc6ea4ed025a15be1c785c8a6eff5788;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fb935ab90feca451acf354ab67ddc0b7dd1a2b96d14a6217919462f83c2cb541a21a9b6681cc65e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha16dd303be800273b7ea98ecd34fe77814f0e95f023acd0d064a56d183c2ca5202eff67152086d90c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5accacbbf28b6979e7384131059293162d2f2af12b10e09b14bf11ce8edf990a8c1965f3c6ccedce2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa2b36504aedb73f40f917da5499d5f9bae6fee16e0b730a1969d657810db016448d4e29eb1e73406;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd17356c590354dd354254bc2c6394ec3a356e6c827b4b134cff9a33dc3f4422cb264ad1f049134bba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ca1a089d43624c9a80423756ba961422fee0e314b651aef91ce98904298e84e644e51a1dce9ca960;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5bf2157d61357b1ba425b743d629530151a20914638dc2a0ea5f3f24c8e229edbe6bf3da62166f48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b77eba4b2972ef90760b15b39bc96f6bf4571649295cb071469f86bdcfab9a19b124262d7d7a5fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1d508a16f34793e4145b6fbbacea79bbd6165f617061ae30bc1a44c6710e2de2a22cfd8edf165a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb12ae762c73d44c0c96b179e5605b2147dbff69ff8cb4d245662980ddf0a738a83f88d8615ca6ccd6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f83cf2261c75fd13924eed0b20fa11817097abbee7bf87ef4cbc98fb0509752c3bc000b1c919dad9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac16d9cab8e7f687779a432ca6d56783b6cc4608feec5af5df49778c088537cc092f8ee3d85d70f34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1a2d7a01dc21f50511bfac0092c75fb363d4f2a20b85947d93731b525ca20ce315d2d8a3e481bce1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h601ba9f8dbf2f3cd1e4729816b1be846df8c927e7a3db4fd85cc7fbe8dd5df250ccf6c5d35449ffa3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59f995a60245b6fc77663bc3c0a3999a2920b55de2705b6b4fb1617d0582b5c389f147d4f6bf997ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf21f89a4be5d0c8e62046e0f182e056a110a5bcb12f7a9473b8297d9d5aa30d1ee406376811e8f866;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfde8309097d34a1df17f57fe170bf76a2e7d4a72574d6303f7fa7b234f963ff8ef63ee0eb303d7897;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h843e21f902c3e4d519e9d9f165064a512eec95b83ce52735553181f5c1ca24e594a7ebca773f28514;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3a02642dbd581083ec2e978ea0c1e0c15ae59a61c7e6d661ee375f9a431deceb44f50d8776909a44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h695710203195ad510ce994156b35e3e4b9a2490583e5fb895895de0ce39968a2423cdf9bf15e252bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d32dd2eea9358165170602e8e36ee62c36a1f902361139b0adb3ec4d2b1eafa561b6cf0d4ab8cb8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbf65487f1ab62d3f5849994777e39a05f1744e798451a041f142516f5f54062bf66729d685cea86e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c8c9cf07ab621f3eb664ee85ab5846be4f1d418cb456e0985d91aece798214fa8bdfc6723fddd658;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51baad7b757f2c3f6712f6c180f7860821cbf659d159095dcea07c9a8aab87cb6f6aa155b26fe3184;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18c9bdd7e60e68627d56796323f305fcc8fc85e83ed528a172af2f50280675d8ff0fee1341c4a2f37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h967607bcda7a95eba6b0d055214c9c055207b2f2fca035156e2c99a6c9b8aff3cf7caaa2fe3fd7963;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d9ff09dd821f91ee1f6b0a33f75a9ce4bcc60c1a5c5433ef151b8663a57c83bbd4ecc1360e7f44ed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18a3036788fa5af3546d2ba9e74a8f945d5de331786ce9d4b46a3cea47c2abb573749be80575c3b82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h714aaf4493088be82e4868c07466c37e29d5db63c2b0657490794c95a19c60b16440127480356a790;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf482ddfa952293be3ac20cd0018337b1264d631c4b78a3a6b03c488b8ac8f2e2aad90a90113f1958e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea8bcb33f4840eab45c8980e2fdadbdde9ed091d8dd81df4b746dc852c674d9cfa5e8eabb639cafb4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h455988871fae2ffcbe477fd48d3d05fdd31a06a7038693933431d2c5e83136387dd2570cd9002d81;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha66950051aa1781514ec9e94251f08afaa2bb12bcc1316a9287fda014afbe3071273468e04400e265;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61831e22b606a2144da48e6b8d2cad04e055bbb262c1c9086f58726970cc78be110b2bf141ae650e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c718d1233a53bc1831b1e1cb8b5218b62a23476b087deeff2e69333a3977c937c411ad39640c71c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7971c031d75c749d9cc3c37b8807026496eac0d75ac5e3ddef135b693993de5cf214e94be54133177;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2f6b93059ad2101955bb1f7073a6a9e2ca3cafa49f975ec903b170ac9ef0fdcdd5cebf505e25b418;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde3d3e653e7b2fc571e2bdeb0c5a4e615ce912c2fdee11488014fabfc78bb3a15461ea5698baf123f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47f744229f4ef3413c70cbb4e053e91da13137aeacc97cf3368d44b36888d87abf0fbc505d0f168e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b68625c22566cf091989848561a8af28e884bf7992d9f18bb2c36fbceb35d9a7e8e450e39ba25fd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe8e53795b1a96a860c4119cbb81513c59f2da44d386f9d78f493693d799a2ff9190698a4982afa20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he77a8b5499ae8fb8a94d4114963e95d70484eacdbb0f573a6f4c2a5977bf9a44e1079e98108d5ce5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84e8f2d0e46fc884c8767ae4225357bdc26ed66928257f5d7362d6d9a293b2dbe0920be137c69b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18bbb49ff175a84e052ae5ae0d04da80180c09fae726254eb7dd0a6f06f7e88179897fdce92809e63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf44832d6e45f5b8d9e1b1f0e9a8707e8329345125311b39ef6dc749fdd10f373e4d9b7ca05f22d0bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3110f7811ead59f202c388db7c6fc540fbaea5aca5e4bc18a96375825e74d05a16f4ad87258099bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51448099cc6d06f6b39b40d5cc68f69746cff5f2010c2f06c0f4126dc4457fe15653e34c965689ee7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb79630d6b89efe9b45010ee0632d2c5a7317b5ea1fe509b1a32559ce592707d16b9d4e045044c63ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1bbb1e932e1a04d742e7bd5921117243d156b55cc78261673a1f4391c6978b364f4a2b5f9a9c29b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51f5aee8de187610bb353a435737f23c10299bb3d6a2cfec99afbfc029a2c9a504b0523c7d0cf866d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca2797bfa42709c461721e71e10f16e7db8a62951e449b79f0a0d3ef90cc8c6cb440393c403d442d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a3e81c3a1f278089a8bd04f035e887370c36d4f2c2040724e7c5448914fe7308901142d9c47a1797;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23a515c106d5c57304ab5f04b72e0d0a47294415a1ef32de918c72abc183dccdc0cf4f93910747261;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf79aaae314922bcc93a17f79a15882f13d63801e10ec21a7b737865702d24b6444a118682749a5da8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ac4c11ef144aea0dab1bbc72566df4afbfd957cd047123c8813d696bbce5a6b60f458a5c59844866;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbc466d6544153d00f6fc061c121cb6d3518b3a92310faccff7e4de192270cb44f1ca471084fb7736;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9f9826516bedbd3abb360a8111e5f05d711201f83ee352028e87a0f2ecd359925d000edbe16bfe5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa75ddfb88fc1c59160bb5a5daa0c286caf5051f79e1cd37ca0d7d699cc2250a1b4e353527d7596a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde31ce015d0540bdeab4439031ec618fda1906a5dd3c4ed7f2089e27429070be580ad7bb226925a61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8ec135a2c8bcff797d54a681c69c06297e01e5cef2dfc0881b6cb62ef4b3d99518ae495bbfecc849;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c3fba8a130f4cf1cdc43da9e9bd0633b2543dec9c370111141ccf0d2dfc611fefe20b8052818cbd3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58280d2d4226d27644ed710e2a89bfa3d81aa9ab0a73831b3d50106ea7b1625417538a35da05a1e96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32a126cdd5394a9f9626b27ba307c6a896625c4bc0f7e60f1dc01a6d25aa052af0a6b0dda0a24c780;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef5ba2bf0426a92ae6c57c7bc595258a7cbed0b22b642d02455f0dc29e850ebb0742f0bf4f46f9b0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a142a1ed3916f4290424da574394f7da2b07e3c05c93107fc476716b9c3b615928e04ab8f2aed7db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had77c844862a9ae0a55d587db03732dba79bcbaaddde82fc6ef636ac436435c72c8f101abebba1a47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b81d8c9bdff0416778cabdf53ce96b98f3abdc9873b26d3a4a64b2fa9f596233c95f305f91a147f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f5e4663b87e5bbaf5d53c161b52bb3c63324afb78ec0cf3d0240f647a3d45f6392983599b60c9f39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h805a610f4a312663217c8c11520e8a010468d425c9074fcb140e5ec14653ec05a97aa9aeea5a51bb5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h897468005c562294c51c440b413bef61214c86c6a5ee581589d7914d50754d1268627fd9621b7cfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb2ebcb22f461fbeaa96b3626cb2840c89ca7f1a6460f080a49c6c7da9d12c6ece30e2465235aa90c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66dc67d58aea13525285b16f6c48dee29358dd918bfd183535d938b2bcbf57b90c24032188efb9a18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha00cf60646448b26360491b737c77eeffa0fe98bf0942fe321ca1f587ba4b430b62f894d853e6c794;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7df2e039ebdbcb735fe3365e49da0855e9c7c2bb99f28b6d8d174f0348e338fae181cf3bb97b43ac0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a8f3e8a25866e19ce48369b63b1f60ae703b8f4e24e6049d70f94a37352173b716b386c2c0238866;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff377d49d6b216c4b90f21ac06a6ddf38e8aff0e51ce09aed44c1fd5af8e9718fcc483e541aed346f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18b2a019ead05261f3ec7ccc68e167a1aff5fec840f68912d0b78e9cbb84e33eab81067f87bb6cb22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbbb6c5968660bbfff74cb9d11e19cec177b288d859d876490f5ebb61d39a048ba955378fe48b247e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12fcefa973a8029c67885f22ee7725c956669ae150506dafd2cfb0ff673f516c07fa209e071073c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h760f358250b7ed6c3c929f1f1f30fe79c08b2cf3537951675db684f9d43794f7c0ac52fdea65d0156;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h610004263ffaa7c80aca5832cb4a615dccfc3c734983edcde9a2d4aa4a4f05416f95a0c5f620db3e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85e13184bdf11d5d243165b543dcf934279d92c74bba99eaeebc024929e0522623ad2a239ed4add21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ef13f6660096f8c117faeb54ca11a4f940cd2a435176687358a41f90d13a4674d64a861591fb2b11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fd58adf0711581daa7c59093f158a61b817565f1b1b120b9d70327038f9a822d9421ca343d6d353f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ef1ef472b36c05b18212ab87fb7f4ca1109127e2499c5924984def6b5effff1901c6d9dbd7112a25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dab38d10ba2c33d7fb19da4caec95ae1b8764e1feb5386ed4c76305b912a82e7840d4dbb7a99f650;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8077f99219eb1ebd6413fcb439f0bcc776500cf046a421e3abbe99776e64f40ccdf3306242c360d4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95f2fe71e86fe60ead0e3405566edf4ba1a844d5d7152f1830b3968e9f12fb73f034eeea1c8b3b80f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4372e1d1688ea7a8087850eb26d0722cd6ce7df0bc633991ac6ba566c3e3312d67cb1407d5bf354e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6da788c1d8b617a6374ef543c800e0c319ec35b6b3bfa3862d1cd216a9c06bc0e4455619c0ed83b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78c1c54466e9e233bf6c8d05bb13b6737aad1c8e250a6775bc9f31da9124bf7e587282a4426e4ff5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bb02a7ebcb8128120a832eaaa68a7da9f8a10a1bfe638fa1a5a3447f8a206b4f9649cef897ada83b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b8a8ef7c9c906c8e5f1da3537284a259e6636f3aa16da3f63872a893e576033aee0b771d43c605a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h439adf68d5683c90e035448b7e8ddf8aa3cba457cc81aa9860e6e175260fe76730e236608250c4f4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h180c9b348fd5866cd6a6a3e04084512897d18e212095a9c59db00978fcf6c8dde700527289577be59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62acfb4aec671b44923de2c9516a60dfbbb32a7f079e04c9249d590c8ce3dbcdd4c9edd2646629981;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b8ee7b1ee441ef82a347646f016c721a8221b1318d8d0771fa7b47169ecd130eedbe34ef4418d319;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h225f50905bf22f70e55988f3dbf25f31073c4569dbd1f94899d52a5f49e1c3b8a577d04cdb0c1d363;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbf3b36d4fefb79ea1404a18332ed74d0c62f82201d16138fa43a27a336e9032acb5343569aecd0a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc32411bea1e29c706e739ad1c10a9b9d7e3df35a3d8dcc2a3fa4dd50602ea11a1badebad32c1843f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1901a45884a2e6dae2901d4d89444d9ce4bb3b071f2d8b56362ba265215f9042e82f60a1f0dc6e621;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab5a1dd5d4d9bfe5b914275f4acee64d02ac6444216111fa4c6be6932c04fadc966075cc5dd218108;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7f65115fabce853b33f6f7aa7e347c8f9b33371d448ef28342d3a372b37fa4086829aead894822a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h326f4efa024ef2f9b546990ae6a45a537fd8e19134e193c29a5c80f6fb115d6fe035ec0eee64eb437;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97546d541d530372105033731941a49a7a6bee711edb2084c123f97db5412012348dd8a92fe62ad91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f7757b530e590501fd62b1f912e1a77aec1666c7bb550e7bf403ecdcba2eea604870242a394c2c3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbe5f7af4597c8f58762bda6a41f8f7e3b43ed01bf28f41f465bd8b02c0ed67f10141e111df23a5a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3ceecce957fab622d1ef8f1c8a7d1b47c7ba8c9df3844dbf9e74b73ee26007db2509ccb6601583cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64482fad07b7d644450226368b51c7cde8384c6a36ff157f80fde351a9bdd68e796d7dce04dbe6e1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6786198e9e7055dbd12dba2a547f9ca71d90056eb4878949eb61833ece12d4dbd055f80ed447fecb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha93fe6ff277f613c51213858dc56c80e32cd42dc3cd324bbbb0ee5c82412eb3f46cb6beb0ebb771df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf52e1080fea09586e792d2920f0f9c1efe58f9ec712a74ac26b628986e58148f488abcab68954f1d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30e314b7a399dab2f1ac6a8a6cbcff947e3f250b3b7c126ddb22474e6b2e416d4c5428da9bae89065;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35fd0d2d0eb78e5c02eebe6994f2e18f5b0cab0eaa4876e2f4363deafb7df3754bd3196fd63bc36cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c127d53921d3d300239fddedbd6a0383d767d675053cfb6d9a065ea0ddf717f6ff5e76f8cbf0f277;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he234559ce2531582332266cd87bf081cf387511b455dfb2d3581039db6428c5b13716e6671ca314;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a421321ade71215953443e7fcbe91ec42db4bfa8d853480aa5992d771bd07f2bd87132f6263a5aa6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40b37846f806de2078ed9991d4e30c4fc828b015ccdcffa71899568842ba094d4a676496646e2d31b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ee9d1c37354e8c55af14329735b0499322dbf65aa36f33c7c4b18669385aa51ca1f0aeda70cda14d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h294c15d0b10c85052389e9cfccde08f89e3f1dd367f17bd8d4cbefc41a08ea132972dd9ca3b98439;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0afb908b91950e2da588118306ad7f9be780bb61373d4a44370258157ff27db8239b36176799d2e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ff84baea8ed4dabf7e1bc615e86b615d9f5e9c56939600caee6db1f254bf51c5d12b070e28a665e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fbc230e7d46446db0527da9710fd1f9209638ca65874dff299e39bc0df80b71f11c0c66618ad531c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6491b2b9055de4fd461c505429b7a5bf967600195188837d8cc739a9200cd3787da0be2bf52f35c51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecbac9b521e14bb747b04c6ac00f08a92790d5dd9713414049923e8cc9d93f96e6d82cbfc75d97053;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7e2dc08b96f03cba65e19a02d283cbde98483c4098f3ac24f3f348c2ac490ffd054a3fe5acc984bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8110f327ae88adf8d99d0fbab11d5a37a0e19e14f64cd442a58dfc8e385358e28e687f21851a0080;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7134246575a48054d1c8211742be599ac75e9bdd4e4711ef3ff164676541792568905ba16122a0c7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41c9737064b9b01fee0a68eb5f5198c7f60d569474e285161d3b807f60ba8516fe7fa0d9f59ae1b1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcebd895e725dffb7c49d3dc735bb01d0ff794cbf6717a4ce7562c54943d6a69898307209a410262aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f116d97ee024b63647b0b5e42cd3b5f294444a890e19e27569eca892b89c301a1a2311fd397034f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75a569dc117d7434d282c37c0a97d0fdec321afe6bbe9cd6cfd88546d8d35d189c4a6ea18b47123d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40179d686d2747ccb4e01aa79d2c7f4b4da34400edd938601df81489f3535d72f5c51d0422ae95309;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e1b1bf8b10196612405f08e9421a4b20372fde6b645e221a599236b1d60edd416eeecae6bec8c306;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d73771092a13fa625cb6817d08fd61a682392c699fa67829db7cec9965ab51a87faf35460b3ba9bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedf7ade9b8623c7581682fc07ee024ecf8fb3fafe0d1f2a230c04cd15e2b2e2dbc711bf7d54689f8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f20b932b1ff88910c5a779ce783e8dadfac9930c6ccf30c990d2de24611938b68ba3479a109bccf0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6389fce036c62300ec9d522254f532eb2d3b8d0e5616dbc271c79f9d211efe5eb0646a2e46f3fc76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h527cbf4bab20f812cbcdaaa0337e6ca47087ca3b3e1ee207f7688deb3fbb3bb0973c2437991d9926f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h825ee2a64e7fca1ba0b3dc5e91c4d9a862630ab80ab50910d1e28d2f4996998106d82315df424bdda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2febd90556b4ab61cdd7d4a1da73dfe3373d6f925c4db231b2a6abf55e80f1543a8ca74bf30f036;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb9e1a5363e96430dbd0e96af70c80063d02961bb2dd9fbe2881ff759e67dcb854201bd0978e8b4b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a0b4d10443943d661a51c6523d200e42d49c5e3c0793546e13a120a7d93857fb7a94a9d4619f8803;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55c5d5a22a50117e2e1dfdd1c95f20b0ffc0212ddaf5ab8769a38dc5c0c21b0e0d56d0ebc728c7ad1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h772e52430640ca5cbe62e0821e6f07a4006ffa1219d4487daa7cf6edaed2a3e8261f95599a6489557;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h957dd9886debd0d5b1cf03fcb9001e7ba335e06fba36b96863f1a6253ca0a0e1ad7174bb22bb7c81b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba1007f7833c3bbc47ec33d0355d18fc3e67f38e210b8e401af14510e2c0c746f3fc091eef2e080be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb93697e8bc70a189b34b877f690b53af01e5baa64e2484e33c7731453b0986fb68a9bd7fe7e5a66f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb33279118bf200f2d4011db4a24e732637ca60ea063824bf412efb5a525ae1f7da3e9bca69f47332e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca30f1bc0ab7ddc1d3e71f5667e98cd223b397b65274e5cbc5a22b32889725f5b892cc3a6ceea6263;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h173c0c155395c6df0617af200121a44de110787a13fa76f69eb52b2669801507cc3fe424d9d44b3d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he087ca945471063b0db2337eac5af61833134fa02bd45488b639229987053e3e48344b9428cfe2def;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc88cf4f79c0945fb21e86349556579460439b5885f985cbdb379fc9776cbcf985129ad8fcdd8b0e1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf7fd78b2ad327bc9dd6478a199feb6653ff378415ea37fca4470377ee5bf70243111ac72022018d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf3cdac3ec40b9858acfa5d18084b967b13ea4c4477693f2df0622d2a689e1c15f350615543e1624;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9901cfb062b631f908ea18370f18c86f8709f66a70ed7f6e0fb6ab58a44740f8ff2733947400981dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e26f753bd0e31bcd31944e23c5a30c878860ee79bc967bb095037ffc9984d216f6a8da620f320f09;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32a949dc958fe6b509f87c9c684cf78f30ae5e2a394267de39405b9a07e8731de628a0556c2acfc51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25ab3082648333f88b0d503f618796dace72d1ec5bd677e00ae77a6e28ca2c07e4321449f0cb82047;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fb471283800be1f389071df4950e87169d05bbebb4fbadadf223ba66fff09d031276d0015afb26bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec4e744cc9a3bb1c6a1da758a47a919a1a1281b8e432f8ad93173ffe6db4d7c295ae32123dff1b8f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb55a8b0aaf285b1adddce547e5771a47c63c0412b94d54c595766c13988a094ab29012f2fcead0292;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc5f061831436fd98ade1bc46bc5005414816ba710faa6e821a47e26c389a2969259dcde8e7d2336c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13b9bab1e42caf506cb64a15089906e329d4152073207a0953ccf31a9dcab4813483453021937878c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5de51eb27553db14afd4567929fca61625d92e13241e2068ffb57cb3a1927f110561a7e1dafde7642;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8212a13c3947b1cfffdaac94db12be4412e0a735e83757b187e1a47e57032e7a949c68c226703c9a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e35b477f8ca40492ae7acc17164281a16c31f94c2c215a9f0af974e80a530fd6cc1ea9bb5e239b0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46e519b15930c0fc7a9f25aa748d80954b7ecfc95e9d36568ac6d6e4924ffe4a5337594a780527663;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe397776e34c359a30341f774a42f9aa91ce407ec6fdc9cb521a17a56337c74a4bf2754cb2bd580f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0372d95abd887b0578c809612ec0207846632b5eca96ad73fbff15debca5325c533b5be20a06c4da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb23c09c7a34acb365ae8947345e0051dff66adbcd39f7f9abfc4eeb8e9c32990e6de063ef9038b9cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f3209c3f0e7c6624ef5d961f53d58381fc6b5ebb2b051c6ca71ed59b5d4ba2787073cca1f1e5337f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf44f7b39bb01d683fb2c3dcb79a37e6d6e01d0f10a874f0ff1dfcd12438baab72ab1e4d76d5fcc916;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e54065b580a947b18f3ba12cd4aff990d36ff983a5b030ce541ac850f2db48b566db086a1e0f4ab5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12bb02ebf63796add6c354c5b18a53f476b7d0ee0d9145a8395a2b1df75beb0dbdbfcb65e77250d92;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcae8a35145e8fbc833ca2be925bfc979e99247006ed1fb6d96cd330a8695c92589bb4cb1fe892bb54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac946c762ecb35395bf6907fe7f262face351191bbdc1e15c5b92f0b7f0180cdc361895e02cb2cfc9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h210ac1659856f5e5e5de0ef062af30a236efaf6f5c64f4c2696ebe4f58d68a4894647f0e50629c814;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e40a86f925f6adf3c3631cfd4c26de0a0e16ea4cdc54f22598a59ad44a4632e4d642ddeb0e69a41a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4de449cad3f76291006337ec1cef6f29d2842d0d0390cb951f4412b21c13c6f070a68ed9b532dafe5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc822b109c35b558ab120590027024c9c4cc2864b378caf98002f1c644414e4eafbfbcce64571a098b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40569ea590335d80945870559171c24a676b664040c72af636dc550590bf373f06e3f513c580079f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7e9864cde3efe3e85867b6db719d9670b95c3756678afa4bf2bf18c0f00ac5a19c8ccb15ec0beba8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0a70a650820c5412c2165c0602df8ae722df7ba65e5c5b2ec25e13ea7359126666b05bdae9115511;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42f2ef78e0da4d1a778052b3a0a9001e266bc90ee0378c6530d9e47ba22036ddd09f88f9127da7a79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2f35b1aa7024a8395f89fedfbe1ac81fc1f697065a269f45acdcd05a75fe5d372faa2f08724ea106;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h576129c8cb84bf5c382311954e6df6446354eee4592bd01840079c385aec26c3b962eba193d0e99c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1b4f25f5b7aed9f17abb824ff61dc336960e59ca32fa01481c210d704a594050dbdc489ec1295418;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h913c02600d34eaadb8682fa2da9a3ff9e4fce50a27b9804fa98503876990b504019dbb210c9300197;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf10309bfe7239c0bf37388e767dd26f44c07329706c76aefead222695f74c672d505e73b9a840fbdf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdcc9c8b0105ab97dff242df13eaf8a3a3a473ccb538faaddae4ea095e26db6db744475e15daab39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd051ec7f957deb5b8e6c93bde1eb6d41200fd70abb23dd4cd3cc60f3ce490a13f7e1cadbb050b3482;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96ffb879e5b83a28892787de29282ca52752134ddd5efaf0e4680693e7b5b6ed5b39210f15d22b19a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4006c43de46fa5b6b8a3eb3368d930c7f824ede77f8e642857dafab13a6e67afe5795cb873cf0fa8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc890887ba3dad816afded7172bc698d27c068780fcac7fe0eb1b68fd32196873bec6f848ad55a3bb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h974fdea597b3dd9aabd8666f1cb3f31edc6d78630fb8601cd1688e697b1150d914cf661b0ff04b249;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h886eaed1fd6f27a2d228c76e9e8e5f82348a926296aa91b7e9cbb04e07e88062e7b079c8acc65fd1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75e98a7ab2f2e3bf1908741f140648dcd0e90049bdfae2f6a6d9b1f44b7a5991c11d1147657ff5cbe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddcf167a7e45934a964bbe21b066f402bf07b8aaf98170c18e460b5df48c4bb596cbca4746146253c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h974fa8e458e2c5f150ae956ee595a950d63165cafe5914bb654483307df47698e6b7c4ae08c7b8300;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ce8d9ec3bebb8993ae34f34d0f8a7b692da427862a75382c2f231710c5b91a3b5de0ef948961d92b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h566221e0e8b9601ff5d079874e4107a93d1ade817fcd394f88e94d00b5130d9f0b64b291a182d8621;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77108182041b90104742081379fa109cbd9a249cfac5a2298ae67c2fff2e6e38b82796e61d0ecc25e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda51ae7c8334d8926b2eb2652ba12b843245c5630b8b9f4f7c121ac15b40f0509450548f3e9a819d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f4324ecee05f181070e96a1d949e6e194a5cb12c335912b7b2abc332e4e06cafe38966a0d054aa24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb317f9716dd277894d45cfb0eea6be794d14819d4e00206108ac58de0566fb3e98db043cfdd073099;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc218c4053c61a200f6a1c3276918e83161c49ccfa7a0179d0fb79007648866b8809ee53aa906dcb47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeb45bee5817d0c7f32fd0f656b217abf9188ed6ee0670d28551a4c5e4026e46285a0900847a731dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23ce26048ba650b46d120fd4c8a18d59689b1c06e8cbf08bc86f5da6922832008f0c0243f064f846d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7c7fe28fb40b418da52b3876eab4659d8805b9ec34bf90527e832533a25da59fa5f77820d4f47950;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf843a6ee89e75e119889f15d8b9466a10748a41899a91a6fe13517ac4a0d4b5f99c985ade75d3416e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6c7d4e402238de3ba8e50cbadc94a106c8e6b76e78582c7ced6e08296d3d15fa069667f7b0e795d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1030435976cb7532528a9d581e02e4cf8646168a298bd950263f6d25d143fb22c1109a554536cfbb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha93f9c4e72c8c3c3af497971a9dd95343fc7ec314f73477cae1776889ae5b243e9941b921b1a435c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9fdd14d5f57f4f7f6723c9c74c73d9125c6db2e90c3ee13c11ca03eb581116c3717cbb27ff8604b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4d7ecbbe208dcc688579cfba3e270c6bcc988ac59c5204cb3fd2cf2ba159a64884b6a4e45aab4ca0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h231b88f222267ab72bd73c5ed25e477339f2f3a1a14d0697c68ce3c7d4a8457173b33de1ca975c38e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a9964f2a16f8e41a56b880335eed323d7d43103ea4598b7e2d7435b43f6402cdeda82635618f26c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h973ab04e1369df8e708dfa10d8fba6c7034c6a0e9d9d63f784d9f50607976fcf908b6b39834b59da6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d961dc2e1f2359629eb5e11b911a729b781550970b899000218840f452af25f6581ab1c557c9d064;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d99bd15f8890413e9fae185380fd1daed55b477844acc7757f725deb6478714665f949b4ec14a2e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1d9c0f2f2127ff90fed4e0ea693bb05945306a5318aa378583d3f7c0a075dcac6c0ec2e4dbb91fc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4415073f90fc90d548b2870d9046ea2ded3ed5962e6059e0af85aeae569b0644dab8cfcc0ddd8ce10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c0e27f594087b2865ec12c2483f4df69ce86e34b3eb94c8a26fdffdc628f0dba3b870729bd2d81fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h482d64defba3b326bdf1994ee6062087fc84beaa7cc10bbf82463bfc9d44ca2956001df2f7459310f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbc5a2d37504b2d0ed8663dedc12bcdd403f75192e91c1b345594e78eb58d0bd3df7b56b3a6496f29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35a8523e826fdfac518510ffbbc56290e1b67ec621ce88e5bd57a1911e2d01fc8c744732d6fa7e1c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2989eb742c66215374a288bb02e768cf108b4d9de8c19dd8989a92bf97e678071ef31cec8319013d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5ce759cafa0f8d8cdf3aa8f6483d123f43c40ebf43e5a240ed3a98d2e0d4fdd0e430d5c91d59ec5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eafc2da3d26c800742c9386c613e4e5b7ff28b9c0ed945ac8ce16eb4ee3c2cce70c5af7aa48b7ab4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e095425beecd641b7d64f9a009f48db8fb1849cb48944970eea27af50cc8ddac81d2b520a8a57e48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2d7cae3b2c62f3cb113870c127a4c54db7d1452f1742a646d12d7923ee927e31ae93551b4f9df0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf82d48c6e2e16b8d816a704fc1b811e20a1642113705776bd0daba7ff463b8bd878f733b7132761f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ea17d402b94f5966bb35ed291a92768422e0ba292a3287d24cd1018055976a429ae372e49d7c1e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0513016328101ce3202243ee52ffe9db82e0148d02e3d4249bc122a87aada3eb2aad5414bff7e155;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf30392c11c6d6b45424eb6755fedf3ddd7975de19431c11eaaee0c391bf276f7abf2478a6762235fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67d27fd4eaa5f55bb2b80c9c7bf1dfe117f5e60f39f90f4e5a3d722e1c3b79023ca939c9e56048eb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1a55807700c0698e4511deb2b130f316d0c11ca1b3e3b83ab448756b9cafaa855c398d35f7ee37d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13dc298d04cbf27e627ca11adfa2c3daa0c53b75ddd4e7b05c2e235b43fca26cb29016bd2db5c5e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0059b25df1630692921d769bdfcc035b1cb009629a7c7e9b9444d8d3d780961d1081a255dfcffdc0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81ddec158db0c1f749b06fa4157227632112ae6ba7baa411b763c4fdf83d2479bd0db195a3f0e3fde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h657feeebae6e91cf25b93d067a197a316bef3c2480e1be0fd837713c2ab99a9b7b5c647a7fda0958c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f0c126a7dba827ca87e44dda56f70f7c90c020be3949eca78a31e704ad2a1a70e446337659c2b4c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef2e2a4d1905e890ccda52f1404eae7c102de8edb2c810c8a6a0953cc2d2d95ca8b476dfa4340cd79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3620b792c49798bbc966dc168f44a110c7e69214d670423a660fece75cb4431da56af24b22e32187;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c8fb2c1e1f83c04c96af01090bde206ef3937953b42bffdf9d1dc01f6522d4d41ddbd5adca64b79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h995d1a5a5652b122092d24ed6e0328c4490250b9363a5c51635e7a4f95758c063e025e77e1882dad2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1a2cc6c10263d1c6aa073a53cd0f08f3bf2c49c668ac5355c055dbba20734b240334eac7ddd343f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68608ecb480d8fe2a3be1e24fd82a4ce1c7cfe8eff6da331aadf88ddd505dff2b7a65e15b1c9ff8c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd2926d410f3f38626211fec7f58c4cda6023688e216ae2f9a03696ac3787ed01492a41ab773b4f48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d2fabdf05f32ecba969bdd76f74c7b5fa12915b5125db5e854b1db9e82af6dfd15ac3d184e69ff5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47201e11a55dcbf3ee48618e0404c7c98f0c950849ca1d136173261e5bf1822514f8a4582b79e01d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa3a6305ebdb8b9edb1a83dfe953ff664d9c80ac3182182e9c7dc642246f175db3970c9a97029751b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h423236f561ca786e5c38b52f9660ae357ddcfa6fefca9e4a06be4978b6090c3c2a62aab20f241c78b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h563426b942d543973a403cc138b087509cba205ec2375506ad3a8008061e30e7c451acb17205ae6ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b600e636e3b1291e15266b4f256077c6993ebca92cedcb922325a22a9d6e5b207d1e0d117a1f01eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89ff991bc786826920a6ea98d64b2e9dd6baad5067e4ca490d957626fa7b5bd8ebdf4031f0e352cc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ef5766b8e7731b42a9ac47c240d087e547c59fecde56fedf25105ef2ae44b544383bed32410295e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44092c784b591efab730719d3c623d0f989cc3e7e2f3da1ca4fd81bc6c1d00501bb4b8c19a8f8287a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73e5bd8464e9e6a6c46e4d2830c93ac4ab060cfc7c25c3794a966478cfa2939a2e9bc53e0d32bc384;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf54171884339c93d96e84350f99ce88e603a3ce31bfc269472b853f9c4740231b11780854b3f4e10e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bb39daf8bd54f42dde16eb31f803da290e2e95856431af88733d21e1af74b205ea591f6eafee324a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57280009e516ace2a3239415f4137240cb38880a755ce65d82597ce4edbcb7fd3e0dfd349b493e295;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c39828376d8286bcef3555559e096e793d3b6a8a32135019da11cdc5c62b9a24e51cf3fddb3eda82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7837a99e4351747f68b10ab461fef475a9de87c7f2a42d4c13c8b3fb011a3651c8dbcf4149daa045;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86d651bafb5639d2033213f94fc45229a98bf14f995b8f8c6f2584890069b13d2f2e8e8b1e962f403;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcc30d22b795c1beec1a1e78786a4fdaa3d0b20b4dd9a6540b4c8767ce1cdadca70673bf052cf2700;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f7bebe7d68c75387505b0413b3c45fec73d8d0b5827998d46763ee59ec326145971290fbea2ed962;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c04b19aa363be626d73a0f9c406961ac59ea2f03f41772ccfd36c7dc3e2d2ed99a5e1c782819feda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6f29cd0180beb7e0a4a454597986d607cbe07117e5f86d1ade8beb9f0120cc6138c47a8d551356bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40fd7de1230680c217a288b918fb1bc7b8a8a39511cf46ef616c3949edc1f7663a2dcba4c4e01ee46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4437e08d8af732cab8b07783bf4567674cefa1e2303bfcc7a770722f400365d5dde47ff2cee4fd523;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h797ae1ed73733fdc81cc446f17cc7970d4d37279cbdd1b4f04ebcca6320647acfa3a61c98813f86f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec60f6d38f744e3b5e605773e3479ca0b3a9f9efde656e4d95812b304fbd8ea2d342a4b09063d6461;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7ac289c3da4bfd9eab39f2c88ac4992731bed922a0c707e2ccae83f80d9390e119d57f55f42ead5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8805b8caa336b5dd74d545a0f64bc726d4b8242047d6e2ca6b54a9f73cb4c1232bb2ed83807abf49c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b469f0ce19cb6d68efd2e5fea8739ad6f815b961a41368dc259081165351e33b9b3742a71bf2c07e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9571684895bc27b85073f5c533d4b43201a5daf68e87b28247bc41e77d98fc717df2ea7b1c2af2bb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80e12f7781abbd2de1fd42a4126a820491b9e5e3c6af77ac4ecd9cfc9c3ed58931a9b16d45cbc7d05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61f06fe3b1333cc1fe2cd4387560140e8bc47897fd6edca1256c40161a7b71053f4e0b9d89466dd0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8697fb41f2e8160e88cbb6d0f889b76013b23fb723376b9fa8750219bc949994ed2a1c999b5b4b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5227ad5f1036f6cac194ae661da6b8c2bd4e8381a8d8ad167c7cca3615dd15e5354962ece7eec7651;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43c41feadd90f7827135309c57b43a8cc2c3c6ef1b430be2102272435e898702049471b8e9cf0f00b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h493f9ae30ca13538825196184e34efdd6e93343856ecd7b04851b8e1a9c940bec555975b288d6a0e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2695ac733f684debaa2f7b054789bda1175dd48d5918e95a7bf59797033902fbf31b6484e0a8845dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a9a69e54d56d42cae8a0b990a4366e57b684311771e422ebe91ca5f71478e9b4f7cf45658b1bb7a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h750616ed39c866d4c95a3db8c5dab4497dbc1bf6b54da373756e1ddb53a09d12c6ce0d083dd04f09a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f651cca7fa19124e243aebb081827e80a3f09c28a52b929759505664159f92d177f78b4bdbe9af5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec3d81d6e41d88689a30b09e7d8ac4a62b88efb41a4cdf0a51dfc66239d517292e33c2055d3157f6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee64a240f475abf185b340e226c40648e3fa6b2e08163adc3dd982d4b07c5a06a00f5d306fd400f76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5c23c3372b5b5379268024ec71b42b5c8fcbf38521e3c35062a0c275450b0cadff4db6ccaf9f4708;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h571227bb8d597d278f79e1f765e4abd6b6516228b0ee8f96de1d13da427fe6aab49dc2fde3e4bbe5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96358c6ea755b5e4c5c30469fc2a2da40a978b2f08a79b1b094759abd49aba1b689f0d83e81fbac8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d34d7114a70e30e95df7db56eb854d4dc38e7ca5ea8565b06bcedb4ce20b409b89013e1c18ee93c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d0d73a82e87224290f1c8294fc25e28192862a2320ebf77e2106c7d11dcb41f922b433adf00183b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb62118021dc7424c5c05cdb8316f318b8acf2f2b21cbfd9835366d2ef5f8bd7aea6ccd515d936ecb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h633396e3b5b260ebad680193b8c6f365c5f19fad5a3e9f5ca6b5fa0c863f74ec8013f04cf097b71ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h997eb82d555307f79feca761798e9a06a971e72f2d528e3e1624fc584c2f5894d97306c92393a0dea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cecf9fc78081b84e175ec11cff20ce6ef5a9f9dc8337b426f8981ffcd0b7b939aa218cbb4c206ece;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ef836ad9fb93e998337cb5c5bd058347adb9ce79683e4aba51519d46467ee6b8347ce3987ab4a575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce162972bab77b225943e250fa52337315948f174d0f5695b90eceb302228013a0c23019955a4f3d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6a8b14db0ececebcd64b10c81b80ebdf6f529b3fdf18187fcc132e91ba22ac8d1dc4e241c87de227;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3347fabb4da78f5bc732b9c7c972f0cf91a427749c43c3b52ae99fc82927c51a492be6243644a169d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h283f11afb7fb05c3199fb9064736949fb55ed1084d13bf6f8684671629ff6d7572b90984af37be03d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f06855ba68f4fa36677e7028ff4cbb9f8388682a547439302f2f2825033485d34bdca307fb776c0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7370e44350a965184a7d15ec495732f157256ea44d6f70d5a99ca6e9ce3043efc953468ad686e422;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6167a3691326c414ed6832bc0a41ae8b483a2ca7faec4a17939cb121437ff5e6c26416fd0b4c2e01;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h546f1744ac5bf9974e179ff64affc0b60a8cd8399f0c1b2c2ba8e60630a656e3617c2af09f09447c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7fa8e790076fd26579b1fe8a0440d9032eca98b5427c9951b135c98e99b65b7372cfb734c8c5ef8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e825451438ff05ba42f65cab2bc31e9efec8f016e1fccbfcd09603a47fb80ad0d7ac48fbd14b9cab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h690c3f8d6d4443ff3ffc062d6c41f84fda5c08b11138934b645d2a7de6f36aabab0ec38e81d60f05e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be010c47d11d2f9b02425d91beff4d1c295a95cf1db026b4de5950a2e39e558d6b450381347850ed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8caf9e363a58dda82cd3d5bbc6816fae63ac11519a3209a93c81d00fc616f4eb87d59234447b7bb89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ed371c61cd3d05a3c359a281ad0930a9491ee9347e9db30dca5a64bd38bc7830ebd68bc5e67d534;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8564828a9a35ce2718b72d1faa021140e9b69b96b2acf49d59019efa562f20040ab363a394d057265;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaf0cca0bc007c3fda7b07e29673c1e2bf5bcff1c56813e4da2f2c31d16a82b51cf72a847ea7fe86f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52314452f23abdc4a33ff54b7d2ccd754217a0f0c35e73589b97557ca74340e5edb7c97251e66c3b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9ed6d953079067cb3800ab307fd26d2647f7aea0f0e8d93588d1a69aa6398ca8836ccc4d0973d957;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6919d469da4018023ba6550e2053e62c5ec9a58251660f31322f55ba22b2f226ff6778020d5bd303e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9f48331b88bf03100865f694f4e5a95729306fbda4aef14ce127631bee1a63f846ced8cde964e860;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85e2273d020dabfc498e5221400284225806d796cb22db652957872d408b711dc7f43329ee4b80165;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he88bce594b52bb150de3673d2c17a3f7ebee42c99eeac8235021757ca62d4923aa184ec3342fd2453;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91044f0d2bb1727b6fb4eb6e4c871399e7847486ccd75ceacaba596ef5d072c7f38798bbea64fb765;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c9f1ae66ed732b4d1d79a3e3157ebfb5f2d5694f791ec0bfa92001d8a9d95d59770dc368de28ab68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h335b843e662b7b6aead50607dc45595fefde2d620f7f991c6ec909e369beab5f72a222f83cf533fbd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b22ffa0dd8964ff3e49205f0bb42f334b73583db577ace1d4b40b62e93cd00216b1db4e7cf89c73f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h180aad07dece646baa31ca1fa863b7193937118cb2758762eb82a68eaa93d73b7c8b7e0583afa5421;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2901b8be3706b6228a90ebb4b8498c4627c4af32636b5a526d2037967a4145514533702fbe10709e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64f7b3edb34df42f77c67177289593680610d5dd9998b92431876b049ce7d5a12c50103e11bd56d2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h330a8c998bcbcb9286cd1311539f3d458dc013d6542962adb12603a8ed00c62d711e2c811d4ba383c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88b359956d6d271ceae11a473748ae7e653a00b333b785f689c564f15e4e0ab17496da2f1cdbf245;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4952b94f83658360778cc9dbfdfad203219cf99414a0090b2e5a63ea96dd0c79b7cb374fd6e752576;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca74202ca0487a62f6a506cd7424c605f6f419764842abdcf7e21ab8ea9bdeb5eb4d8490431b9bb84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc37c00bcccda8130f5ca3503e914d7429943ec53bb9cc590c516f973a15012bdbc41a68fcfd124f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc5aed76f17e935907186a1738b600c9d5e02646329a8268e0ca0594c14efe62b8c23ca4f3f1f1cb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3606d8fd4dda472fe865d4efdc95e7847cc1bf9e5a4f1eaf9b442e4c5bbccf332ec3c534e302011d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcce493a1e9193b72acf92f14c11cbe052b8d5c9e98d2a8ac31cf31fec596ad87b614575586289f16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd04c8dd3f308625f9fc9c4c0eedfab83b84f5956dc5984888abc6af2ea0a7f64ec818235a5781bd23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdae86c609dc4623d073f063d77f8f3202e7de75f3f44a2606d1cecac05ceb1a3837fe228dcfa0455e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddccddcd58591f832eb9f56ab424147fa261fcb64a4830fa2188be33ba9a1b4e24945333d5b22e9b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74aaa5aeff9c72d35d0422b6eecdf9195ada6dbf7fc8476706c65cc8492b7e9b56bbe932a693b4cbe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7329bd5f248b9817e05fe2bce204e04b015f34bc5d15c37364285ab0e1f556af9aed187603f42c014;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9729a6e3088d8e1f97e446556ae89f430d15cffeb8775cdf9dfb0c060858064bcba452e99c0246913;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce9e8abe624d1b76c0445a08a43f382c387a28ffcd17c59af17005f9d07700dcbfe17aec8d04ba4f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf45aa168c44bbc1564d894548e119ab741dbebc1af394080af750cd69cc591252b1bad3cae725f668;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9443b1977e75e96b1062e30b3ca5a563c89367ab9797fe8a49d7a016ec871bc539102eb44b628d513;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h674b17b4521c7443f6e7aae4cc8eb87e761257bac41dbc1d7ed53f4ef522fa7c6325b2eb81134df1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfa4e5a386869292ff5abc040f4faa0ddd9645a7679afdd086028f10f3d2cc04e95fd77d25ec7f6b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65ca9215542eec580be949809722dd0c7aceb7cf5b563777777bc29fb76627581c2c4c7edeae34ec8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ce3b8135ff003bfe16f829440409c204ae2d2482a6eee52f8cbfe5b06291a1a2c775e448b82bc8a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd733f0d6519677b646be82c8a87800943a5dba69190967c0071224ab079a1d96ab2ca4363d76feff4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6d602a2bdb1c5e5b8a336747536ee09e82ba00c7e51236b20a44436a120ddadc638373e1a42e7760;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h366540f07af9a55917d60b76627d6a3399f25e9ed895a7318a4a6645f0de3320b7712af9cdbc6395b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha49ce39b86adfe766d299694f689507ebfa6ec68bbc318bdf83d53c588443948be2118b5d89e0f3a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4de1c22ef0b38267ae892d630b67faf41e4a06ccda3ff00c8591d39e905edfd3a9649bbb29083c1dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h751adc38f29f8c2e18f1da04b8d537cf62a5ace7bc9a54d8f73a19c50c1e7f2f5eea775dd24dd6b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3121f8df1b1f241289d75856f5c38af0e1e64dbe2a20fddb5ae5a4e9a0c8330574b2a510b4078c400;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b598019d061c73ac1bac2fcadd79619ee38d04c3eddd045790b3cf12c4148719976e54ad5074114a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71edadeea6ef4a5ee949d70ce10272e1eefc1ccdb541c4864fc9a7af65449114e3391852c043a11f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0c22cdb9e00dd9778e734287b7fa07a30cd1119e9a948934701ef35d0490f5be1c46d429cb46c8b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b071584ab1e3c84d7ee542eb193750221e0459271d2111e30cf2db99ac7a20e8e3334adb568149ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76ce2c21dcea52828b56bb2dbc6d283537d1385122e4b70815af611f2509f71e58a1edf8892bf63d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h852b33f543c70c10dd93a7af6a36c46a9df72fcba46a1af43de2f451e6b8c180f452dbe40272402f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6411dbe5f25da6d70e23689225d39e168156615c96cffe8feb916c7bad6ec272a7180b29dde54abc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h480b912cf18ccd5fe82129a7ee4fd2528abca2a66897a400a09f0eaf8e2662a283a1f3357ae1d0607;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39ca5a596310d42968c396a4628f4bdacdd3ecde298b7582b7dc73d38927204a53d987bab5381e3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48e09ff30631e47f95b46c031ba55d27251bd955c457d935f5a9acb0b8e7d1824045f82ed8ab2ed29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77216bf9ea0d3d8d6ae490725ef31417d36a5dde5f0d23d0201bed032aad7b4c944b334e616219636;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he64a550a3b986693488c1e4cc8662717a57eb5dc0593b2c9468f6840fa4e35808e478146a204aa04e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef7d7c7da879f8e6f63459cfa13ddef6b80999a76506ffe03042d7e1ae1ff3cd809022528e991f455;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15c25433081853ec6abce45478f7c3aeb7d11899f3575dca13ba4f79f549afd1e103c08293040d16f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6ae818a2376bb24dadf2206c13ec1f6e8fbf998ccc7ff4cce702fb0c6753d1b2b89673c3ce5047cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8cb1828b7fba8eb8cebed688a1b5783eb4cffcaa8a6d54d8fec3e428199e64584bc61b8d01802c756;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bbad069a0bdf90bb670fd1cf74d562ccf4239d61c487f0d401e74f2a2a89179a4c3b0f3dcc72420;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2dca57aae680b7955727828cb067821ccc9249b9b519b93525b036ea9d16aaf28b6a72a9003be9c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c2474982f3faf04f82a48e85eb47b638af9e438c555b29c4afb114d3a9efebe8c57ac6b2aef14ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h138f09f444a82386e0b708224e5bb03ff5b6db1ddfc5d8fadf486399183b65cefe3e39997c211b6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe5923da57589fb71b7bb8edb2554880f0666e58d6aeb86c350861bfbb4b8fb072dcb2f062cdf7403;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4c5882d432b11fa0a10c69059871c912228ab355af3113fbd27bdb563338498614b5101952232750;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha64ee868c7cfa7a13b051b12cfccfa4320845c1ccee3fbf8178a992ea624f34a368acc219c6522174;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h269000a5b91fac981d7287c84bd3e8569b13b16727c155e0dd10d1520ded8453b42f077e8f9de5533;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heec8d397c222c419f8b5e913843f0d4fdb9ea7d1cfae1eda2587c4415e090e68d99f981a2b10b55c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3796d3ad0541f3f8a444f0d58b895625b21544d6f99da45a5f0d19a589ebaa8ba8cba4df779e4388;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23cacd26beaa2489364c82fcee4bb30bfb73bb398e33e8609cfac45e53fcbaf0c3ec348dddb19a6a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5b5d5631715658d99ebe32ebaaf0e1727439c7283b01bf35827c84fdcded4ee891ad9e8c9783e924;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29f9d5bca3d823e3073b5b40381753aa34bd654e1ed0b3dfae516439686eed62b4a4e68d424225a97;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h663928d901766b8a9e970bf4a611f7454ba75c93bb439d200943b1d8a2c7fb8abc4d679957abbd972;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h672d31c4473baae081fd4d67802f3ce31462c74f34d573ea3595fbd4371cf6fa09ff86fa8222b696a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bfe5800f535076a718e05bb373418f6830bd1c855de6fae6fa66a10c69c63d3d3251f1bd9deb0412;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23614304beacb8cd62f4e78dd8383f036ed3b473a26ccdaa05701246480695d4948d17acbfbddec64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha382aa670fb815caf9b7b5a52c84101ed04403c7fa81272b753c54570679828775cee607afea7f5a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7764f059c9a84d064e76e5407de0fa6c1b2d76e11d9e67e1034527507fc1f253ec28a6ecab111382;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ab4bd3db14f092bdd88738d4242453d26b11ecbcf52b35b5e2a1bac14c984255bb89fe4112815461;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43008a1372c5a3b8bebe4b7f699909800d0189a4c16c145f5fbdda3f4ccc36c31f223a761b5c6aab8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2050d4810fca3143f53a8b222d22ee0c07cad56fdb922851c0e8d17ccb56aeeb7f05b1b2cfe8bafe3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1754e780e2c7862ea8fb433f8694e773da5e91357efeb2de73ecd02ece7e7db0785286913cc63262;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h533c77f36e3a11d60ae3d606ebc6fe7647e33e308ed5c335481e161bc9e41685df865b351b95a8694;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ced0d51c743b22a95472f47d2e0827a0e6fb02555939b9d666526f69ef5c8dd059d6acbd01a94436;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac76c0fd64cab61da3ce3b305ade4adbb3c16d88af5b0fa5797ecc0cf90d07262fe6027fcdb0d0329;
        #1
        $finish();
    end
endmodule
