module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [31:0] src31;
    reg [30:0] src32;
    reg [29:0] src33;
    reg [28:0] src34;
    reg [27:0] src35;
    reg [26:0] src36;
    reg [25:0] src37;
    reg [24:0] src38;
    reg [23:0] src39;
    reg [22:0] src40;
    reg [21:0] src41;
    reg [20:0] src42;
    reg [19:0] src43;
    reg [18:0] src44;
    reg [17:0] src45;
    reg [16:0] src46;
    reg [15:0] src47;
    reg [14:0] src48;
    reg [13:0] src49;
    reg [12:0] src50;
    reg [11:0] src51;
    reg [10:0] src52;
    reg [9:0] src53;
    reg [8:0] src54;
    reg [7:0] src55;
    reg [6:0] src56;
    reg [5:0] src57;
    reg [4:0] src58;
    reg [3:0] src59;
    reg [2:0] src60;
    reg [1:0] src61;
    reg [0:0] src62;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [63:0] srcsum;
    wire [63:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3])<<59) + ((src60[0] + src60[1] + src60[2])<<60) + ((src61[0] + src61[1])<<61) + ((src62[0])<<62);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb372d30b9656c4cc1cb6dfff834aea18575bb379d8c6bad659bd4fd5348386f64a605b03b430672fd79204a537f04d83389777c1fdbe3564465d7b653c708e60b563bbeab099d2d56de4564890d634eae8a7ec9083be84495afca237730f944403dcef0f0923dd09c8231eb1f353d8b03bf5272cdf8d017222a53cb7ddc0176;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9e3ba24ff3da0c73e08c2f60182b816fdd0cae2cfc07b0412105fadd4897b9c1253c9489aff817ede66b897b28fd7399fd5e81b570b39e6d0ee5cd15128805d8564fa419b6d2fb6041823d39dc41c9f73e87581cf3f435118a39d4adfa77d7a7cb20191781425307da4e93250e5ade7d724b2fde5b212039093259eca42b980;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ac4d003fac6e6d2c189a6804080f2807c8d4178a9844e57bbb26bb46712562f8fefe4450d81410f7c218d3807f930332bdfa2e10af437810822b9669eb5bfedf91ad397a78b21a3278ed398f67737b582b04ef41187e594c389cfb596be882a973977a36cf73df54b55565637285005c72316f043c30c9c325543b9dd782cd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h490dd6b734eff04e5fd3370b84f7ca305a821764a091f0d5272ada8ceb90e8f9b1b788cc3659f5769d8f91b48e0639e5fd6bf62b1e5b479dc7c106f899918142253c04a9035067726c42982e9482e25a8705b4bda3ab7ad09fb85c88fb9fd157ff085a5b78b3e9a56e5b20865ee35627579b1f6255e2180851c567c67e5ab959;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb02ffd81efe4d3e9c91b584ce554f11edcea404ac39dc3349887cfe561488a69ef0a89ccb561e01f8ed695b660025d4e561e4b07e3ea3e0e6b3346bf48f8c8d86714bf6ad7deaf1662289aca4068bca90c1dd7cfad3a5f25c1318094474de6752021c5078e6e1d7588b7e7553fc4ace39dd8517452f8bac4e747c1c8da0d9c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58d0518bff0daaf1d901fccd8d906d13eb60f3a7a59aec960671481e5b72d7a539dbdc4e8383134784f124023d645e7cb3a060bd0ee46b7345aa92bb29ad1f8b5ac2ed7869a912c1e8bda457da3bc7c2bc0ab249831d523b5d7e9d5c7dad793d4c570ac4ca8196c81eafdcf0032eaf83f8c168eedf0d8529fe0266f3393434db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14f42aa94f430ada99ff714081654d7c42204c035f1f8a983a82f35088ed45269feb9cdd23c87e51932254f10ce3c128a02057b0749ca87a5ab6a171c42deaf1f1894d72abb4ea52c2367a9edda8c778d0e8923a571f60073211c1e6f9a7982116f1d22081684fa186bdfb442d563bf7a4f0426698f9468a6dcc680e56bc1f38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd51a95fc5d283301eb339674d7551922ffe0f233771df3a4fe02d72970c0d5c2c18b84b797062df56c5f2c7e569ef4229ddc44d8fc7b4833f6656c0fd888086deae3054af20f17b74a6ac236ede64294906d7ca9e58820beb71c18141a4585c8eae04d54b75250ddfec9dafcfc70fdac5e7b51a0e3f5feddc00fb9aa9f0bb38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfb10077d144a468e2c53b1b4cbe0e200f4930d76505f53c5d4aff044ee040f8db46e15ace18e095febbad21afd236abe2ec11a8ef19704e006e9ba20a73e0889eafac0332f4f032306b85f87cd2c61b9a9367c068c98ecf24f60dbecdac7cebb4c344087372a28b5b5f194423a71d0b6f4e8a5e8a15ca3a1ccf2921b987d6ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf843578c3a595d74ccdaaa6a1bff2102dc390670a2173283497624e3c1aab050f1eeb61a461dfaab230cf2ca2c89ed0986250fb80c577dcd3fd6a3089a87a7d28a10fc7557580282b6a0ba32be8b8927011641c814b7edc01e9ccfcdb6f33ef5a38d5ce23d046c523567d18bf6e365c88fcd5678cd10fc83be767f699a50ea6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54713a47f56867380417221f42348553188f0b2d901b733e4b64e7864d037ca31c773018d2c751f07c7d63a2698ca1c3e783699c98472889e1cac0a42b7fea924f1de5a9114eaad7873eb49c459968cfa6c07428e5537de21ce02abbb0d9bbaa4357d7ed93ddc3b072485198ddd570f87360edca5b5d49fb218dd293b6f69f12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h991285f4fd5c56b7ccd7fe43d4fbfd5c2ac1315b9eca3d4194548f6336b7d229726157f7d7c3238c865589ad38ed712f287a0fbc1e7361ff0531b9e9f8b6af78641821177598870899ec675b2cd851dc0903b9e80dfb9b8d479a1711fc28471529813397cfcbe327d9aba7ac648b5d2e637d5cefb1d97f33e273cd7d299c9cc3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf7b23f8e33b37120010ae30ce110a50e5885299de7a3eb1d27e4330a2469b9e9a9c08922647dfa4f0744f77e981308578dfd2f1567da85a3ddcf3791a0879e48c13460b94ce11b07cdc6a760af9394fad9cdc1ad96a09b124819a90af8d3c58203bd4b74752b1bf41b8987c65417ed9f1ec9f2daf11380d654e5f25c1591400;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c147c95654293d9361b87e26dd640e27d58e18761c160c3e32709e0fb033c0fb7a95bdce3733a873424fc5fb16d9e1af3968fa1dae8fb1590bf05076d6f7f15c5618780510df028f70183741cfa2d94faf6ceca9ec9a17c1792b6e8b7bdb0d29ed5efdcb1febf92b50e9a843dcebebb8cae8c20cbb97a573219dbc06553572a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb66b13847ef886df2137a99572551d5184e97f56748acadee16b1c29315d4da394e603ddf0c2a3a3cd562c84dd861fd2271e01d12ad0822fe69f840ad0e6a51768f47c54492ff84981bd78c865bd9f39b6a92c01ac0937cf262a0d9c736ac05a605473cf37a9a93b6334ce0c9e89a32158e44de6efef11ecb6c52c9a72f58b4c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49aefac5074235d9b8bfd67bcf48ec1a0f034ba0c2007ab9177f96fb0fd5820fc5d348df57933b9e7fdffbd39ec00c351a82d1ba72ea9a6b5fe2e47e93e7082df4d409df8a551c0a4e8bcdd0c7c6d72d57883e341158c208d74d76663456cca8499f6ab41d3a754506804157a9f5ca0c6e555421c636419d4e048e1f235ae9ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3acba12d09b823605e725db42b0f46940fdb2d7a3a5ab6007f14f6a61c6920aea8f64d7e6541bc932da1a53f569de10929cb5446738417faff1f206bf5aab82d84b8550f98306620a4aedc3663b2253f9fbaae4915e3634764eed4875194608a5dbcde7852b122d4e4048e7d3ce3a683f94adceb4f33cfdcd4d030bb736efd4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he08d8eade491ef460f49b2dc895d40965f8245ab5156652bda9c70139f2218bc55cf59814c21363c0ab1eba022a6ac54f47d591eea8aca53dcb1d6a6f13e2792cddb608e402d84e48edd5de21b2921cfed2eaa3e0a96f39ca562d1389a0d1ae350880014da344068065ba32ba0d4d86a0c7a049f54f31ca5d8e921c20baaf035;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc85aa6b71c3085032c1ba7d716ca1c458d9e972a24318d68953ef9dbba41473351c055c2d3705428e219f34bf1170a84d4f9aaadd53cecf7486ca43e13880d2862804cabc2a6e465277430805b4829d646c231a31cf20e451b4fdb082e10b31778225bd1ee3fc6f4e99c977e8859f283c060f3c16bebe9232785f002938cdc8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf650eb80c18968a067ea36c360baa00b8eabafc7f1332f5bed413f44dd5a1f3f2e767d1c41189b264a1911606b10fdd6dee692a02846e63bb7f1dfd9797f62d15e2f86b661a2eb6f94f6bb0078cd3ee1ee654f3c19d8352e67aea285fdb370ff178f74d7c10d6f4ecd69977affcbcf1fa1781bcc1ebdfd7b4f6447a660f8124f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h724215be8ef53f4ec0dbb3aa942b99601661b3fa2ed3e0859ef27e6412de9efd77caa4fffe7d1c1ca39b077172408d36960310a74641faa00393fb4a847b0ce5c1a583c090028f914a398df816442abce2b7da177972a8297f741ffe953cc9f9fb7428093506869daff886c4fc6d1ff51822fe808c384a228db8af9631a0896c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bd9b95a633896c269f1ff0d3afd7aa2b53800da8fb117465a611afc76007b76f38d711d43b14c3f0185a4016eca2da12dcee64155080aa9b6d6f3f841aefe5cf8fdcc21a1f68995160a85838741a796f96c3f8683ad8e23b64ba0501c512e8d67d084bd30e9221738532b4d748db363e67dd1f7e7c930c3b31112f47cfc9850;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h814b8fff0c88219d601cdaaaa40cb2a0560b2e8c6642c90191cca6687754559896dbbfa1fe2e16fe959c0b5808eac53325226c68fe9903a24d72d0bd28f96fbbd1b50da1b62c4db599eb65d543216201c615fe43572a64b44894096115d8de058258598cb2df3d90acdcd7039d8b509716c3ac513c391500e5ca6c8cb9f21549;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h745989013f5c230c1887e4c6d547c509955fd1f9c53daa70147dbf13525c8115adf8e08a3600b9aad30d50df8ccd528eb65c877e7f6c36d164157831718c331f688b41dcd7ede9301b1ca4a1cfd9f55348fc86b636eef9b3e62da6ad580d42f01a9544a78988bddc0c1fdb7cc1022fddca095864987147513b96e3ad80a91767;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ad06f3b65c7bcdeee38de59773e6da532f3c2d0cacaf62eb0b65de10fc951ae3baa9a12a41d183d52091b73e2dcb3dc9ef26b158654689a8e2051253aa3dbfb76916bab9e97c6a12f49b546d4692ab6c3a7c4114d926174b750629ed057efc8196988a2a9c9dac53b6b7409c4317258786dbc603bc209a1a3463eab8cb520f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcb8cd4abef4e95bcf75d6794a3e23ef709374b0569ffee390709e556f3dd656541eee5c3dabdc862d31beb67086ebac8590ae03a076eabb6714a40fead4b8140a0beb3685e9f44a58b7cdf820381e62e221de5e75d17a15f8ccc5970cf7a5e658529a511b3de08278d4293b71d32935cf7494ceca5c461ea4128c0b0bd1bc0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bf2a1ebf04276e0fca7134f6683c1f932960046d83a540e062397163495b407e00a946db8e5671f68efa8fa95e1be4346d27d45783631a044a2e06d3ffb371c967bd58c13c9fb0a433d831f4fa98ac010fc65396bb7686587d23bfe6891cb4ec53d5b8b34d84e91618b0db89096131ff2b4a4b4197f54360b11d4338bfe136e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2202c86942a50c39bf2617b6cdd434e771d3332016fab5846f7357aeeaa1bfa2deb93c7663e6bac4ca47dade12f46802dfec124681315c9f70ef551d8339667a679b85c324b55eb237ccbc952e476e6359b63d04234219113c4f1a62f2c35efc5868e4c8f799510bc88e7c7bffbd5d5ca8c79da9980d777b4814c52797e90e18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h472c996182fe3fa4c4324eb30805479fe390c2a177cde95419ed7aebb0573ecfb4c6bfbc1a2e70f7aa4e5f7c60a796a3b39a4d4ded42df17758fda5fdf197046779a1f5fd897ede2854183031f112be37b8352df04a8cd61f2a7c53c0549e1e6563e5eeea5ca453c3de34cb3765833316921128bada8859a0e84e4863007d104;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf43174140c03e05e09de86f8b18f99be894f681cbb48ea31ef1b29552113d8beb6e813a48cf4c3e52243da294479dd9ede734e5c0488de79079da25a2754ec3050a026f8d273dd9405e0ba053371efb4afbb811ab4f1bbed2010d09f27e82b9fef3a5415fad57beea39f14c2eddc251135198bc30b88a5073e2cb63b260c9041;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc12fc9011842343062ae478a3b143e11c2457223f7d4685c1fa16cb4d945987f13301f92f6a0b17062433deb2ec71d9a82bf008bab9296e8eadb457cdd3fff0bbd899a1cca07725b894b14b754eccd414697d1d7738ae126ef955539456e00dd8c2d453a631598c0b6acb52728f17c6bef1f5c2fa5cda4211761d43a77283ae2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h119dbdce9ea7e2a6b902ca194bd5f1e14a5d09ca38c1415c8851120b29887b1f55a0994428a9f6e2c229ef47fb6536785357ee305cb0b2144be0514c3b8e69a98069993708216dcfdcc98a26ba58cf6cc875aee864a8c637dee5a3bd0b95db8ce9ab7d64a6d136ba3a08bd7ddba5e14a062c6087d7143c827f863ee8c8a73cf3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46a12c325aa55a31cf33efc38118e63f2f1e10ae1234fb25e8e3ebedd2053391e8a200a07637b073c488849ce50db465a966a6ae944d85bd9a15171325d33721090cc759e729fd1b7416df4dd054fef09fcaa4a59dfdc73993b4829526dd9ec1e3e72d4fd209cf170fb64701a54b922f4b53e0da1622069818166f1c45583860;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcc8733c577cf6719076f31b1717875939ad15ba05bd81c6c93cb4baaef735a81620d519a0b9e68600b8ea7d1ab240e41c5c5268cc1673e8cbe89b2d2314f1f75fb1b123ed6210293072e121c3437f3df65ad14c24549b715403bfe9ab7db166c67216811c19ab4dc6979a582fe52cba075a9002c68b776dfa10514cc3ccdc93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h339e7dadacf7c7bbaa613e1f649cafc01e0c0a72e34d1013c460e09d8865b1d71628f11c17e905fa5a9d30f5bbd8516ec6487da82f4ce41dc32ee2eb9fa6a1f63013169f3e33eafabd945c6189d0f34d20f1588b94c4634a36b8a5e320bbcda02c4fb0cab960831a64d1cb8d533e3995b498b0b82b77e90f099fe25d6665588;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc3ecbc893abfcb64d4331b33adbe5745087e2d83f2b522a9fb03f279797546517ba2ebb86c8cb329d230f2e571238750d65b2c0a5c01abd484b8af271bf77763a0f6618517bda81490b9940634f3929b2a1cb23826e91c7a749cb8f931d602a3fe5e7c63d7723ebf02216d9d69b1c253718feb7fb59b9df4f31e15e064da007;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99859f576eebdad30c05bdde34b80e271beb395903f0f0ffe5e9894cb87e3aa56b15b48cb87156056923458b81cbacb373676fa10f87bb301668d3bd0de9aadf34855069677697ea0c018cefc7b09f037582f399ecf1d324f5c7db3bd08bacd6c05e1f2a80162c8c4d13f14bfdc5a259b5398e059c20f9c0cd42d05200491129;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcb5dc9d0e529825204d568be66932fd9d8cbac2777c1ce8d0a3dbb380bade94a80cf65f419de761aa42a4adb27890ceb918a1dcac627aabef52757452be0e64342632e84423a981c4849d1f9ec9e809babe6c0e402ac25dfb807bc9088cd7fdb1930ebabbb85fd9109b31099940e3ccbc05a74f0cb9c912d14f46b617d81654;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45007c3992140d1c6ff8dc2d42e3a8c2fbe7d5f1f9fd65841641e2b7547b35c64831965f725887e0becd70922c0af097a29f5280a84da9fd09c52475bb5c18b9c4aab20dd9771f792a4bd0b1963f12c5715ab24b581ac627dfd773fd587bda79bfa51dca7e77593e4ab19c78d3b96fd4be0dc72230a5463abf7d3d4df864f16c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4090da3f99a1eea018639964a15fb4587d118afb3b4d01171a3d566f920f24442024fb1b25966f4297c69e42f894d63cc47a413466482a664ddf7037f8127954e767e908f8cdffea03c4f3dcf8abbbf351991d95b270c4795ca2db99dab43ae1a7b159958ea3fb45784e1c7c851923e8bfa7b9ae9fe3de86ae684df96e52fc43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h782874d3ac6b8d9626789ec2ea9b0c7fc9afe10d0d5fdc109cd39f23d92ab8a8d03ad39fcc37c8094e3d2a1404d38c2c25d71b9ac4e51a551f21626097a2e858aa76dd076fa48f5a471e0648a08714a425ed56dda5d264f9628c656b35b49d974ebb9fe4173dacd166f5bf97e34f01fcba935d183c397f2aa59df03c44d2403f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd09cef63dc219f6ffe4fc8852fd35d4ad8b09ae828b6fa01b8872099ddd01f5be54b79632c1d9c902a2a9a127f1a8d5acc911a997cbd204c392c3599f4bca03a688aa37226e850f910816442222d4b9089f2206c818fc5dd767b5ef1219e5e3d8e268a96983d87031f54c07c926593ae99db6cd203489b1a45d51b95f3ad0ee6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5085d6a2b8bfb0902506367a41e388e189484748881794fd31eb389e236d93bf5b4c94b33d2af00bd5c6d2807c114d72240459ccafa21fa36fd2013971040859c074c4fe8d1aee1691ed8b95cc7d66c5ea1b16e5966d448142baa535756d28b55fbd1063072781a1285b4819900a6f223ea72c59c9c32c96eabe8ec2b73e1d2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h875ae57a7113f2ecc6dde7e7e962d39a96c6ce2965ca2049b965ef1ed58c222bce2ac6b127dbe8fab841d1fadc9e896db24a7abdd5e9081bdbfcddc1a5ed0d532d6f8c68e3c0095635e0c912c3cb63b5b73266d87e756be75170f3a17732471b15727a6e53a64c4f973bf70251bd8087d39fc48429fb94929cc7000b8b97a49b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e4c9f66fdfe3cdddf1043c3c89b30dfcca6ac3fc2fc002c1795ed15ec00d9337ea7647ca72e8126a889244881132eb695f3822986bcfb3d8bde9807347d49a329211300d16f1659f071451d5f43175773458e6cbb3bc81f925d0f8b2d21d3ad4d32af29b9c13bc2f6ff483c544cb233ef013d48330b7e83dea3f58f5dad26c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83d7bfda727c053b19bcf9394dc86382b3fc16833a66369df982f964c39944e75a677f78d703a2831f5903dbf45186473fce3e4faa72c34e4d09b83cd2a03bb875ac56a12fb6eb27be8fda799f739f5c83c6853a58a1d4a35e121d2e8e8495843c179956a83ca249405b68b9dfd98b01b4ce7859c9fee71b15ae6ba5bc640532;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bae04e30ac201602d535b4342fdce7fdb2d07c25ef413aeea7cdd105721efad6fd2d9b5f29ea1d70f8c2ecc1bfc908278a6fca72814d2cc8265d7ad4735b0604c447d544f70437624ef45a0d687fc35d30c583252b26713365179c183109e88fdda073b5837533ddc475158e15338084ed28a83e11bd0cf046e5c59e86e56e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b4b791d5c257f7fc20b673432224a2620e05181a1a5e446987294a7f95224ee41094f504695ba9d8560dcdec51d3918af41fabe3289bd5eeb5b25f45ce5d89df0918bb214ad24b6ad8ef6c2c06faab9b10e7c497bff6a06c07b08401ee91894fd94b81db3dd2a6cbe8682bff4e48ca820f0a0f277b41bb8f8decdb1f207e367;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h716d7e8f6cbbfd4b162c4eaa00b5660ab3190477e97312a5f5238dabd31f8a63780dbc05f57bb892e4647bd28a6d207ac8c7b7f37260fb6aae8364be506662393747c802512bc6546bf20a59fc7d9c83b0229f7c5c1d9fd2f10ea599349ac0474e684fc8b45b85c6f6aac477cea429fc10e63edbc136ca58e20ec782ec2147e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf4e301626a1ed10d58d48977051f7845c0b12ae846347681f4bf8a65e853237d50595540cd64fdcc6626192df0b3ccb57a096d2481706add8234400fe2bfec42c68a2509fb1c0c77f7fdd02433c0a22372c47b494b1a797aa950133ba676bb4e5dd3bc2679e10e75c2dfb51410a570b731e3db39e0f02e9740e622812d242b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43d62b9d5d3cde3cb31326ca13b43ce1a6174842b6db8d8fe1176483f4221e5bb676ca6427abce1e6c3f1ce50733317a0fd75da6a1c10770f9824cd98e0be726a8712786f7b991eced303a7d0a6556cd81c28a6ccdbdc0cfe5dbea37e94b37efc68f77466d802bda3a52b09d42a651867fc0914a6c8d2d5a03440165d555af83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b232178f664dce91f4f572ba5d5545a6fd706d737e621b2d23c275b91073aec2b5aca9e1a7affe4752a20d0003d9eb658d422f03bc07760a720ed312016928ac9ba0702dcf8975663369d8a219c10b1a4b9a7fec17c2837d82c3a86ef281547f4aefdd2720fd20a17ca94f1bbcf7838c775beeb424a95c4855bf681205aacb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffba7dfc5dc22ce189d8b4c95afa87876c06a376f7c9dd400b564c92bc40cc04711a67d6c744113a9cd27cb1f50a5ef1f6c232c4f9d09aacf406078df4275acf3bb7b8fe13b9b1e037a6fa11315583e59f23ed2ad6882e7c8a8ca54d1dfa214bd7093531d4a92c2ac42a3824dde4093c3cc37e8f497172ded87d7e7c364d460f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54f1c36c88a32e4f9d89268be187a69905e7ab0999a352aa4a8e1d1798a83da59c7b5675a183724db69917c103f37d17e6b4c493d028669966a333b5d9f0d0ec6e3f56959845ee6c3b4e96b1e4b477be63f1ccf3f26830202722616a2e8128fa054196069e63b8aea8f7d8d8f24c6a41710912441027487430734461ab2a4239;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d15c55d1f7d10ef0ae7134a364c94c71425e6cd5c608de7227a1695b6fa6d846f3e369ca69f8877ce18d0f2d6e783231ee3c7ef1a604bb428e5e03eba3bee65d791fc90c9ddc4ef01c3d03819c9d6828b6776bc66a5283b5da972140c01a3819b8e00d6e542b25edcdbe78d650f0dbba90fcd52e679987d6b5502af14c9601c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85eb0940ddcad13161cbca18848b020b952835d5d658d9b332e2a6516fd85565c7bb0d946c89959fc5a1c357d309c9f642777b76668580d682d3d77e6e5fee0da7ff2222542c8e8f944cd7e580963265455cf4922ca2ec741834f8d620a8709365e8122cc28f576ee24e8fd489f554caa1df3c4bf563881e55525320f8e77e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hded55a30666a297ffbddd65da2fa5cf69be95fd77b6b954aff760396717152d5ac8404a4d1077f08cc3b86d79d920ce4e9391914e5ddbd7e61e58b03b956613705ffc652e0b2f3da239e08bfa1850b9b45c7361f5c79b43feac967f6d4c39f93031203184211e93169af127dc3e874677868c8aae3fe555521a680564a193fd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he57c0c7c3ecefef068fc43070f48dc24f1344865969c62f0774c986c6fc045feef602c3b3b94f9c180d1a6e81ef4143af3c7298792526438417a3a01b5e3543aea3332650e27412b15e4e15554c0eb2cfc7005998f191b4f293b96415fb531e8d3408d999fb142cbd2605f9149f5b9afe2158b36d8761b5f2873eaf6c43149fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3055ce982a40b09d950015d66e9892078b01bd9061a45899d98cd8b76c45d43df4e856b1dc99bb7f4f01cca513c7c9c856b93ff7daff157fc111b3d0e2483ad1e6e52f31265ca8211d66aea5e47bb1b483049fa8157111adff264a7c9992bb476f39de351328d00f8993d4d79d458bcdc6b70118a4b21ea81db7b671a2b802f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8acd0f06b0e9dcaa3c8461de8fcee45e04fbf4f9bf7283714b01b28e2f593c28e149d85030952054f6098326218bf36f3ee8b7205c1c3bdce5fe1d774802d09d42d660a3a9788c5d4fa5ab2574e1005f7b8f2fe56349d50f19099148d5fd0024d8cfa02e01727d15384aec89760c6ebef6504724b4f751cbf868c632baf53014;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30f8e5a193d549f185ada769677f5f0db673b86433d3a4d34881785ea36c37e78a8d2b4ccd6f96109c3fcae568b67be1f25f66b6793c91d55e62e01522f779938bedf4c3ddfbc21cf3ef2f5ded94b183e0234863c6984d8a86cfc3e7ab0c05775920610c862313934b44a41e413b47be65734fccfd58961c71dbfc88cdf7e668;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h272b467c51a8e2352433104cb1a3c48bc65944cafd60bb47155d18bd1c4291b43eba45271037ad6f77fc601be7284fe54c04df2b899ea5ade2d26ad9a5ce68058ba0500829af510d1abb172086d292941bf96edf00dd7ffc6802f0738960ae821dffd00f14644c2d9d35945cd26363b635cef242680d4c73db817c4cd805026c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda05103a550618c38f8db568e14ddec3b5d46579e52d502640eb6b46be3b7f1aef1d23119acb71fb4881edc17bfbb1b43baf78a68a5ab423f1e1e52309eb54e3efdf42175a29f4ef0455ae2998337e446b47f77c400740f02056daf8e3ae65804594ebfa0d4ad81ca941982a00ab94d3f2faa3dbb3d8cc8a95e6b531459eaed1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0c1aa2910ea3f6467a3ae4e71b914c5fe9e424503a686c328797a83049d711407bd2a76265958255ef4a57763ff0a7eb2f866e885ce266ee6e0fbd79d0fe2147cbc92be9ef0ea5560542b0fc2073fc92587c138f445488f079c176d0eb8053398ab71221e5bae513f73216408d0d9d8a01e1dd28636871e96d19cd162f27f58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5552b22bac874f68da2575ac7d6000b5dac432128b87d0861c3678ea30cc8585961b3a584cc58e7e4f4985bb327e1fd30dcb4700f71fe7c470e42074e90cc07d8d71ed2e502028158925082950af2ef5c4e835b2869ab5fccb6939984648f4d067b656b09b24893512a1f80f98077087cdd50690a216007fe3d6d7553e398f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13a239057cf8ea6c8a06b895b0a5b980806596c215ac3b52d042c2838a145842e5721c5de4956444ec983a10df5617f828aea2d59429b40d453d9fa530dd7ea679e0c0983aec854a3bd9efe50fdadd2ec25e16c76ce034973574b2cd2d97a6b5fca6dba56ea5f0f29676baf51225bfc045fc793cb0ffbf07450ccbfed64575bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1501b46f1166cdc59076b059ed355a09dc1a877e9f60a37554477a031ae4fd6e28c3beeaf700e4427b8904a5063de8f2ea40d17c621bcd6346eb078392f4d009c04a9c12afae017f5b2664e82ff399e300eabaefa56ae88463117f6fc8b4cba5971e26593198866c1be70ca2fab4fd1d58f10a56268d227f840e3ac02a92cea1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h206fd2cbf9b73b45f0e8cbb21948fdf76d288e50048806ea73da892c1c888a4bb9f2c5ab89bf9939ea7f6fd9cccaa6ac6006c62605af703161027da1d5d68970c18aeec40e3697ca465e9fc93a133c4f3af5f046b0e369efd490926fcacdb06d49aad5bfb9a1e92a484bd595f7a3511037680c80d77cf5c0ffc95537bbc14ab0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf98471171a051d0c5fe9e0aacfd67c47e4db077c5236b7ff0eb907a2c9d7462b7e8dafa1295c2216d20275f5c6a93fae6eb1e953c49bfe854ae8c3425ab513d55b9c8a415c1dc3bea6e4f4942c571c0021e8c247f2b9da44a33fca7eb236a703121c0a7689bcba2a6aa4f8bf2be1f66c83af89cb04d0e76922dc3bef42f6e61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70c187fd5cf8d102cbd9b8c9c97557727cbb6b08804f7236d8c2229e87aad726bd264917602cec0f46bfb40756bfdbb3fc261c8c2037434baf897cea25a35916c86d882e95f1d18a89fb841cf3b30f6e0dfb62e45f6e7082a2cec04af35d9174a95da21d0d50eb5c18d849459c30ee536376858506b445486a8f91e401b33d24;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5086694ff600525732ca4fa358dcea93f030b9f58798a9645db6f6bd008579458410c865fbf7d64aa40266ec2c126d3a824170cda77aab9d369561e80d29d687de0d9a268fde9da70cb6e6d270ee27b822d871ab8e2fbefea8cdf9af17b4f8b90d2975611a9ac06e7741ff2d322d59325c2a0669d20817363df5bc2948684f3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbbaf2d4d4e192023c9fe4ad7d510a1cfa405425531e011331d467c760d486aed421fb1aca5ae92d34a6a39cac3d36a7ec88aa302f5c782ddb9edaf26a5b6f2d81fd661767e41bf8d00be576b168bce0d263705a616a410f2be795be964795b490ec47ed2cd97946cef5df13501603e06dc4f6a1ed3c2ae86089b2bd032842ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d579208b9ce451066ab3cffa9390b9b8444cace1846f4bb315e385eb71b418a9d8d048578053153795af67afc31f0fb3b48ed7b99f83f4d85a2fa5b26af089ae13cb671cc6f610ccb3db8e1d2ebace17edff344b8a4cd169858481bd6827b9825b3a22bb72b8a42ecd5ad1d257cf15b532bb9bd49f3bdba153f5d26450d7f0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d1fd7a883698544824335cdb4d859f5ebea8056b086fa3fc2f29620c969475900eb9539ecee06c3afa8a496a225359e5490126902f39f401e62a9340e2040f6a90cb6b0fcc169e6e846b378a206d8a46ad61346c152c865a85563c9879b844e3c7fcaa58e3f4ec4ebdc9d259b52d1c8e8f59423c2b688b37b93104400c914a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66943a77a80c6e3ca68213aea2f8b603aa2b08f0445a1beed983dc5c359c855e4fc28a2b4ac40700fea63217a121496305e8d4107b51610068b036a597bc14a7bbe8d2c4b1b433ba82d102aa7d4e4c0204ab3a3b2fc24947019f6e58fe3eee146bf3b7b201b116001074bba9c5d7f9da698f06673511c785715144f2df19841d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h397874183cbc173d98cda6e5a4e47f40c76add5ea5771ca17f3076fde7b473c9757e81b15a5ff14a6590e3c7182a83c4f9340c648e5c34b8148d9bfe8f1788cb39100e7454971beada1d12091f0f2217410315f9ade5e4c4b041cb4b258b593b6cf83a6ccc7116b041cc9a25324077829d2f69b496e16ac835f2d52f484e9c86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c7bc347532b44265bb87857eb2db91198687f2c8dc32ab3d50e5adfa84134b5957b782e47df60d11be9c52a07d9f464a9539b6f71ed36daba17d1ae3e6db1c870fff4d1bfbf5176de16e2787dca21e63604142f72f07f88b3514dc1f631059bb51bc4986741193299a08c81a14d5e40c9dab6eef25aca3a12803da3e33f450;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54035ee2bbecc6811b98b91923f1d14e83cf4d2a48e1a8fe9a3834e07f056fecf6660be990f2e4c6fe35bb3cb7c2f04de11fe31ee454a2a26a7e69906b6b582193f32166b7b2f4ed66bdec22484fbf306bfda1f9ee64bf42ca682376e2990b6125f52fa804cae04b998d11a6ce3ae3d5cebdff82c91edac55bd4618ee7110bda;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b63ce701da779dba15e52e8fe1c0d4ffd697ecb49b6b3f11a5aa6fc3c291c0738f34992e59b9f4c3fe9fb6919dda10bdaac5cc1cae0dea68c9d4424338d6b6258cb475d76f866fdd37755f74b34c53a795d12ccabba0079de7b2408a4816ccfec6702487fd879dd89fdfd497c8eab5568541490784acecb04370ac96c47c178;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2833e59f4604f6b7d14830bf8670f93b7fac640f499d1e5ab47f1dbf2f58807c1ef1ec1fbddc6b853173b85df2d5326d4eb0b4a07700235c442a3876c31d0fffb5aad7892458ce9a7fe13bf3f96a5a271fc54ace7c9c244b68b9278928fcbbb6e79be5e0133c09ed41fa0bf85beceb9c77f5106c355a784dd7b7f421a5c8449;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94f4a735af81274e1d8517fdfea2e0d5526ab5687faba212cd53704758d363bc677504ce8ad978f5025411049b3590ce6e2ecc93a6ce646dd2833dd48e9fc9e44da04ddc0fa362e26ea35e593db338f50b1d517e2cca80c78aca97848fab40caec0e382af0e1e7667a566a95ce9fe881e77c6c2d785fd207ec7918dcb6b00ba5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h597bd16f54ff7c414167edfef72df5e203a0d6765470e30bdd5358dfbea5902889a8b52a347f7893af9e1126377579b90c19ae0aa88f842cf4c17d3b4fb924160d2e8c8fc211a66cff727697f0e34fdaf3a9c1431a329b5f6e96a20f2d400c63c507ca4d9fb9be2c2abd5d7939c2c2d4ed5eb7c45783cea7f5e1cdea966c0b6d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf47477c11581240f25b55f762d8a1b87acd34368da5af9d0f35a584085cb82d9a0b6dd517d90ce49f552c9c0d770def55cf52d0999faba0197f0ac4e1d0ffc7c49876c1f6fe446938d9de5dfaa1144aa433dc1ece121254a07dddcfc7cbbc0208f0200fff7bbe268c1694c0cb1028e67c118667c40bfe1f59c4d1c99ed0d45fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcd55537b13bd879311b55a364dfd084bdfccb37ea07c0a0bee2656066d247d28e19432d704ab91ff0cebc56cae13a45a87cce008c7b7bc22392387346bf02fa63c880c79c85516618ff02eda7bc65c5b00dd86e611d2b301899553436c4c3a3b3cc24b5e414a7f28f19e606274cccada33c8fcfb7565adc8742d56c07637c05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54a9f9d7f07867bd41c017ae4be7343ac3286e6c21e41c51f31b55dd87b42392e843fb4ee6c137fb733dd811aeac7d2957b53547e3c4008aa062385b6f8fd9d201581bd1debbc6fcc7ab0734de1c0c99678ccfffee4be90943685563d3f2025487419de337e5c32ff81cf000706e70f739fc86dd3078ac426b632b07b4bb81b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3878634ee020bcbb9a0d17df131f9c3d4ea583e40ca03729900dd20a219af7ea187eda20746084e882ec43004bf96e6c1333406ce275aeb1e3157a0ba139202150bd01ea10b91f48c3010c787d6ec2c995fdef594b75f124f28cfdd37149fdc517093d6c9e26521d4a03bbc5415c08fe74d779736f2493086e4b69cb848b2411;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d5738b12a173c4cee9afdb55185503939e2bcd4fdeb5497769df764c6a8525024624e81b3f44ee9deb130a14ddf083860b4d4998131317fd75548803b57bfc03b427c63965462b02feabf17b6c156c67ae6517ee5fbd0a1692e45d8cfab9aa0dac3b76450aca1fcf16a19108c14f6d4e39a902d067b30ee2d05a337a009155d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaf29fa7d3e3480f93c0c6c0e051d9bec42ecacc1dcd8efe05018b776b76cc7d16e73432c038289eb2bd8d861b727229d1fb1bbcdf8ba60cc6a0469e1e0832b4d84f3825718efe86baf7e54ae9bd0da703619d0705ad8a4de273cc84a5891a128f77851cbaf246effdd7e608c76ea318b32015348bf014c149ae766afba707b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h411a4f60cefa6771da313d3af64e1eb8fd6c3702c2d1b55c8d44da5ccc3c69225d261af2368e0fbde04f8110c25acd3340f9f7370d650a7c0ee45b827b8cf7e0856b6bea96d353825cb874c825007e1279aeb6dbe5f7a20303527b408d7851e84168ec6542035b726849ea9b5ecb23279eb5411938bf81148b70a474708709b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ca25499c71f731c0ab63da93e97fe9270af9b5090f548b6b77725fde3aaaa447088b0e053bbda35974d5219871473f27b0ea2e2d739f40dfea654e0b2c804e26be5985f167a595a7479d2a4e503b3340c584bb0b070ce6d2ab2dfe40d433116eb399dd538483f36dbe59fdec2283d23dc987fc1a2293e3ce89634f5652a895;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5a68abdbb2cc2ff51e0bcbf4ef89559292069c13dfe69ae7219cb41e19be9f67623a8b57fd80cda5550d25f4fc8f29ec8edefd6a0e1f6eeeb2f6568be2a7a84ab73118ef5d3156f275754ce394f7222b66529d7f64ddc733ea91c9782a308172ea6eaf9e53589654f64e9d4328a66e1573ca7d43410e978ce8c0fd3b2b3f051;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73145529a4e07d49d67a7e70322e7d8b4f0bc33c87529c244251ac3158faf9418766b206a48cf2009b1728cd17f31518b1d23a6fd010eddc5db57607e666b24796418056d6d1ca5631ccd48dd3f3ef4a7d67630b545c451cb15cce9dad919d4790f7ef50efbf6ff10dcb4cb32f8c160ca2cfbd43f48dcab028e5f1926b3eb441;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f3df7f784e758d1cc40285e02af26653dd6fdddee74714c9caf3fff57cdeab9f44b99dc263dd621fc483ce5a60b206ab349ea2a98e90e8e8497c710c7a36e40333ef39cb6ba55ec1169cfaa5dd36d14d46a52f8bea16a688b8cac75f3034843b165e22acd781891224a3230d68c219d0916cbb5c63c7f81e3c4763764b1b886;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cb7f33ebb18fd1d21d36cdc0c96c596899d59b2dd0f7e8e91f340e2d49983a9eee700332e2ae99dd4857524ea7058c1fe91f0ef5d9445de49e08023fba4356dbcc3e264f4d3c5977eb48fa16eb14087f6431055e2f12db9510bc84ea4393856ef94e2968563ce83e76ae0ea928f82fa4af44d2ca19786c507eccf15a6728277;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39a3e80a449ff67e1d6d42ba6c367c5451b7659d4d98079e285a2d9e541080a84939ace86a6af77e9b5cbbf83eeaf7a53ab268a2c4919f35960359f79951104d67b28c59796a83a3041aee67367bf568d378263bc698d0bfbbc7a24407c8f3a16a35dbfe590be00927d98641cc087edef4a69eb74c98cf4842c25965668b2398;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaab86e0a50bed4ee63fc18406f934f4279373b32343d7858b4cfbbdc0f8f7125e63b730cd1c620145d29d3922557fde5874370748fc285fefc10277f658045cc58f6c224c43fbd8688765e84678278a2b8b4ff43afabb8edb2f784aebc4017c38e70448567ee4bb5da24be21639e2c1130b7a45b4a4761cb821f6a5c0921363;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1ae43220adcc21dfa4976ba00732390231881df71a964b913cdeb2abdd266680e088f80017ed866f2287444207298bf81ceec2b75da9dbbbcfe4bbab3cda1fe3c2d563be2ad6265aee5741711bf47aa2c4f238d2b49b20850d5788dede3ccbe3d600e93519d885c21c40dffa504d560758f93c3e7417379c5895b7438361657;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b9fec187eb46f4983355331b36b711ad8b55168d8455e842979246fa85390649dcd21cfcff4c4de900d6d7ce7e8cd5aae0727d94a139a43464d8c0fc3d9e8576c9312ba4acc952cbc846f95217adf6e1b834702fd56cda65765091788a7dcc01ef637c7e51dedad87bed346af1c9010212f27414dbb4cbb85920c6d1bb300d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc9b0a4217a16ef86bcf829892b2390ddf1de0ef8bbbb2a5615a0993213f9b805853d50fe3a58b6288d053e80c16f7e5d52abdea6b8c59cfa6cca655bc9d1a185878e5ef86853d8e811e7088febf8a085835f81125b670574fe902378c1896b67ab603a60382c49317863af51f3a2050ccc04e7cb73ea629c97f921bcb1a6a7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1d6832168352abdd3f913919e7495109bfce784c7d226571e3b71e286b97a9929c1850de9c249042f5718667ae4a1daa68df76e624e0e9bb0e441eff220073c2c3dc16c0c5fd8f8978b6b4c7ffd7b725e880a47f3be386dfe056afdc7937ffc1210d163eca6cb9d4725475b3281821bd365fa7cd1a8a3c7c633c575506355d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30228db175b0382b86f936e55adef81b636e7815a17461c5e74fcd137579138688509397775ae592481aae170701c8fcdfa49e099a36100d7bf55a9726296ca12700dc039c178aea1d9281d32846e083b74dc82f04fe1a1c1f89936d04647faed239724729874a141b82bd7da6252d2731ba4ad880649b9bd62669170b72654e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf183baa56491d8bb910fa4089a51dbd48026cbe78e4f6e3877c478dd75d9fbf041e38f5f29a2935a33d53eeeea4e4cd02bbc67a3261b4601f92f0bd4511170cd2bf43392f62be478957f2f4709f09a64f07b18146deb84888c5da93466bf80ca85bc08a8ce3ca59dcbe713b58f2444995e5ff7ddf202d642786a4e8f4ef4953c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9108fbde5abd8c24dc5061e261d9ce4831a77935a8472f351afa7c34be7ff796f1879963fd40d2f1d10730dcb1c96ddcd96856cbff4c379aa177d878a2d03c025e1d78f9fe9cc7af5091b63865f629b8ab11a721e78166ce6786fd8b0916801fd38713d658532ba9b2924005162b76a42386e5d175e6d431b2671879d1025a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6213080ecb150a18c72d16f62f2908557e867368fc04c286b100fe3c47e45dec7b7eaa258a0a7abec4d14922ced7a02ee81e9e09301155bfb7fc313a5647815cc2ec6b865d64b209817a3936be2cc6448df3c9e6451ebf189796334dd2a5b23932cde38fec2868125674436a94fb0e54f0c42d8361f2276a33cf29e5d660fb9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1308319118ed8368917f214373ccced1baed2b280a3dfdd215df5df996932f23eaff32cf7ca277f8a3f92b268d6cf95363f7e882836affde728d0e3ab30398faf7faab33c392ab086fd7bf85b28d2a27a9a0bde14f2a42d468befc88d58c16c2b4f85983dbf8d4148aa3f8324b26e76bdf74dabf98bf92872947593100ad7280;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87ce16636e092e20ddc03bce62fa81fa7b0a8497f484fb60ac0ce09d967dd45fe168d07f67e51fc28d9ae2918aabd3adacf162eba885ab4608df1c0974631f41734d3477ac4a18a2637681b447e0cdff7d451472d02388cab0f490676fe03a29965527621bb8de1c0a33e44a5ea53598e84310e85396b04b73b9a9b6e0c76bb1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he51afde1dbc0493944ad5f1132184af72f56c6adb55d9a3b3f78a8490f7a1ab576069c5aaa5df075ac1c7569db1211a124523ae8ea4cb31c216327e23845ad735974b1a21881b861a6d5769170d3d5bdf2309059afeb1c27dca7a71077d7352feef2b2ed4c5e970f205f6f5d1ed37458629ccebc1a7a75cc5136e8568d090ff8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3d5f2f4c6ac1be9fceb03fe3a4d15c67269fb55ef43e973d1977206a330008b05806460f76b983d58859beec9593354f6b0a41f330329b81199a56d34f8095af709e4739b8d96ef9d67220144224fe8bf9d9fa5cbeabc122383dd852cc4d1273dbcf6d6476b1dd567369e563c4c30298b0f64f33dd2c6d8e77c7b5a728be2f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h657667b6317cc01400e050d30238b14774c6715af9a86c94db70a0039669ec992ebbc4ef62900b9ebb39f15ab17c1792fbba6de51fb3d8a522ff73c27ab6e690f3f44bf3a9be570194f7a48ea8afafc5ea7552f05638fb87d8adc3446036928870c8b6406a136405f969fa7154f438f80263e22a9fcf32b068a92abd2dcf9b83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbe0f0be143a9cd7e24bd9cc90264f1f7cac0d5faa8aa97ec0790aa7e672e44fcbada5751d9ca45ff50d2dc532ee952420b0b37e1dd875ad44c423fee2223fd9e6aa6531aadb2cd8fdad7b4c5276b5e17353b522350c4e7e5cb31efea0b8e1e3c76c2db0f3dc8a8c973f5c9cf19408e420a88a2cf385abc35c51cfb96a29e705;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27cc37e1d88c45932814fbdf4dfe22c601a8102a3080beceb09d4cd82f27597d360571cbfc5e6b94efc5f7cf709ed20d3a35bd01b5db477228e8f95681fd24189c93378efb525db8ffd8b7cdc99d1b5cffa56bf4ceee63dc726c887df0b6bde71a834d5d785a9d48e8cc68e8d398bde3e4a4b09c78924c7f7638d5794b2944c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28d036faca7934d13e704c228d8775f73864d6e371f8c83af8f82c1752cf189dbd3bb69994948050aca9750ec194ae3f6c3da9b9cc0aa5d79212eb2f1f0cc8d1b65c38c860b6e8fda21ff149fbfb0c83ab0d84e3a0b26ecbb1ae06550d5f97e4227c0886d24c03d75949f06a506683cf26b60e3f48efb024fb44232edb5eca06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38e9abd11ca827f4580815303aeeee02b8261f9a8a5ee133c4a614baf43f6b5d8a2152a6a020f55e3a2e989b40f27088678f92aa5b6d2800acb7969dce34132c72115d10113a7eed08be56842e49b740d7e5e1be46becfaee40da446eedd1a34ef43ad7ac3c470b8dbbf8cc8976c2ef1a5265b84c78e561699a41ab74d587cda;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d37e5ef3217c875847ba97abc8e793f159458244af8a89de1605419dccb01580059ed01215025fdaaf5537e6268b1c46a96a07c2abd83d2bdbcf7fdbb5dfcf1a1972a6629277cd31bcff369e4f92b5dc578362daed253d21d9dbe9c9525e08c8bc0aa235592783794ea95d3e88e7398ea85855f5bf1fcec5284e7b60a785ca7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd8794c954b49d912cd666209c9e23af684e22a13cc1d21e755e87bd38e85e8f7b2388bd32713227716eaa5eefda85a356d161857a8ea2f007d6da0b0743a5ab30bad48b7d5ddc3ab8576258d04e584751802ef21aa805c917f4471d53fdfa423d4a5e0171aaea9a59be27c57efba7f8c54ffb533f98149abc0ed4984312ef45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1de8ea62b872c2424b80f832db711ca15a76db8a5b54518967ec746348924c9cd2a2b25505de7ae2bb0ac9658e0244e2aca651def75c55635066e710dbfdd307981c00d2dfc62168b7dbe0d319a98512cca39e6530bcc8cb0eefaf71b6e051e509de5d3bdfe418dbf935d1880b2a5644e4caf85815b602772d3e7173a2df26ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45ec06a271f041e09a38796ff6824d099cf5acadfd6c93d2c7b46742dc86d9fc0c04531d12092f0d306a7f5cb19578f166f1a85fad103662eaa7d6f4b82c8b1d9eb534b2e13ca7453c7d99c914928c3344aa76bee2c4b93796266786d531fb869380ceb7b20ad2ff9de0c4bae75fa4bacd16878e8b40ccb72ee4ccf8f96fbf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h878b4873de901aa230614278846358cf5ae986ff8aab79c83448f7b0bd5c3bb2f98c7c320e6f4309c48137858a72ecd7d77d7b79c6967de43c608e7927bca95d6bbd419767de142307fd1bed46e56782dd220a4541503e745d213329735870851c71c66d261dc1740f12478abd28701f3ec33e456d5a39c99ffdc45fe6698957;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41f5117e1da40839c0fbce02e9804389910f726c26305757a431dbd050ecefcb72b6f9b2c73b4679d1679ffc4b433a8c17fbd5eecfbc8f9df1b612020874e4d557f2d634245ef983c574ad7302d392957405e1299bf65ca4ae0f7a67233b3ce422dead1bc07bcc96226a0922356d4989cd7650302dded2dc12cf8641030a94c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c06aca547c6e63a54189231cb17f1ab77f29b1aad561508db7fda2158357da5b48c1c042c6a9455f7acd5bc0a8bc5ed2ed433f10e54bb1eecd1164191b13f1828b4e72f0e01279985a4de20b0ce7a0d60ccd148d268922a1c721bf3a78a336eb29b2e4186c1536d58760843e849e2b82a7ac607a6f6d7204d2b0fe42f855c1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha58319155abd728e81a82e8bf2f28313888d2ae650f5c0f2020a251568f7e13111b4e2921c74c08b80ce6b79416733574f9885e99d81516813a3499eed829b40097426d9357ba7382ea6671dec4ee574e3585a2252fe3f2f31382e64a31905bf0f2f3a4ad15975715b1fc6fdc945e6c2435f7ba9d5d8aaa9f693734ff7795520;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h233630608d50953f1b21ac6dba7dc1c1189fdd83873323edc1876e824a7b552eed33fb864f93797c8e279702ccd7f6fafad8711215e6e07f5d499766e15950296b3781b1bcb10016e69ea62576e22d918eacdf05da7cda5f3d069ccb21017bfa74524e8540cb67ba08879e6e5d4c326df7dfc76cfa1764ac8af41bc0798a3646;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h513710e683662c21cb0cfb9ce5c669bd6ff03ac50e61394d83554fa1cb75b9c4336a683d7abd3150adcfc39c801fdc6650be969e8e77302cbf849b8a7bff6b51f6d59c6df9abf3a306f1a408f5953f70c8c00ed6228888d5f90f9620eff7b1d1de53361aeec4511ebc3610fd08872bbcd8cb9da8dbb6b39463a3c37d0481baa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8e64a76f054df6b27dc01eb944e00bb15f33558b23c715161f5be4e0f46970dd9526afd83cd7664fbc4a4f19ceb30f746dc8a30c4c6ba53658b04e77267373f2fdf1d5afcab2186ed18a659aa61435fded1e60a66306f2bc85d2e35815ad3278a40410f95e7e011c35eba2147311c2fe604d8be7d8acf30088d1e69e973a4d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8fbf6b545c3e319daac6952606f60e5900e3c75b3d5c0953f39a41327bee72b73af0ac4e5e3b36c8c290fcd631764ce327e1b8d04d60e2925c48518f789f2501d33d875ccd49c3b5b24614cbf98a066176f8439443c9ed2d02632553313b25ae3a7304f21d39b724bd55f2f8bcaad3bc422a11a1c2af2c3487deb36d500b53;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f54dae3e15d6d69cde9cc9448faab054b98525767de3b1f47a07952031ecfdb2264d04b117c50cb1bf57bffa50b694be175bcd98cb36d64ce471257b275021d6ddfcdd71c8c2b934f8588f738d80dd091c4dbe9230f11a47b640219a80b7d1112b24d990ca68101da9ed57d4a2df1f641b16c868cc7f94d94a01715752c5a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43e392e6e8c2e4eefa15811f4e2eb0a503145af0bdd8d9c990d4b981fd79c3a909e4f5c85c94fab2d7071deadbcc07763fab3e1080b29abbf574e15ee1e79a55e87246572fbbfaee38f3dd9581de55e842b79edaa5c475ffacfab44b0c086e699a3ed9458e44d0ebfaf32ac398a03b17ed9a816095f2297d0fa40a56e043234b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab26d79bc4e1457dd0afd2920f4dc0fc7978c01d3ce8c74447d2eb35530ef1e271498a0c967f08df28f545ee65b9f90737cbe10287fb5d58120dd2571b58dd0a526aa0f7f3f5213d68e8a7dda35535a0da0a009db4d6c1288a02ede819827d0aabb1ae659453aa74c367356ac2093c9c42f816114fd20327cd13946f73745091;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72bddb876088b31f350f6ed4c79050383f8255b33ff8dab46f44013cfd7c78e72820857c629ead46d31ca4cc714b236ab8ba57565e0fd40ce773dafb120a006ce24eecc018250e7d6fbc499a92389d86176cdb60ae4616640042648ca9dc615980e10d12b36bbf7febd04526904727be6f9edbde1adf7ae09549632020458d71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a3fc555f6fe629c92f66900558ed66571445e107f1aa2ed5619a347b26f2d9a2dd0d59346469b374272efd02ae83995082af01775fb61a50ed4f11bbfe978110973a83d9d2f7b96f76af98aad9bd5fc8cd91a8a633ae79afb6ec233a33f6d048ea2fa082467c6bebe3e4cf6897b4f21aa3c6d8497890d5c314be7ca32d49bdc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h416b17f93e45b8390be7543c301c93b0860fc368ad8da3e542605b4599bb1aae597fa78c49d27718b437d7e41fc69ae80f140a24b990060da5690b2e006e3d06e4586885112d1272aa2eeb7f31ad2cb960d060c947450d31a198fea830adfc707cbdbaa5de3ac37f0baedaf6a2883e1de775e33383e122bac1aa68fc6fd9da5b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he62d16dfd0002299b2fa7a3a4f34fe1c8f40bb68f4e9cc368e16106f30843c4c4975f1c3962a44b470e093b8f60cb2a55b5b0a3fdaf1807a33cf9ae163c2c670bd420ae6cba24ae92b062b4fe3131e30ade63fe852b67ec28cdf02b4c13b748e37335b777b60c636801fe469c3bb8f7841f214c7b095d60f91acb1ca62154d9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5196acd7af005e8a498114d1b33f683ec9e729f778154598f2f53da4db51b2b4ff5135f2815df4ea6cf90a70353a21fa0c282ba2ad94bf472384b84f2801f7c46df35166439bca0cdba3f0a9c857835c90642fc61bb44f9550c9fe74c5e71eb8ec7a1863dee203a65035cd2b57642c20c322f0ce3ce99f19d07bfbf15c96e7ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha546109c90b4e98c82e45c600deb81e03633ff838759f831fc3104a3026f1971703f6968ffc367f5dc2389b59751f908a3a40cfdaa44adc2fa7cbdd1c441b1b92187e7de80269dffe9f78de95af38c3e9cedf35f51945fab791e734beda748fadd64e8a6861c4c353c62b3673b0424fcabe8373c93caaf8f8ca86ebe7b4ab301;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb460da7b32bbf012e2bdbd7d6264c15b9dcf3927ea150b02ab3c44202d5df38cbcef4580f4c318d0aa070ae9e5d7334663a862985be8d2b8db3a2843e57156c99fcf79fd8a0108ad25af8731380e863c7f136f303a88347d713feae3b84c4507907fca01564506898ca54f032f4f080879e46605b01e5edb1c871b956bb0e256;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bb3ebdb19e66d936a43a7682093f31c2d1542ec731f6f135fd76782ff69824bc9ff09b153ca7801563c60f73fa0e6232bd3b00fc2bb12da001c19463438d91e51d187a6a2c64a4b4f9343e49992a59452a6944240609e70d06ab9272218575222f2083f05bd4e9fccb1d3f441a8381e1b53dc6caa6017e6de15d9756d238fc2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h239432b2a90c8dd95a932cc648a3cdcb0abf6d87304651b6140f7361d7625aae73abcfce15bd528bd3f299989401516f1eed1f372e0364d24bde67e8175fff057e411ced4a76a673f771f959722d4e22027d83db4e5076d9dcad09abd0e2ed2660a59687bf83f580c6008ad144263b93adbf7c4c21c8d498def6680d1010eafd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd505bb8bac0964db78db303f5b394176dec935612d6a0d46fd2362a8402bd89a3c6c767e0994dd475fc530315ac465b96b0d0e81abfef9e2758e8b06c6fd2b2c3c515a8d6f974b420c2c84d38e81d7384173f101e7b4171d3730c9cdd6bc3481b2b901d265f2182f1985afcb2f6865d13e3dcc923c6f378b8230f4a338a759ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ef99b9b9cc7808a872b83a6d27bc1e6f6a77803accf7415287c2c739a5d5521cb75fe4e2687d1b60dba361d5ce682282446dec48adc74251b64fb351858dfd8afc1143aeb0a3751b3f4f59aa2bd8e6384da5f8d9713ac14205e3e085917959426ab4e6f8dd4fbc80c83e32d9779bac0021045ba555c8b65bb56e8059452013;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h366375749757184a6c3b5decf21757f19956025a9e3e33c1fe4e6a9a9a7d2e2e4d6095c5f4d385500f08050ece0df295024f8ad76c52f20ff2e4a1a090cbafd85dda860370d95f1075f83112166851cfc08e8a1e3863c8e3b77c21e98118034fa0228a72df5731a17fbfaec1244fc9a95e3cfe2d500aa85a1070f60380070c04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6ca6cad88248e6ed33ced3d854f550e512f120812e7695383b13a0e83d6a5c40b1c1ab864f90cc109177259287afc9fd281b5a90f4b57e20b02642e6895dde4cb5032113410c3518668687fd9833fdb82b089ae016a00f6f82b4fe4c6cec896d30c3377319611969dbf105a5a4369bca11bf5c7706651d3312941163acb6de6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e145a23741f1e3d817ffa38c46728eef4a72ca8efe1fbba635a86ef47dae2df1a3a6b4df352ac8311bef7656522c5f9c2b0ebf1130cd466e28f998530ca45450fd38cdc55d8df4f62e2c50ba66522731bc561d9752afea729857b566efc6b4b3bb6ccbfb3934d2d33e7cef74dc2d3653070f084b0c9b98ea2630e4232d48ef1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1dc7569e3703bc151c6c293730518efaf28ad8f36f3ae77a2ab57655ae2194400c432f3a43284c4d14ad8565ace92f9e5d1153e8c925ae086a4a5e9b8d95bb4edb8781eb6d2c1064b8b27844a42a5f57197643ff32c632a5f340ca9ab7e9d155d2511e9a0467e42ba56292892f4031a06ca7e47307f931e9aaa380ba488ebe56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd05ba0fba9ddc471c15d03de73d3c98f13a254c2847fb660a5ea408dbabf756686ba58088aa55ea19534c4e7a503f6c05ff0cb47e69accdc67f1f3e7fb667d6d91e5e7d773a26c4d5f86e96cf365a15b59833e1d268cd1a09876a1081081604ff616afe9248b676395512863286fdf59fa5596fe3e83ab812f0969ee3039f909;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4b40c0d9c9e88b2523d6ba206b776d566bd38fb93517e1998906ef359b176d4e7398722d4fc690ca300dd049847cd892295ec267b2a8d3f109ca64564fb60939a5832c57a6c9546b8d608052574621e9dc04263794aa87dbf146aded4bb595aaae8ecf3720e62719930091883b5ae7eec22f683e1edcc3e5ce45d25776321f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h430100cfb4bc797abd7f4e9de2f94cc51841efdca971c0895350c41f80bc04cb4b94cc400ca9a469e14ab385e375fc514a2eacd11191e0f35eda4028762b1156566e0d5355263bd4f501b61482ca0344e715f5e423ec571713d7c20e190368f354416477b07f2561fd3e1b358bfc12728f514427ca771d83c1195f4c73aa5f69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a43b6eb404c23d6bb32da0d024e35b382e9c77bfcc17b7ef2036725b4730e9a78de8cd5948ff49244f8ce97fcf6e6d56850d199afd57db6ce509910e8781e854ffd0b36be5a9f157021b3472b4c03d9b11c01bdd7e00c1ee39a1547cb0ef75875b7d180cfb3d59ea3119295dd948a8ebff4318cb221786a3adb7c099a0a4948;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b88820fb7c2a63a44b346b98ae1c508320c4cb396f8aae47915313fd5f27cf4c83be805aaa7dbdbccf7a9320facaf1794be68cd27636ba9c3685c22b10e4dc4d5a25f1033c12d63ac01831b28036ee004362c3f73840f269ffea39d07f33d608ee59fc6dc9e423fde2efaeb8c00e93ec5b40db73cc64d3c2c08be6f4f1fef97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he077fa8efa9d296e9d266842815f8a6339a9f08869198ff86104244e451a32b506c9e2ac07f350dde1fd343cc8f2a22b90f54a9e7b83bc3869f75b1f51aef5f4d0945dba1ff944b7311e7860a8f267e860b5f3e1f0b5c83a02bebf4cc800d8d5a715d45821ed98b24b9ff6911dceb65871e95aa7776e04193cfd3ad001abbd30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8d70bd9dd46d6c39b4010aa0a5fa61151502930080d05699cbea37f817b234669d82c88e7484d3bf68659dbb6167112baa3e441632256cef8daf57d8c8bd846d29f78ca82dc16dea19ca658bf1b7d5c452e3109bde38078224e7ead04cc6bf1b4187e3c482b1984ac1476496ddedd577a69437b590ec64f411cf5d09fb60579;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef88d2cb9af350c37cfa1b8e3209702a431606d95ba3f8ae0d2cff6702d7de2f2f8296ecdd6a51d4d96d4afa5b9367c98f2e0ad149f4d2dacba2395914a09e6cd68649c47c20ba99ed8d0459c48b46ded39a0e063643bb6d4bd81212a2acee77dac6b36444722d7b0fbd0e8bf9a6b858ac23cfcc1de03aed6743a65a8193c7c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8b8e0f79348f24025658eeed1d5c714dd4e96384ee7729c370556d855e1289dd55dfeef724e950f7d432dfebba5807e9856719854da5c61f881c8b19847888f8612cdcb4995ef4bcbbcc8c4df309301e77e664558fcf5acfd1f380bb1916ae541693b920054e86db5b872cdebd8446eccd64a2d8a4c30fc74d673813561c534;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h471cfe5d070a9c049ebea10a0890d161276ce66a6a56fc752a9fd395658ea5bb7dc7b3b2414bffdcd4e5334e6658ae8f8d60f3911ade429013d6eaf75c73407c5a9814761f6de7f0ae258cbc8788fd696ee7baf575211164713d18c3fb5e1dcb113719fae885c71730ff872c893759cddbfe0c90926bc1024ef86378a23a8335;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8edda7774240fa7f692aaf16d9243b36c404af21145d80c0ac6c0c9827778b0ad39e6392ac7c13cb8238ef207dcf4385937cd464848df0447295864799d9a3c05aed47f01bca133b4106d160defb2cfec442b63b15e940820867aacdadfafaa1ba7a50eb6a1904eada0d320e1496f386d576b5d05733e0bc1f62201e7bc5d5a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h398cac4334f71c2d09ddeea97cb69521e1135bedd7847068c8581ca645751a5f3a2395c1dd033e6fb7786b9f5e44761476a43c754b307675bbf59f714f2686b7216207b335befd81eb903fea689806b21d51d55b6146ddbc463a0163a6b2cd54a95f1613bead65ddd69c9efc37c669d629fe881643c9d556d53c646ca70e60d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae172e0ddea06c2e361ace8f0c46700f073f89582b02c4337f6e8f2fafb785babccc8a89fc267a3cfa83b2e4e72dee1127f5c2131bdb68c082b1b999ec80974416c619b7181772380566d8297013915cb83d75234d0e49832b868d62cb7114008b13cccde6c4de806685e5aafe3b2bee02a9c6a781c3ea5278460971d4f0234;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78b8d30627f846e4e752a54cc4a50f9191be006d600b8357bb048d58d2b4e8b0854829e2e711b9d1defc5c55f1dfcb4bb2aa9cc8a64377084b61e2c2defef7b032d613f0f59ed2ce4bc7dd9d64ca4d0425893e51284db74d3028d2d2822491c7e5bfa2a36817d92818ec9c1563d42526acebf68e2d09d10ad3df373283eb6d0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6416872bf2d0079bb7d92b7904a4d4486880218cd4415bbed62a228c09588af3ffb96e4542ad2bd95a5d95d81402263a0c52e94dd0221b421285d9847feab95ec5a39ee9f9d295b3edec86577253465abd981b027b17d83a75a34e0a1df44c898e12cd137946e22a6d94ebe0a6e3c9275f7cf8b99edeec19cd86b01c948dbb3d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc53fadd15cd270f34be825e68a67eb8df66a836e3e43987f7114dec32f9017bc84154ca25131622f6b6a96352b4f1f55b1d66df3285f11ff41fce02e349b683ca2628c00060cd9e05515381854ca49a71aa20e31b1a2ca0e8a8721fb55ef1a582326ffb6c37de6452bef2364817647825526ebeeb3d09438c7de9057f036e23b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h236b188f3fd7a990cdc4cb201c1a87ed5c1f58194f578ae1728e10a170b0faa4d5d482d4ca34e87ba0160655cef42cafda3ef59e40911de9aced6f3d954ba56d539882f103ea70a0c10aac53e3d589f33923515f85a307587cd630f9f4eabebdbdf4317d3a02d6d46f3f5f45f26629da32c63cb5db9b80aae8f02be1f15cffc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0a01ad290999e3dfe81a225c248e2916a4aff8f972f37832f0db3b1448aabb605e8908c304bb91b6d3e127bac02a1de7f3e453df2b02a3846a2cfd68a364d27845fdff5ac55ea929bbb9daa6b6bcb0291bdf30164fca3f2575d2adb5e0f6875c67f7e8a5de57d46c40550c560bd15f9438529139535b3b8138d307af2a76f8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e6756fbba93a43a41c1423a4ab399f0d164c616a4428e67c79ebf97f65d09c45265df253204e5f523a772265e20a6886606dcd6d3ea6d009b0484bb88dcd14d04057927a90cd9273f3863b59dbd3aa03917407d262ce67c1f6db54a50052e875cd7b8447ac9f40669942a432cdef7a07429484af700908f5c9b3315343cb6c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77a583896a1a3bc33896e8acdcdd34662ade87d4cc8e376fad0767dc445a09dc4528117e76e23866490470176c09f9cbc190a76e625c60eb697227e8181a1af0ef657ced9c8403b8d3949e4183d4a0a88a446d313a0c7d91e954eceacb5ad3d4c4d551beb913b2e4a19b0d0b6249d2a1caf1ca798decb9523b8a8a6708d23f6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h724ec1d47058a1747fbf7bbf139103eb6283b079d0ad3eea250bdb90b8fd76105c772735e03126ddaf479e41e35c1f66857a58ef1ac424c15d3a47f2476cd14c64fdc33a344550679312556cc574cce4fe8eed5dd6786183155577de40e42d6239b63cc6ee093341d12ca57917571a9c2d2d107a813942f942d1281298df6a9e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5ff6770c4291e2ade0230c8c0b8bc724723a3cd1e6c114683a6e7eb74acf73f09e33a4dd57042a23a6d24287dff2250ba4c5e3521b6789bae0de9a20419f81bc842e49245841fff9d3c0582a95f862972ab117a36693105c3a2eb1b860c0fb2c9ace7dfea9d5b0f4ea64875d5ae9ab53bd2aa105b051530a7e77309c0c5448e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed5d93c66513a905957d6c3e7ce1df0c26e15156ac2ccbefb7d8fbf667d3deee5d5a3b40ca86e8c17dbc2c71a796905fc361d89abf711fcf2edaa55a207e6e2d9ad0615cbdb5d79292c9b3b24376910ccef0258b2053b63b05ef7e4c4335dc381b5533ccf9823f7cde776ded4e952d468ac04ce34e5655b2c2da8d9aa2e7bc10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h951450d3de093518c5065cfe804e5f63a43d17bf99fe70d08a22d79bbb6805387c7dacc52c034bd850b3d37ca1d289cb47cae82050675cd6e8be4253fcffb07d7f7ae49885950fb3b911dac69df514ea034b024b4fcab5ca425379fde5eea8ea825b1c3a0f1dc10447e0c8bcc95a755eb031a7f750ddbe16d4ccb7dd545cbfd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha092b13594cece10e3d672454001bb9eed540645c4d0ac0478543d87cb1be4f23898505de8b0393f640237819b3779ba09aecbcb7e7dfaeaece082feaf6497a720601672b953bda545c04cc682a24c674a46ee255f543481260a25d0709dd213ae9ef161e3951e11dc088aeac7dc9bd975ee432fda9645c2691520963e665df3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a6cd913da601a75ed66dde85f2ece63f12a4d8a8fa613132aaa76740f9b76736159242cf99158dfa966e42b9fba35de97a3de3784ff04935939f4fff3a00f07e8fe37211994dbe93717b9d43903e2531ac4b6f1c8d0b23e35756b990d44e1c4d4d7ee3a94b414e4117bd77937dc2d1571c9ca7af0274ecbbed452f288f4c89d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1165d3bcbda3528289b8a85a7595fa7c95b874d11f966657b972d5af8f2100522d5e6269141e03fee05032134ea7019038fb8ec26d94fd5cc15ce4e827f9a9a030ce644b6d9c5367dfa4e5db166478b8b3d9f0ad0a440e7ccbaa44ee324a6f681ec988c577af5e2bfc41b17dc61a9fa6f9ead927680cc929f9032b5303570574;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7704f08a91dd0bb5f38061cb59aa9caedbadf016a60eee6fbac1aeff41a35341bc5803d236025eaf95c11f8da800a2f0def6610236d3899b551367decfbfddacfc329e2ae96c3cb252e068f88f8e4ea7ed2efedfbbc6aa227ed09eb712f91192a91ddaa8cf3449941913f28c5132b53a6af5c5455000352fb8ba1396f99c0b0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3acec0ea685807cb912960feda5fd3df3b924936921ca8d8bf3874c0e693f5d6f8f8b4bd60d6835acfa1685074aff3833bd936e142ab0e19b414d4266bf035ade1b183649bb80a5abcbb46f405e0196d8e7b03bd5440adfe1d233435e0f9350efe8fc4f788353a402a041287a61eed10203ba241b6fe37feebe5f93e54edf2d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cc0f2d87ff845b7322898e82c7d7c33f2c6badacc2a44390b31db5ce77158a2860f5d376412b3d10951daa6d3dfb22e88a72f0409cb42f433089f5c71142c627ebc8e80c4350786f9e5f6df9bd21f64462f323258217cc7071bd3d2d12c82d5733a327ddb1fa1a53b3a9cba7b5a4674e585648514564b4832b5da2e1d128b0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76c57b8a03cd17b9a93be4493ac884c7dc64f09f039ca62b8a70cff6cb66af747f96c9bccca7241e3a9938657e18b14eb1218b03d1fd2401e4d93c1e54fbd1f9aa1da0207ace87945160f0176cdb42669a39ecaaa16847e565a7eacdd85e0bcd52a94c4950ebe04ba165ef10ae55f4e3ce4765b9356eafe3d530f82a088a7d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8edafc8ea1a2b189c9b842b57e0aca26046e1f4a26fe294b0d0a4e4fde8deab88a1625e9bb9c3e835e7bf2d98c119d320f9a9aeee7b002fa1b32017b18bad8db9b13fa72c54f93295d7d55438a84e720d3f9d402f8a2266a3f6038cbb540f4a43b5e082f220d93f34d8c270cf7eb1eb98b3927569771781f4ba9bbd42ba99c85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e96f182395de699f1ab58e6184d0402db1c2f230ce61d5f908844ba9694c77095053db53fbb4aba6c628e3046f3690eeadb541c0defc2853d34bf3e18c991e15d680945aad42dfa7954561e432a473e67a18a370573e90e951619588b5f32173ab73ef2254cd12dcc8ff75f60c017cf7b1a2e2af8d035b2d78c1679e1a960da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8d92ebd70f390c46bf1e0e09a8b58ca1633313bc0556b0045215568e3eb15711d3ebafcd17f30b15b69cfcc68cefbeba09f7f11e0f2d4d724091c42abee2035733d961a9a73429b9d82b5c27934fcd57de1d255623f8066c32806dffed8bbfcdbe0bfc45374a668f2f3f4242e43fe4155b65b12f7170ed40ea84b8e08b99d15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf09aab3121962d14ff5cd8ada3657649a1cfae6a4d3a0c4af701d6af715f2daf3e6dfd990a82598bfc5c6272ee7c25b1b9bd6eeabf02aaab54c3197945273ae41a6ef3d0cdf6b97c5125161a1d23b1940efc0b217194ebf2d411a9c6bc5ba26933df028e8c01e9eab66585eb66923862023cb995dd87d90b2d56163b747c6eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c5f1957f8189bda6341cd1d793ba046f984e2cc0e04ced33a1ac0e5c2d1ae6def276bfefc9cc2704de36398a197a05514092f2a1f33557a634ec7362d1780f3b2c11730d09ef836bc555a340fb3b28edc310571a58e7053b99b8b75f835403a01db3d308d49faf42852dcfd5e234cb2c0f8e9efbafa21e092bd89c7b533cf8d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5838b48f05a8713dbb199e89c54a936babfeeb01f38dca9ae39716a8e634163281f70ca825d243cafcb0df63f1ab7249f01f4cc1b5638e7c3bb32cbba12b1e0c2511152474d97dc8f54019b30c12c5e8770d0a4b44de551965babdc86e382e657c1f463a6d0e9a9785ada3ccba113e6552a1d24b2f2a9bfab5d0338834c6eb0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h371fcafc07ebe7d923434c05b852dcd5a5a2b4b443663e62c8cfcbec663c591b70bd60d4d056a3633bef4f5ad0e7f6e8a87d4bf46f1841ae738e784199a32ecfbd3bbc9a1d964c8eb7582f73e4cfbe0682911687309ffa21c5fa1cacde8de3ce8abcbed4cf72c4b8ac522d0be19e65da303b53638bacfe3c1603eac370f0999a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha86b257a4450db0fe2194537d81da43ae8423ca7b93a62b56aad7be7d44e09fea85031f762a7510429e90a601d7912db99207ef023e0b7be27d8d6c950785659e32b2d94d06e370865c670d1ab8a5b9a2c1ae956c21c3f9f9db959996bb7364d778368f0c52e588da01c5a00d22866cdfbf4b546ea37ec210ee4cc7ca04927c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf09f27d7080106c2b68adfe3f3fc652a930d2d992ae927789b1bafd4bb15c830af68097874e87788b12587cad9e83fe3a2e5c5ba56b87b2f96ca6b610c9a04535a295c5e78f07d4504fa6bd130c2b5f8e92fa0ae77967937215684321bbac88d0dcff068d0b38e0166c47a763e412790b57a6bda21860bf23adc4e71273f1fea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae0fcc362276bcfe5f96542b69839c44db0b000d83a86ee33a1d8de79e1a39c3f437434932d1dfbc2761c1c0541b56aedbb432d6dcb298a3e696cdeb6101aebb4de9df01ef9baacdb569d27da917da52e663bce95bc30a621512bfb7f53c22d82c5db5244b792c7d250ac3473dfb86ac50c7a1e1b6d580cab0084e18726a4954;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd061853d2048c1cc71584bd61826bc39f496899b0f9ac6c42dc7771f016b45d86ea958bfda14fc1759286f569c879fa77f25181255005f7d09d1d1223b07154491ccc4ddc22c71cd0425152a176fdd35b133a54550379f89e0070d4f27f213115e78cf348018a41ad69d7c03501bd986df568a070073f6719db5b8db1fbeed1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha24aa48d73184dd91f701fbd79832ee16f53a87d419fab50783334c0414040bd678569fdf2a2b10c88860df98d2acf04eeb45e36e851603454837bbf92c0d9cef5137ca4a5da1ede66616e85e64d9378990d05fbaea9018c4a13015a9665ab07c7c576ff5170ff6a0769d82a83115587dc9233090235f0dae7d91fa4d60e6fca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9a6ca2f56c10350eb6ee92a5b4cf3ffd67275c1b05f87c99b1808819dbe1bc5478067a2dd31dc7617060641c5590bea95651a09d0c66569f2628bcfaba6f4f9700a7eb7a171deb182444950e7c0b467e0478e9236c7fac61f5f93cd3e9974a2e80c093e863f205a6f7799694a55ea540d158d0e113f3898d87dd9090f00e292;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a962c12f29e2b41220970965b0d20e3ec77c9eed99a7351856fea28602577bbf8b0a5239505be9985bcd2f59edb65d54cf2bf9450d33c55187f604ce5df7b3038831a24e4d1f7adbfd7eb0f16cd5a0fb94dfd96a77d39772959a140cb2c5ff079479d571ce8acb888ea6d40ebc01ee8c76d5e3f45cb548cac772efafc61fa28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h884dcb852ec9654f7409bcf56a654a5933dbcc85c5889e5bb74f2fbc64c34a0e0a0f261ec7752dae9f21220f7954551db193681f517edecb50ecdb12d595eae1348ed24baf264e2bf4842beccde7ed888162a6cc86d78cf7e9a12409e6492c1c2f146949a7e1b47c597f5d9dc518ee12f94d7bda4bd2ab94ac7f774d940754d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c863ab874a9c72d2861b60c58cdf297c1e04c04c1d78d475aa8637f3a4049252d7e2d4ec9254886b56b35696e47fde26a4b144dadc63b3471ac0b7ebf6a29cf1ed0c6f15e061f2b72cf0cdb41bf273a87de8975cc6524f9eca91f032ff2c5e186fda2c8bea5213a7293ffd3cd956c4576d200070b2a45bc9065791dc3035c38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c3743b392b5ad3daa42aa49d7719cc792c6927f885cfcc2b8286f100090a1e020a46861b9b43742ed5497f1aaf28b11b72739c4d68ef1d741b9476f43f3a6c9d363e7d80ef97e01dfa74f700a06fdb68a7aa44961ff4910c9b8c377bedbd87102bf4f4ecfc7188b9467abec85d5ce57cb1f50d19dabc68feb28a878f0b53324;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3336ecc5240973c14994d276697a08dfa975373a45bcbac71af3b20f2541d44a8aae8757b07b0182548495e29f9dc25d1ce66b6f49d9140eef1e2ba32901628387a845284b4e528d6bd035c6e6b94c23bed6b5f9d823f8802eaa11f2b95df5337553909a0f81f205abc7664021a27167aa20d2888d343d06f1a5f807013fa75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he404b4ed734bac0fa77651cfcdd15026ed800ab76ae9414f4bc1cbd5e6d0aa21293ce57d82df46c4c8151a0a360bdcc8252825f88d89f645c7ddec08eab222909c88dda9957733124a951854d525a054312aa274bddbb267341758c291694fee394af8e3088290a06dc2fa90a8f79ebbcbd0046585bb0df8279cec7d39607db8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77d74917e7ae09908629a5b6bf93539914627968e3a9d63fa491914162044e4287ace07759ce146f2693f4eb53c022445d90662930856b96d4e40a01cd62fdeed2ea0394033e74ccf463727329f4694508f485f89340f67335b2c189ce2574e0cba8c4dab9cdd7e6dae33a18774f7586a896eeb4b64d28191a430b6150ec2f6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22bc92c06fc7a1c4fdb7c762d600f477e0f9ef18a0669c66375691aa0fa9fb7a2ad7b4f4dbd007b10a1f793bc6517d32019c303b3b3d6c4ea4c2c5b60bc70b5f71537c9ddcf5c45dddca23ea843b0d91c5912a951d51b8c0625b2188bfa76c04490c00187773d7924e2a036e0ebaaba5bf967df3caafff698bc094e96b6c1fee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42babb52a2debe54cc3c2f0137acaa4154c5078fc3a779302562aeb36cf3ac9c279a3c19aafafee75abad8ef1ad399f558d2ff3141186df7a14a852c331438022579b9d9f8ae189efb393660e4b4000eda3e062067e59b85403800cacc589ac1c1949a084111f27a18ffb67c558faae7e5632b05c924b2bb0004d14bb990dab7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8939d6534556b71a3cdac58a18a9f07a77c9eb51c4d45d12b5eb73b014219bddecb4684ad0cf750723c92454e19461972e61be51fd21218fa2381ee21924b9dd90a0b03051d3c855990ce96488c466d5f44b7d3d3cca26410cfc1fa2d39d4f0a92246ab1094a8d10b39c17487bd0d73a209d093326eaeda65e779d7b1773dcc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7051387531fa2efbcd5c6a02931dd6cbb1794eca74e2c1df863fa294c7647e388a4212578504d9e2e31a9618ace676717965a609c0f80970b8c60312f3113f72b6e6aca5029df74cb8739c15bd4c4725e6e313b9b60c81a0efbd3787a87ace40d7969bd6a3de6edd540ab67bd08d798547372ae3640afce51562abb83bc68bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'head5ad1ad81e2228052437c826576b21f1113dd623899e55fcc2aaa68ae49903b054b46cd81acd7b45d8d617fe0e68db7c5691d988eb18c416f634a7688ba5a056ddf58882c17087d98aa88f342d05dc70cb7eb1785bc4619ee9377ca838a9063eaa80c80dfc5c1dc051b0526b17f88dfff20ef7efe8363186d4f452823edf02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62fe50fe108dd762153dcb59302e00a7e8bef16bf08e57766bdee82d2c1faba3df58b3bb6adefe248eab0946dcc13fddf58ec4fed2a9d44728d8b5df68a12d371d59ea3cacfb0bb7a48685431090db2dbb79f9e8595b38a30ed8f38006b7f5c1f384c3c3a6a39211350fd3434e53ea2237e47419d145d81e332869e89a10ee14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc04bfab2bac8a8f6eb842bcb9a01aa1a482cf3b38ff13979da69116d28dc1de297ce841f0dcf6fdbc5c5f477931f3f77f160b8a410f51ac740c82df9ce7f1e17f92fb9550bdc179c637e1102a20fa525abbd1265f67c7d26687d3fd5dad69d23bd18bed9bb5faf70f2a689d730d15925fe443dffb1fd3d4bef314452bc603a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19f1f04364fe5f06fbd248771720dd03f84f33a81b066d28238a9c222492a19bcf9650918e3522bf015880705cecd9ea2e554d8f7a193ca8d7e95d77c26ed5cd7572f9040291fe4d9e2a85d2c7a8722dc707a02ab776dd1bad6d6bb51e62a177665f7ec054ce2a000489f72065a28150d242a4df25f934bd5327ea4bddea81c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cc52c7bfe04f72336901406249a9c23ffe214399cfe6403c97d698e5690c6b2c3289eebad6656a11484c8881989b61fa880617e3a5e59e65021e7de8df1ef09eba8647123c6bccd0d4836eb05e9d739171dbb8564b86811c30618d38eafc40b8a8c8a58ccbd8bc6303e9d83e0d97094685ad990e962b896994c37a59fa11ac2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c49aa774d03abfbf0db256e2a66f5687463b7f56935d8a416b9f0ad5d360a2516d112d97e85499cfb0fa1b6f19b470bec920dac722d91399cbc5a4e66e9e127674fee9a83d565861f755e33f943e0d4797aff2ddf90661ff9f19b68f99c61dffe27e82fe523bb9548b23e464b02c834a80394de7130e5eaea454867f5948e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha77d1436aa805055ed9a01efc82dd37fbffa4b30ed628cd57fe3a6651e665c2cb5e002fb555a49dcb4f95c8c5ee084a616dab64508c8d24720fa077fff39c745090bd8f70b2edefe069d3ab68b8758259d59445064512875344ea57701d9eb6450e342389411611a86b0cb39f9e7962b5bbf06a0f63fbb3614d5882e601dd41c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e3320f2a33e011c473d424c7f0d8f8a824ec075080ac529055e73517118ea6a764a9edac52d1f7ca5fdb663709409b5a6f608d3633d6bdb9ef771fa1ce4f9fc9322f51c364846a454a45e4970acd23d27bc4824fd2ee7ff07875c0eaabf2baac51f1297288ef905617756394a6f17b875e8f393fbc8134083a0d0d8648f496b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a15389f56006be005213cecc13a4abcf979cbec3a637ec58152ac6128d598c2b6e92f94b6699eba9241a2970b8731238952bcf4db3991b753ba2c0516f6344fc9e00bdb0c7f2bac472c636b9453cf8d2c05ffb7dcca018a11c57a0ebd8d5c5e8dfdf0966d4ac4d2f11b25e0b34915881bef99053358b907bf8e6fd35c8435d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ae398840a7d01c2c70c320d58c1a576bdd46d62175ab5e01d759e159c1b2bb05fa8fd394456446da35ede0d2f60f106cf948b8820bc9857c87724fe7716cc133a79e2ba868fa83f2f7a0f967e0e06b5efa29e7410af71ef3926aa2fb8cf5e59484a07bbd7fbd2985dcd4aff57a0243f812e8410574fa82b1ec72043d8e3a908;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4590afea02aa7efd9208ab805ae1c2c32cc08f617b1b112b51754a7ecafe9d83aceb13a6ecb106c1bfcb7fdd412b8d151bbf85f2adfdc458aa291c9fd4f52dc3464837391c31f3b5133bff142ab9edc0fe4b2be8e9dbc42e5a66e8e3d0c1af43be65ae49aa305bdc17418ac9c0998de8a33d61fd83826e2da061446d569901c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5176647126f61430a393978292b3f77faa5c33f9e5a0ab126f095e9170798a4f67795b160ebb6df01f61d39df84120961216f822ac555b89f535cadbc3058628625249aca7e205e1fba4ab166953eb246c40b736f84f4fba8da16df16750dca2de8bd4e5059ebddda31811022de14fd7d6eaadc6082a9729d6f8514474cb9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he65e4200c30c2689f69486220a409d4949bead2509afab8a49ef9978688558c5ebc3ab6a903ce0e5037e771ae2b074e651b37b691a12134bb4e894be662add7e853d297705cdb2855ac7c9502ef753eb5138dab363daa9b5fb4b1d1a4fa3d4e67bde46a1c63c9246effa4a7945bcc7564325eb780dea749c45f04c7ba125c8f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2baed4267d57e2533601de985fb690f8bd518ded49d962a8d7f7aebb9c85dcc1df758df3e55b130dc359ebed6875d58909d4eebf4ed38b9ae19d567f0b456da2137f5310985c08a9d9c0012d677091fc9c49ba9c91a53c1f7d5e02921fcc7803bcd34c94b153fe594eb45190d96dba4d6c17678da203fe0f2a3b0718f22d7a56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h708a1b23a42301747c28fce9c5b7d0f93e64f68e5f51412415bb2b359dff4748ce7d2062bc527b54a34380591025fe71a07d0ad4b9ea0c26b83dfd9749252a8a014424d29ea2b2ec801dc109e61dd9b47efdc4a0b6934719cc173a90f66422963eed9cf167a0139c78099cc29210088f4871af053fba4c5b66d860cd5b97dfff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0c88221cdb02fb50b32d59df92e9d4d98eb43c17e44450a58aec9fd462b70d857e5ef13dfd227c21767777237b06303876dcf114bbe41b014b1893495de590a053bcb2deeb1799b862ac12c976aef1d0c08f5feb4141ca44fd84fc2a463aaafa44bfd07525c25c22a99ecae1fe38e6f1349c17049ffa0cb39e383709a2da92a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64f6ca783021a5009f5c393497e9e15e4b195f957e06c66ed2764b4c210bf9b17d4092eef47a9a8dc39cebcc678fca9b9f41fc44603759cc6ff2aac3ed70933fa8afd3e2065f9aba57191541d62799780b417962df79ba976a54d3904016e43cdd15c185a0c41b935cb9ad1028d22efd930ca8b41acbf0e204a99a8c96ba7638;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb1e7cde5cc3b3443389e4a6b5d3bfaae53a69c049cff1e8c99c41316b256fe4cd5cadac6c0c3e55dff01dfbf413fcec80cad5a1813e263cb06f5df1f661f0c0dad5cfe23aa0e1d4df5e9ece1766533e77db5ccab2902dfdae24476e93a884abb0319b3532a38480387df1f3c55917196ec6dcd741532600fe1a5ef5a83f6dde;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e6e6b250ea81184368a85aac5e990aa82b455c4414a558e1f8a942fb4c17c10f3dfbbd6d29788da7c252d20a4689184e97442b82bec3de145a7e85485e9ce76b305264d5143668c6d0a4a7ebba85fb422da527f54808747ef8d3f7160b511c86565f2cd86f699c6aefb7774ef6cb8ac53bd425048be0f5e40f06d213bc221ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc0aed360568fc8ffdd920150eecd183291797bbe706c0761df42d5b83737af6fdee849c58a8d7457669e91366ccdfc6fefac643f1237ad60c70a25f61f7a0b4cbea866d19abc8d12dd777251e718886ab77b9f99f90ae069a4b3a389af4f23297842754f6132f36e5b389005d20678b0490f84ad31effae21dda520335b6fe1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bf0fb79380c9e61ab297486fc02a8817b38dbc1d7f346b8f63e90d273dcb9e46df5b60e8d67c4f61525a153836f47c3b1af4fa06cbc9a7bd13ee6318b3e5ab3ef09479d44ce000aa196249f2723b572241e2a3f77ce3247b8c6b2d150907deef8e34746865c8f0c888ce9ec188b174b10c33533bbf2a282ff629e9c0e6c7798;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36ca5e756dd818439f4e9132589182ff730d78f44f1169623238e15f32970245bd05566fd146c2e22fe070d2f18952122642fd4e9ec196cd7fb756d30f1b94fbe69e40c95361a82ed68039989a4f0a3d76845274d51e1509ed1128370f5494f605814b85a37c2bb61b045bb0878adb20cdc33f42f245b875e54c61be6454b291;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1ce119d413f5e538670f48514fd76559ba9149105395d5aba65c4ce82b7b94ea3e7f36821eb0f66a8935fa609eb51bc7c632f374706d0db35cb585cd5dd76498ace9a7fb6ef7e81dc84a7b1e4456972de710bab986edec1377cd23aaded02521be050227e7bd7557b9c2f9c7a3e11d5f1adffb974810cbd19d47ed05d850a0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a3b2f8a0b5fa3fd83c2cebc8497e21a24a11b331a422a00f014b6449ef88a5269bbca3a2200629144f5997c1bf6a4325ada9da02a364be3d088bed43fbf6ea56f14a81e03a7339ebe5f9f05a8943067b9ab000f3404024a657daf56e4ba466bd8a9bf1c5c91a4c2e40603a067b83a4e357cb8187e458ec0bc0607c6db1b0782;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h944239284cc69a5ca97aadce3cf760e74bec97888a8c8f8da7f5b7b3661285d42efb73caf9e2ee2fd47ee3c21a7f2b094963e73696975ae145abed56f52562f6dcdb2f3cf812d0425be8d1d682b791960b72ccdc84061bff23990a761215a016cd241dd3b3d5735e9776cae8b7473002d628bd5e2203f43432e9de430b465078;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h830b9e471443f9ae77732f5aa8f498e92bec249ef7fb4aaefd9e605fce1013fcdb7199067ea620e2c846900ec5e85cc6d7886cba1095908a56b28bbda25ccda001864c50a83263e0efa058f02515e8af94bab744eca5ee13d876509eab5553263f3fc2ee80454647d3dc2f2c3cec38f30943c9cb108c4c97065cecd87e6c2f18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1123232d9b52017d51cb182fa7ea1046f1050e1a3756a259a8a87f287647e502fc7bdaf675e830febbdbc96c2c69a681d6d80637d202bbbbd44512efaf2e570a27a81c303624105f3bb408f94460b94e9cc3af01d62ca31ef6db660db45050e32dd47723e074c62468fd25bcb6c26ed16945169da6e44a347a0494f2cdc2698;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f9ef8f608758cca40cec99ccce18e834cf35ca0c07255aa25d28cb031d1d73fdb9e76f616476ae11e412c3dffd0bb23767ce6fdef9f4c3d6e130970d9fd8d85ecd7993b7995d696d1a91e0266daf8f7e9f756e5dc3dbf8f84a04fd9d95fd430388b6f952455c84948e2684a2c62e9958ac1d3ec81a537c31150db373e3eab88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a24ff5c8790c84aaf9dd29ad56c9b8fe713c27da03673cb3f56deb9e470061593329119f3941e77c476efd98b1905e22bc4cce707cc328004d856b9862db3ec0b1186f4f590621fe3eb58128b68018062572ee6155179aab3b10e6f5659549562d4bb9ba8a6aaa11bdceeb3cb9844c53224873606f6d5f0dded27cc6e5efb4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d7a264961c7fd2f8a3b7e89b7f9ce7761447842505ee83ed00397cbaa1c3cbba02991d26af33a024bda55680aff171e132600c31012d8b044dbd734e71cf8fd730160aac1b82e854fc61c3e8a9371150937ea3a913ee1cdacb02daa0f948f209d658817f00b4c82445b04159bbb57e609158ae72e5fd875e6dc69c0342f06b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h498ffd1a8bc76bc29ea3f06dfd2c1cbf45468677344d02015d7407838d7e23b2fb160085c6da35f7ff7cfda601f3c0f8ab03ea5fe7a9ad9af7553e36ce196ef2115887f6973dad10bac734fb8d615c09d2780b4f78eb7108817de6bc1c279bdd4796fc16ac34cb4e3a2a31ebfb6c4ac8d9cf6f1842340da1da8b1ff104ff1ff5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8fad27868cdd5acb2d00b724bb5998554246df9addbff8b70093ba52ab62e0802938e8b67b07d3388c7cc58b352fd2735f1f38afb621110aa28c99f0ae1e70ba83c50dc45186d645e694674a375c70b6de99587b2837c71443d819963c620137f7073e507220e3954af64fdff9e29e72bd85ae9164346a0edc812d244ebe10c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cf18d5dab37125115851266b82f3e7ec5933c05c5f5f08f809ec805ba432bdbdd1a50deeadf40e2863a7562806bfb06e40ca43b34d0414ecdda6aac46b4e1c07691f54a772130ae7c5a2ad0c1ca656500855541b1da8e767a3e314be32bab106eb70c791c8de8406125c1e2feb72976dd54bb6cdc3d5dd31e48bfb096cd78b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10a6e9af85cf223a94f4352fa1e38283a2b7fbf23afb2a0085df53774a4e1a36c0dde74e6d536b35cc404278a97087a83e0d541215eea5b0b16d5b1621fc91616868fc084e1751a5a3a615dc252f5b3c1ca122338d82cc1cdb1caa26a5826fdd829c85c0c8bd328685a9d8741657907a257e5489cdd6397c92dadfe775d8c938;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80e2a885452d628d0fcb9b77a93d214aba60698acb430d897ca1bf06477179d0451c76e1bf37238d740160bf3bff3120973a20dd3ea8f2d5067359cbdd08a1db96a77209e311de3854dc12525e08d4b51b3d10f35f429138957e13d4d92ee22888d99838582bf76e9c8b4a55b95cab28967cc9d8bd8919abdc5270090c50c54e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b418394e4f46216b143370285394a2fc90863159816db46a199bf9266c441cf91542246b3627bf99606ff3712df1b4096c5f9565ad40e860ffcc851aec55e5ec45810cce0be5d372adbcf7b0615c96c7256f1040c2f30f8cf5d7a57e72d030a34733974ed07acc87ff791b8f0e271cbf58544ef0c7c63742feff814d0c506a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc322ee1500754b909fa99d173fdf0f25a194bb8fff4ad147c189db776742b7eb3b0db79f6100324d9b9a753b5227bfbc741d1fa30cfa12613871ec13fb1f621883251f4d3f9054f42513a18e2714d68d77ecb034d8ec59b643f0006a9e42fa37657875b629ba72b6a75c19512b8154b2ce5938686f105e4ea04f0bd507c006cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef5ad2408501b8aed95064769d282084e4d0d3f23c367c96c42761151931e77208b30cae7e807c7e73bb6c025c3fb73d10ed6e886af667e29b93841aea89fc1112ed4a3a1eea75b1fa2b7ddbc531cf10a2002316290951b6dd689075376211b20b3ebab14b8f6fcd7874093c087a4cb91db8620ae5c8b1b9b169897a37fd0e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h819ac2e1603aa66941a89462f0b53817ef7b5a723baa58666f770dd50ff668df0e05f29cc1be5f57f9768b6f1f25a4e32340d13182dfeaa5e2c07322a89dacd47de7a807ca3f2db21bfdd890b65ca0ba780dfd0c2aafe9ae8acb258a431e1ca1ec7d164e93613e6783065aa4b8973eb46b2391d03887307bcd0855d78ed2d586;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5844e851be98dd9e8a83318991091589b9af50dfc2eb887182c043c83de72edc89adee5055d12b4f8da0b9c8323f0c6f29fab9af6a91cbcbb93dc8f938ce5a7682f29ac58356bfd1cf93b55fff96047defa5c62d90563f371e116167c6d02c7eb05b96c2aaceb550b16e918758d2039e535d74199b19fc6501a5fec369f7a2a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8822cc6b1a1a2ef9665eac855560051ab45b8173f2065cd2f54ea096194a19f319f87ba6b46cf8161421d12c805c85a737a48eef9c161d6c1f503c9969efac20eb223a35c478f3ace10cbb12ca9a4ff2429b9a077078456a709ea1d4c46889a7e787ff6df3ab896d2e9f5704983906a7fcd2cc926f773e3284d454da44e89905;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haba79c22f661b93f21545e5c0c4121c6af958e8b208ac28db5334ea7475523802f56e318c5de7c75c1a87dd1db32d5d22e77bf335e217d4eac790997becf1624e169cfa110c2831051686fa753156fab7a1921149906351132d0d8f83f390907d6620cd4f66d13cbd872a6f01f3b1e88d3781d8a140c1972c4a7d0b368fca4f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91cce8ffe7efcf660531751d3fb40392127b13908f2edac8a10daeaa733fbeffe3fe7eacd77b23a4289f088171df9c6a2cc8b2d64bb22d8aee9329d6e4e1ec2e1726948608220c41401e77597927a05217841d488c4ba47d0928c46e41cec935c277f7d8c7b345fef0a9a82d7a3cb2b51444e19896f2b3202b6d762d070d98f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58606e127fb9ff0f9a07f8705b3dea1480dfaccd496178252edb2e0a30bca9bfa9321fdd9830a127f6c4ae9960d38f69df81300918bd4f9a25c481ae894fc7e7e11072bbe11b466c5121b6eb0c3d0e6b0e4f2e728e6da446ea44a64b2e32aacbdd7fd6d64e5963e22c1ac6243c71f360e95845529cfa26a1cde5b81895db1547;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d358a6b00bd7ca46f36ee72ae3f913a4f6337c08a11ceb7438a9423ee87e9011f402b6dfc6db1e8a3ea24ac9a400e451bc7763fbabd0bd34a0b5f4200ba4b40ed8d9d17d809262f5ca89d4664f2515b18254dc3001389818530108545a50b47d56b019ff7864af579000aaa443c84148b2d26c2fc5d1c10c9258bd4be5fa6f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81cd50aabe173a04735529f18c7b806d065d627c56e607a2e07d593929afb2fd8076d32fe914b14c38e6181a62f7141923c012442fe029c48aef5cb3f07b04d93968caa532124e8d7bc2dc452c0eb0f3e88755ac1c63b5908645a22aaf087f34cb312d429f0ed62a6cadf0c43b3cf09a9e7e3be715c8790caa7e875bcc35f1d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cd8462608286ecff94b94f58e592943501cbf01657145bbfe10e22d3173a1b99a55d9700e91674ccbef94cedba332b16fcd8a16c94c526f592dd62db8da60aa3fd671897657a28a44defc7663fc4af79990e9a6814651eb6eda19068c223b97da731761b5f574f6fddc235d2078c23ae1f769f79cd68f61b40d0618ba7df55f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b628bd607475919ce7a4b0d649034f5b725cfcf82cd2924b578ec7cd3db4666db138086efa61b7f19613a6c2542d72b8cf0c55cb64cc5f4b420440e64705cf05729bde5480b7340e3477e83d154645944dd0376ab01346faaad6f5a6287290a89f4e655b8f2e2a88848b86af2288d88304e05f5482b722f78b7f4600da5f427;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e7fb6b627da81c675f7c2ba17aa28d31c993a050ff5865e86a9123f648a1f1be9f1af4dc562f371cbaebcfc820ca1950fc567ac9887ef33dff3b516f2fbf41bea44a43e5d79724b036aad677b9c56242c6b81b288ba5a2fe40b21228f444a0ae3ee8c053b06ab5b8527248477daa949ecd55c57ce9fa3645e3db3385aac5648;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5df1f81975052530306a1d246e7ae67a1430dcdb02cb7712c17cd70391fb9654285199c3fc3c8a916f90e96626dce19da0dcd62056b741203fd97f727a4817e68420c063dfae06a667210bc5aa030b42246b4b3b7c1fcef6a806b947df5c3727f861c7cfb21361a48fa19bef0e21e6c520c97aa06fe705634d4033f7605e5efe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf5d48ad34830d612cde05d5a4c09b640e0d45d8f7516128e4a6228956eecd89eea6b28b85fcf27f3e2f174fb5739cd3ed4e1f4fd4a7d8f131f6fbb75b69fa2fd1c2ec902674d125955396da05fa0df8dc0cbce3ca0a332751c434a14b03630b68a50fd2815422a66d59257e7e15961151d54c6559227083a51853d80d6e2547;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9008743174b3d09a426764fb0cd176724650398f38b0c53578253c4199d76ad084c55754e1fbdf090ee35a6c94f40f6a79de3d781da80ad6a98067684ce4fe270e3a3f1cfadd2c4c889461a21a293aabbb82fd0654e8d6362862e97b0ad268fb058f7b3a3a5cd9eb911ab6918022e5cfc5ccf8488e8dccbde758a5d45b651f59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbf721cfb369cd0551283b308d48558195bcc616a915a95ca2b07cd92c7a3c5f8e0b91a72b0ff9a058783c57f21bd293e614ffa80eb2861192f8fe03bc1aac846ed20da4c28fbd63321f24c10c09a59214a81e9916de7a6c3a16aa3da8c14772a5ea94b16f9e35794cb80c55362e95a74d2ac0cf0e3ae2951aa4f005631a88ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b72889e19cc8418ff69f1dfcac986f7173e3a9a5f5c65fbd6d28a70db80d294c7226347825d30b230e315f8057ccef442ac5d71bc00b8b2e27dd604396292b72560221b60f9bf37bbddf2bca425ed7a80512a717b6919e145d915c80f2b803d10da2e9a4828f30db88bbda64613e641deed65d0ab02f4c081c05b6336f11e50;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1969bab57fb0ee094d733b6f4b2a48ceffa83e37dfbaf97d8f15c845d830b931087c6401a59c9249718b29b3906237fbdb93ce7edf4522b5d788275058d9171c7ad6bb6094df44dd79eb5a9a20d42135cd2708e3d326786da8791ef9314a3416111f2404afe37219f4f8fc75784fbe06dbadc5df48d0b66eef0e90b88aaabb24;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb3512dff9e10b3481454efb7fa76b8cd444ac96c953ffc943373a254aeb4becced322057ca062488a245fd189fe8dcf1160b1f6f1dda4b4dce2d4a2f2331059df4d11513fcafbdb5eb9c0035cdd77db56ca43b3e556b0ad35fa49f7018e188de281cef14ca45ebab41352cabe4f9dc9b4c56e31a0316e740f81915d96f62ef5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h274a298d7dae77f7a03f48679a14b3db446992bc05c07b34a0d56f3589c14b9c79f2ffc346f31a2d9cd99e70488cb1f646072221a50490c6b66cfb48d1e43050d1eefa2bad654bd35fe9fdf9121a1d70ede9e5c9455fd99db5e22e67b24b9ede6a869b60ea0a28d60ec40cc6d8f0c01eb8c213fe685b6ad99322c565106d68e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h432150c81e0d5645a758063c8e142515d8f524ab598fdc103b497ef42b8ac47bf220f58cc1711d28afab48a454ce0b5201e6f42e634441a011cb7f796117d2e5c743fb64fc22ddfa865c36f99184559cd501589466486951d4e7f2ecad0e0ed8a8691862a2b633d64ac14757bbf7cd2725f0442f55e8177902b9408ccea446ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf44317a4a89a3a265b7a13336195f9e8303245dcc419046f7613a33ee3bbb24dee243b18bb417cd7c8eed7b5a74faa20fe4198a85b097099fdb77cd98c994f4efb3ce2d579918fd66ceef70804f6b856b5baf033763417a72faa3b5b2302c9db35afaac391d2f3cc5fdec6911ef541035c81f9dd7ee0490c2ebb30122849f372;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4aff9f401ab061e40705729619e63e9d6d41f3b3a0e7f94cdaeef0ab39e7d169aa75736d5015cff0175173bfe0069844eb389ef08813476d2c9c7dcc9d58243c9cc9a329f47952d67f981c8f4af3962b3008770654ad7c2c919bac03d0e3a8da823fde12dac812eb3716f89db24dae88bef0b59da721f21dce2ccd509c274386;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h815e78252339159a1a2a6c2832468bd11d6fe27810d2a68710fac52bf491532ec2d19a8b3d89d8a250a848fdb1c83f62f60fc7cce28b726482492d3720f632454281c2adb4cb1f317a87251136b234bd62d82ec77ad47487ac63f6b31d89681b431ecfcd3798439d6a62d5aa200b1fed3558a0b54df4d35e5dffbdf5418e61b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc906cf8361c4c1c90ead40c538c90f57f61117b1c62810d7a26114456ad45f420d644041d6ae1afab443e461562c5b66e2d17b6f33cfc38151f6994465ae20b4a1f2bb9166335f85ab60f9d0e5e6f5fe1c2686c26d2316c1b0c16b60b35a679ba0949aeb27f2afa379b5eca730e87d8b3328fd16ad65a80785194011601b04b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e1408805efea0cc0944296b8ca2ad8541c271db0bb58bfd18387902447608c6b6efe6627ecd5ab0e7da2b23c6733f93b9150916835f6e0ea1604da96719c1656d8b847855366677c8483b4f31655389f915f52e3165a4ae5df7298bc21030758251454075d788fcc577517f1a3488ce59c568ac435b211544396d8334f78dc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8e938ae70c88b70a44feff62b104227a7ca6f148cce341d3340e1f333a9ceeeab2c1a9d28ceabc3ab242eea5b4aa22299565abe88e5adf497e0a3bec0a44226b48c1602fec7554671f70a88cb1ac5a481bb7e346facc2c35ec344332e74ad0bf5a5d23da8342827ea9319d461d162b7b408ddbab0f03aaab914a860d06e265f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h930719dd559fffbe727df06c1e0a5ed3240e12ea4c3354017505ead4187b53f3ca195df09034f33b32fc7e78500d90b1dcd092ca7d3496f237dd175dfec5d68abb9fdd9b1e3d311b8f02d0691bc6f1de69e7aaa49a7153b460b9a622eadba91a3158025921fe5cd41d3b813885268433e7e1ca74a2200f3ddc277f41d4bc7dc0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac8a095104851e2c1719de1a331d82b124dfd1e2bcf040846ffdd9cf441c6f41ff56b1fd157dd0b421ca7dec56e3d9984e0708b9c5077044f13fcf9902349ab8b6c0468f0d18b555fe6c3f60950b6c8e4038e4f541cd2f4b179910ec6509479ba97397d60b5d75bd661694c627376e6a9433dd88a9985ab12759e72f66208bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d705ea45b020823691baa0cf84c478710e3dc8a0137968c08bc4485823b5768433b24cb5b29291ab3b0c62048512111441b391979f79a20edb3e711983dac78dc12c89aeb6372faa047bd70c4aaf4d5c9f27f85ebb181a3ac15b8285d0d1c13267437a35a5db132b13544418b3e2f1cb3993c9a5b9c77de946b555d3fae74e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h788735d5bb8a3b83a53163f3d83d2c3fa1371773c698592cd20e492d8f08aa8fd0f1674bb2f79bc44ae35664b367eb818c686718eeb0ce81b50e9ffeeca81a314963b4227b0f0af5765a5e5b7b1742c09c3e83586d30860cfdfbcf8f756e33478075255771f6cc97e0f1d04370e30e6cf6ee357cbe66cc569cd9b1c446a0a7c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h875ec4157d9e75b4e43d068447eddbd3d77e88f6116a3df1283cdd49c27159ca926fd0d3f221a84b69971da6dabcaa30b566916b658a15f44da418697033be5eb012487ff81246802a3097a1483d90139eb29b82bee01fb754c332b2913b66095faaf7882537797afbfa2d68d8d80d945c7f2e2f926e7e804eddc24ee9504648;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2c95bd13b818e7948b8cd977e86325699b71a947a5779e43727ed0cb5e2b3dd61da84a91dae92ef406c5b97a089ccda798f5ae746c6ad04d8362ae37b37b91d61cf275aa3bf733d40523f214b82b24ec440558a1cd1dc45a8763b056651e016a1b6181e509485bbf7a4b1a68c46684b23c9ccd867e537654475a7d5790a827a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc765d5ea7fcefabe577ca2a005bb968d07110f78bc73412d7900b51609fd035a754a18f7ebcbed3ad6b9e2d58b37912a70d19ce44c8a6216d0ee2c88aa559dcb8804ceaffa0e911485ad7f8b4fcdc350c6d43411b603fea2649136389b416ae2d805d77ad7648cea76caeee81fffa2bbeac7f082138a8378fbcaf9910218704;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bf48de3876b97a43b1c218ac9761fa00fa5d077d7dee2081be23572be43faeef56a749086c5df9928553a217f7c954649866296ccf3afaf9b3638904560c0f9c085d3aa0a8cca5bd0945cc44cedacff5609d773d33037ae04fe892761dc88353462613fed70e4d1dab35c28ce7f98cd1833438704050979008c6cdf908aa901;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94012a1b7f613222cb903d0bbb588a6ab4fe3672bb8e3561a5ce7e1dc221ec51c66094f7bcaacf70bede57d39785ce6017797b3ffaa4c779d7579feb2710565d26848144541674cb5501686f2f552bf2c19d8b12fdba929975a7af7c09d026b9f94ebd7c9c0483d8df186122cda4d689ea97c5a3747cd6087036df6bdb0ff6a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ed66b4bfe057977673e8e80729bda106b584eae1e26a9528faa29d1faf49fd303093082900c973131acf16b7b76eda0efe83d74e63c653a9fb07dc0fec2af9679e4b3e41992a9c48ceb0a2bd42e6258f372888d88405b030fc9b5f312c72e7bf0c64f2b868a463dda6935ff4c1d9dae934d900e2146df5c5834a63a85d09334;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4a246173aa51b9667a10bf229cd2ef44c28cf17b9f856684a3d12b9ed1bff4304a9c847dde777d8d7b7cd7fb1ae1917a3b16c8d3136de9dc400feac924dc87254df4375a1822255b238b53905e41d56b0d1ba6fa1104807dd551cc79b90ba11b29580b0ed43c9efa3f09cacb9b3c8e586103a40ff2ae9d2cf7e94e3eded3d88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab6930e4fead385e0548aa33398c952492dfcdfcf0f1b83296537a7e0a0548b44a785376013575b6b103f8e7679fafb3d0926a6fcaae6a716c77a27be54732ee8132970d447abac573c695a33cab67f7ff22881a2ff908cfa178b3bf19ae6e07ab3de422dbebe38e476dd245aed8059d38bb6fabbc320748a1774b770bfb0b37;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b4c184faa93ec6dd55208a95c7c18b314f4cb74e8624e4637d3306a5b24db3486b4dd905b965cdf7508e2663bac848bffaa2ea1b2f8a4cc2edd6b6f83d2e97991ed98c38c5302ac741e062173ead9114f3735cc2411cab26ef1da0e065b7ac91b2b40ddcad368266cf5abde0b4db7a4722c695d992476adb80de25cd862f5ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d369aae6c9a2e33a845498fbbb2709954c5786f3a03ef5f12421cc68f09ea5122b2372c1fa72bea235a32c3ef7c1ef137b9fbeebeb7b5ad9a9c0d14b52886f0e7ec2f03960cd498784f41766cb03264e385b517d62022ff4313aea5a1dff05649fc06fae13161c89bc4fe22375bd48989b8e6ca1a8ab48f38f0d6274432579d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a682259fbac9f0904b0947ddd33807e6866c3d8a92423f67301e2841c32f88ffc5a3185281b553a4fd11a416df7ae6fdcbefff1ed54f7d9c297748f71f373e9c68f3989475c53ba88ec0c1f34f4100db787aaba40343ac922b5f158d0163b548c61094cc3468e3266386b2c9f3d99e6ea0bdcdd5f8144cfc02d5cc4fcc4df18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57ebaa188871b339002860afb0512cef40b3c0c66f1991f6d296b048a5922d2739ab4a2d899e9513a9ca2efbbbcedaaccdb87a64ad638702ec3c00eff6f11638745efa1cc77e75146d30086f188df2a497e34130c985704595dcdef353f40514be90185ecb54c810720500ac3cf8d336c27a05e386e605bf76355b412b2c9ed6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc9b4bf1955f35d79719b52ed153f2cd10921ffb9af1822a14162a1f49460829c7108773c26df26ddc23afb1142b7aff86bc30ea58466e545743660c498e8b6131923e2056be723c0dbd5345961aeec326856a4c70b6c0caae22b9adb03aa99f0fd7d5c3990f756b7f7a1507ca145048572700a6883b573ae3eed5bfa098fe27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33c8612a0b60bc9c64b2105e8a9ff97a712c0150fcafa0ff4668b9acac54243c98f5585815f3948717a86beccb5d1b512fdd3f590370a9ae8f4e02b62ebf213e32c8eb02bac8a71d8998e610af375f466332d4f3c2eba9d62d5d4c47b1962fe8fcea508179c1823e700d171b9058371537d7a9f52d5080b33cf7b2b300866cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbabe84738144c4676ed359dd470c5cc7028787d07d64f2158a581a7449cfd1e82fef05b74896fd0781d97d0c7e15761450b15fa86c57055ea4f72d0ffe8be0a8567657f4cec72ac9e8a78eecdb318381292ed2d183d8c207045c821fe5a4063465e2991142a6844015b4054a2b81ce6dd7d268b5cac88e660808bb1b08ebc69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1695769eae5aaffd9e9ad5eac259f12f58ff71714fd63346a35c081bc111530be85071f7b3496fb263058a6b7f9cbbdcee6f23b4770d297206fdda1401a8722b7336a17981ee1724c5c8fc7b285eedeb15c3b40e9b1aca03844976564b1a06cd94a8e494dcb1dfb6da68d5bf54343f602ed3485f9c8f050aec20c1e52cc06c1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3abcef8ad490250707c77eabe8178de1c670453a3e2e2001416e55b5d5eb2799b9a7f7b0b9edbedacf869db78d09b079cced709e8155f29b6594c9e6a42f4d5f48662213b2ef69902f24f2ded499693f995e81549afed0441c9fec568950689a25759e2f00c48daa6e4d4e9ce09b18a59167aea1281fcf6ba8afedf4f347e0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he45d1858a795636f50d85cf1515351ac89bb41a72836bef129cb55573cb66d46530fc2f00a5da7c2edd057dbf03a278302d14b635c3b2c49c25567854f7397f46fda4bcb117404dc5b76eaaf4da6af1084998b32a7bc11d239b54b552ec1c3b415fc720d3c08127437dcbc210670d3433679ee512a1b0b217cdf32ee4efb42d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fff0cecab0b72a2c0c837ffe3363b215120538379b7581bbd97628cba75558a65db1c36ef0be3307e042b848da66f10e71260aa38bd8d5d0c6d2c782ded5ee6ef197e4142bda46992250f8db3d7b15fc9e3f23f834a2ba2b41f803180e8ef0f7abc2f4ef2814cab95fd7f69b6c7025d5e953746ef226448b6c3a44131335de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d89c15214fe31b57dada3244fd0194f85e253d3633bc46f606407bc5f5f3c9e6394e93826ee4bf7b0290f35c0fed1958b80ba43368e1d7ece31fe433657887b4ac0939c9e32cef9867fa3fcb2b94a09f25d536bdf104be6b003a4783824fc250d259d52983a6fb7f6dd9788d7282d4eec27e01a08a1ca5015f8d5ce1639ab60;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed80e0edd751fa3e7e60830445acd0fd9dea634d1d774cf3a0c31b12c29ad5c3a5c74d90186aa5b83f0036d6dd95c34035babac42d7c1bfdaa8db2413176a89dce50f4543b8a2c2091c1a63d1ac6c9eed4e4ee9900e6cdb0e5eff39d833a0c92d4f848ec2c31f2d2675276596f0ad673ecf0064bafd25ca324e93b043129aab4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22bc206fc8606107e80965179096dc55583c80148900d59911dfcfd7e244e04e82fac28658aaf5a505d638b3595b5ea5168c867e075daf27ea645c519f393b750201833430389f1821e68f0cba835f5ca78683b281f6baef59da4da8f670c857740b57d23d7585ccfc039096b38448f40b71e71604007aea0278876e9c0fb71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6ff664e551cb8fed9dfa3a494944c9093d6a0cf530cddd0ae52cbda06549e54461b625b81f9768fd9f8094481c5deae1e81fdf9cd4ad5012765a72a29ca87cfebbc4c3e59a0ee1e682803f07918cf10cd8034d78a02ff0c6880a804e8a45303e9b82a6e352e2ccaa4487a70cde95caf36eb5039603dd23a477c67935e5c516b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ecc0f61e407451e98be567d173822f30b0ae9377db5af07ea67a8aa47377e0271e9939f5ebbf6cdf6c6a51166f9924a5ebbba7c536f38b40f526f3aff529f202d784c0e92c15c1b7a40a1b6c6b4111a2ffabb3d53c9a58a769cf75b96a94922ed19afb8fe489afd695da1fef8b37a93ca73549e11376366157b4b4aa35471b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7922eae6c7d985e0800fea9c0873c4e6efa68ac356a6adb0d958b265d33d0920f0ee46101ba586beba9b73b070831cbfaae58e1d6b2350da94d5d2619105a1557998915295e345ae1aa8277d51ab084160067c6c5bcf9f8a8671f598ea87a60558c55f09a2ae13ab6496d083ee1b73dd4484d69ffad7d29cc711b3581c81185;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haaf47d3af4fac0532b14eda1337b7dd23472bf3c49bf66b8a5da2ac8ab70e1a71f4632521b154484c99259549195c4fcf108fb2c2aa40f4a5b3546cbe4d45dc493c94c9f352b683d843e8b74300fab678302de1c6204fdbdf82be22bc6c23a395a33699948c5088028a7e376331e4aeffbed6edf9b0e725320de05a17e2d4a6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b35099d523181a2b88a6f5d9c219ad8b2f7a9877a6068236dee64adb21e5d42346f27628167cce921425a469a7195ef53e78486cb8316ca58808a8f6b857485d067b893520a699af261dd45314ae6729eacc61656c71e73c8406f1de79e108be2d3a77846ca2d0121e38d12e95479b5efc0c028d3819d19f7300bc9689e59b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63777d8633ee4b5fd0707b8d5c696bd541f576fbc374f5025ea7adf455aaa69431469bf0ebcf840fd0cf13545924b485abf7002b7e05b99d29e83afc36ac91a8473eda28cc7fdf758b949edbf79d53d5333fd68d1cdb8f581acc1f4d136810342c7f20fca3363feb03e36c7f71f21e0721ea17d2d7027e74fed1ff94a745189c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h256c6481d07373f9edc4ce40d98888367418ff97d5f6099d3842a12d38118ee10dd079474bcc374d8bc9763c7db18cbaabee6b1db9e392d0436823f80ef402f38ce7ee4bd3e4a84e872ca01e12b255902ae4e7fa9e9e7c487826554aad13573893d026dc2017737c263384ce7080ddecc055f87de94401ec7812c8e3c34fd12f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bfb21ffb9548c1cfc9a37db3c3e42f1e2090ff21da02319713da6fd6f1907cdc4140220bd9820925fd5b19e5b859bb9c141c9798fc4ebb136ab5b3d8e88c5dd48d2773933d311094623aad9f0b16d25ebd958591d985b5cebae56adaef8cf85236a3bb4d7dadfc7947f639016a97b75baa617a30a78bbb2e370578dfe74ed9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bce435b75fb7f549eb463d3d50000269872ef24a62b2c8e10d8a895c7e5cbe60735871e9c9c6f706efa298eb17e86230796d32ffa95821b67b2a516f89171e86ec7d00b544d65cfc989275c2917a2fbab5771749a95c7aeace08f9d62c9d2e1541b18c9510ea48f1b736a6f6c3c02c1fbb0061d8bf268db3b16ffbb330139d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59af8a826b2bb01b5628309c3a78ae5ce89995bc5f4853e2384b053b7ec0db7b5ec8ec98a35720f1c7197bc3ac6c6700a2556b5abf3c4b4fa08dbf8dbd69bda9b29a75c1973258a76a333cd8e851269408a68cdb7e6f639881e00409e93407fd8ed47b3670e60edcec6885aa979791258eed0d5860c97c2c59056fab0f74d93a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ec47d9cad7ff20cd0d4e08ceeb13fd755355f038e8366f397606008cd4b0385e3b6a5cc5ee2f310dd634fa5372f7a90c24d7dd7df939d9728e59ba36e94b41af37265289d4b972011dcb2bc368ddcf59af83ddbd6f8d6d7946aa4420d94bba6480381d45b6494882123f23af7a531d6a4d51e2780e3bafee8ac79114e8424c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa91daac9fad18e6cb0ea3e327d9b1e4a1ee8b3bf4c9430ac15da86427104624f5503ee455921d36589ad379b8d90869fc7c9df920886593db88d9bbf1e396d987dc686508d06b3ddc24795bf17ff221401e5684cd61846045387988efa1caea23fe829fbab8bbe82f7fe51a917d57d07458a270a2d41590ff16a2c1a5e4fe8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e3a2a7970fe5b7cde69995aeda29f3349c77cbd250e530709cb5efd55b7bbfe063d10955650b213a9e7f08b35fd540ad480d434fc48d4ab77889cddc863e03a354bb5e971922c82ea7939da37d2d93024046379b04733a6e566ff75a79a85a0ffbb19156ff6d8bc6cde00e0214f286fad6ed320b5efbdb3f0a58927bc2f7ac4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb23fb421a67cddd9d9182cf1d0fcad517dee291eb3fb59215000e6a8599601d09c75169e95b9b9302fb17bb182879e7732ecd9d29f7518b8c5241e65fecdacc391e7f33dd1af8fd44705c75beac7fed1b20f8c6b2b158d79ac1ee3836a78ba30bbec4090dfef5d749fb6eb1d2d6cc9ae912b631b8aeaf5ef337d559974505366;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cbb0979372bad6fbdd42bcac8975ee0dbb20cad3ee4dca4691195202c4780987bfe6bdb47c7c3b7dcbc69c8b47a2137d320e7946f4f37018ec550f4e463e96856b73a32dd08fe3f26e0fe3901016b4ab641b0ed161eadd89f1224bbdd018bf5d32177cca6cd5ff4cbfba7e9802467061ed326907ac30fdffdf892df19c197f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h175aada24d2b070c2e7bbf57ad4b975091bd1b44f16bf0db135805796e8beef97841c50997b7dc34ee5dc22525bff206239a63aa9e820db7664b1e40ce24781fd968dd546c6f4a6134629de9ab4da63f3068edd6bdbd8c80047037ad4078f4a7b044285e5d52b8c46ab2537cc758dfaa2335feefee68ad9da343793de41269e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ef4bed58bb210cf778453ae514d4457f793283f75686835755d8fdc30e87ec20345bf40830803e880fefa420e8e7ef39169f06a4d0500639839cdd8b739775023e23dd8cf028c47a091d1b793d578b32e1a955d638930c541beeaa063b80d3b76439d32b8d018378ed5c22ea51df87d085d7260db64a112974ff4aaec204561;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a0eaaf8ba98a8a3ee733b3c172d46e8c6d2fd930dd72a3db34964cac15b88174bec32d6d616fc9b74b9c3e95fd18e9df8305760ade507d27a5c3975cddd8e6229d662ea3fde05d4fffb667ad3b320c08f2ebebd0acd849df7f7726f43a478ceeef10f603692095a35125e038e70e644357871a8815e81b97cfeb3b6020a48f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h926ff89e39015f5ff46095129c0f03726db03379d789d03f9f84c10055a950dab3371ebf5a0f9a2079197006a0067a2666eaeae3f770b3820a58b3fd6db98254a9d909878227f2e472e41eb349732669398156d3da6a4824f0b2b3231032d8586e481f76305f753ae3dbe6c8eb752e4a8b5322539a79b85af18644b275a87929;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h420161d46637a1d35e54eb6ee102910b5b8db5c65d5264617f1f3060a1f243f0b401305f1b509b33695b04685057399d3a6b6232ed37c712c6704e45e2829f14c58e142cb4ce7c8085c16073f45877a7a0f4a8cf7cb3ef080d5dea5f2891a0e60eddfa9e4550090eac09d566a1fa7bdf46ac93786608dac23a73287406bca32c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he799bb020ddf888acf310cb5db068d4d96f298c44df4176b04eb1014e88afaa0892c414d6b4ae157b1aa5b693abd11052314f9f65ac66fbcba23b2be6af1ca73281259c0b4b80d1cfa9f603172cab39b21fb698c56f8971fae8c0a41b4f4ca6e22a1e87022c64f7b6a33ba0f5e4ab10dc12e9a8b73b9e82f294016004e90b710;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hceb8d067571df9d94a2ffc5e34c0fd3c8fcd25e6e562121f5c466061656d5b19220a8611112e5a57a891aa17b1c0e61714a3e3a687c2d6cd28cf586f0d584bc77aae120be95191b486b01b4a3dae00e179f133dbf0137248f67140fb88029709ec226a244112c6f45d2b55ecc9c6aec51dc32abda2b67bb198320584ecfb7df8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haec01f03a18bb8bd3ce286a24c6504a65175dd9bb5cdb8537d593e0d6274701b25fa0deb706b1d9471496d950d119793bd38c357791ea5b04093df6d99d47134321f58566d03bb7335c855446600fa6ff1ba81a9f5016f2372886b128957f101b7186f2317137e64a3d6402bd87c04168ec7ef61f015cae89cd1f5771896c6a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1861ec3318ade758b9eeb17652ff8fa4591ed5658f6e7eeb26f56e4e3a1831b0b4e463d72e9dd17fd256a063d979bf650dac59066baa67f37791a0dbd86aa70f36713a65dc184602fe646d0f10505b6c5ba6cc0330289ff05e78c7ca001ec8cc8694d13172d8e99503bc1fab03e3bf1dd6d572f36b229f867b2b1d5dbaa2aa0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc16ca014fd22d253c1dfbc692c1005ea29556d66610f2d54884dc8b84c1bbdbd7b9481ef99631828db7ca3ec73e49ae112e96af4916ed13849e83d5e6f29ee8b504af7d55bf85c480d2514a0522c84b535c7315e5b3f73ab27ce4de1368e8df396fb79710df8fa48fa005a20cc91ada0c0820a4492c2d7fda96ed0a0697e15b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9190ea48619e0c3e16c457555e6cd7f36c98bfe05392af278b4f7dbda28a8516cd9fecc723e29089ac2814c65b7ab7c580ca9691eb1006508f890cb8afb6e6fcc8ef0117a1142b341c2798b40499311716f53ca8c28668c48dde07f0c562d7faf3aaa529ea70d5b2e9d154ec30b04f4f9c591bf4c63d3a9e7d938206143e3e9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78a885a91628e3c3e276f8104ac6ac28011cf0438bec75e46287087c81e966022731c1cd6dd923dbefa29d50f6279cce7aafec2bda9597e9626b079e08c101a235b52912408fc834dad4a506dc1d4adb1bdd10200217698224593ab1ea3d83ee15487ec02d41dd626225b677d233cf3f706f07c735f22861c12cabf8ae961896;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6faf26cace6d5d9c8f6c2b4306bafe52806b830bf6f9476e91cca4131db042f6be9a1bd1e4498222f4afc6860026641b167517f6ba4f89aee7a1e80e3c0c03cc506dff99ab3c671dec407146d917e71bb0be2fd1bc647f69904ef7f4727a69d9b09bf72a9abf3d6228f3183941a973f4c2eff3c8c97821fc194b49fee278ed45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bdb8c077a340dc26b136fea99b845676dbd6d461e43fd3f9e0a85b2deb5ad51bf74b242cfc030359f743c5a172cc23c516e2735893a0dd00bc026d74921908201afb9f639e964d9716d68f3fb8ad6e34b3c809e55837c27bc7c7cedb50f798746f37b9264ff812a49cd9550eb276649439b2ae913a7ca76dd8daae6cee17cd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habed3525b5db473b90adf6a30b2719f10bb1eccfb5791c7f3939f4c1ee90f63fb636dd852f005d5684abbc585121d134d3fd6a1d4d3f07ffb5350ce2b7cfd358acedcc2247b26f21646c122ac5af5249b24960ca1fd8afaac283d9443724e9b31a4d1d48a473ba96ad90aed350ce9078c06803cb9ba3bd5a7bc712483452f207;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fd7ce4d14f55cb3bbf7de0f741c4b985b5dc1ba50adf94374b08a9a496c4c4de8cc27a68d5a33b64e17257c5bbf331ccfb2577d9b31117aa310b4e0e7e07265c50a7cedab7a54c33c5acbcba2325247608c54c595ba603498f2a5a4042de276aad021dff8183ee31d1ec2cf4f7756dddb97cc8a1b881b4a09ef8c93f5f1ff62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b36f374cc9bc9575c7a3bd5c7b7fa1a8df3fe9b3fda3ba559bcc9f2e3f8ed5ca0c335df61018d94e66e6669f2f01a8506f09241c306388c881cfcc5c1600cefb135e451c09d6eb18a39a38f8ca047ffebfd89ec493c01ea2f9d410775bf069089d6044bc5ece2966b7b5ea11338ad2f66be78597564d8be0b965eba34a0701a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ac7f2cdd180ec89f65a6295eba049bd5c272d7ecaaf2aaf0240d93bc88ac68b434222ed574f6eaf810fff74197bf91dddbbad838afac9865d8ff42309a183f79f15192578bb14fedf3363c2460f920b4ab0c4af4d9f3d0090a8776a195e8ce80a3474d3b94cd5a9dcce82251dd2013c49897c76464cbc0f210298de1f99f96c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9042480597e4571d6b3ffef1e69ccbdd5db40f1241834a9f9935d7e3d09cfad40f9f2042ad543d0bd799363e6e8d97aa11c5a9fbb6602437edc0c2efcbae19ccd398d332301268731c842f670c8b7b2f60587f063b9929dd6300bf1303df12d81f190598004df243d65ba88f4048c0ccfd44813ac037b091610a4b91f363c8f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48234990e42a20d579df79981b4896aa7d2b78be03146647fdf6b06a170fab32c6b46bbe1079a10505958fc4b25dc927ab182e26857342f16f82d3a8979287fe870345b592cb3344be807860b30485839812701eac83730f5e9330c253b1fa355076908157286ed81d6aade7b8cd320bdf5fd84c6bf07dc39ccd35fb88dacde3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1995d44377c4999f510cd7393243f8bc6a9c024e35b728da4f549915794c45e74e9d8640e8e99e340c146caa495b043c2985de7c861eba9331170f9d207d9bc22e8dcf1aebf6e5c0b404f4a19b57ca12796b37af6cf10c213f48a849bd4c939e6836d7c4572cdabb2abfd96a231eeba03d1baea2db73702344e5acab1810e42e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha27e0974763d55c0863863989d838ac53c61451f5021a42f7003d5d7f4930984856dfd107b7854d4c3649c61a5880c7fcd53788a6eb005e7023f940d0c5f727e641a2b9c16fb571aa53b25b3cbcb107e6dbdf6231a41ea3573341a2f5c860412ba458671245f47ce9e6c840f20b3433c465cd4d54318c50d187b78679b70fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7aab8836a98f1fe0a5b4364358d147717c96210eed3f6a05bbe9b96970fbcc82831eace688b520bc773a082f099a783375a8c0be72be45a246dc5a6e408c28fb3d9217f161535f1b824cd3467611e44e9e5c04d95ae2cfc444ebb4f52747bf7c46384f4dd5398c47ccd0a7b833cb88fc8f1bd4bfe7b8ef612f238279bcc38055;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd846864adcd994babfd1b157eaac3f6f04bc5028968f54c4724f08dc4017a17ddf8eb8387ffcc95f4128318d38755fadc12e04933909a98a05e717a5300823d9b2ce228003dae17947f9cebd893189e88436b37307eb26c7a012a91968cc04c02f5f1b963cd90734b7b1995824baea40f4faa53bc4c5db7aac137b3c39bfcc01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe15babbe736c84694e50a6a0f0adf2c5059d51fae01060def83e03760aa67e0fb119219cacc18040d7b67df5212eeb3d157f3fe40a822cbc69da37a93a9908698cdcdef3fcc75ec28e8d3b8414b4804017ba29584fea977bf6b7e68db6537ffe279042329eba52bab06aac229e3e5621395f21a7514bd7e5a4055910f7fb018;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc612b581b817f1a7f734d75d2db068af30ecf7f20dc1df020fe8fc0c35168f95a0fdefb811aac220091f2bc9e86803ba32daeea17357a0b03e493d2425578b010e0e9cfdf6d1776ce9cbefa783de7c939db851d4d252be3b44c05f714a62c5abc259f647c530781b0b4a7b5af4f6a74856c87fa74fdb8ca31de8b0ead3beb5d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9c98e8002925123f66cc1a9fddb4b4ec360a38a0c2fc3253d5aae14c1708d1a65f34a32c60241f822e8b194714a3aa30f4b0e35be58568ffa55f9287da47ff1a39eeabfd3edcc3220f7db57dd1bb55ac1e4a0cd9eeb70ccbc14dc155b7b5a9ac856f707addb17bfe6387ebe065f135f511d137ca53c5a29825a1a298c0ffb8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b1eeca6febac662f83480a0ebd5a30939043166f184899cabb0fbb8e929249244b261203164d30be76ad1718b059fe4492af51e054bcdfd507e95a9248c302c3a312e748b188fa5becf7a7746ea017d293429cc914b13d5694844f1cfb2587cb4bf40dabeff897bf74085628bc322052742be976ce89deb55f8c60bc4a6a77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87ca8ea0c799fb5f1961a1bc8e0c2a52bc252afdfc7f65b60df1610411b3006523b531fb48d6ba25aa3ff3aecd8f29a1b32d544aadd8a1dce0fcc1f45a4f045cd03e26641a04dc2915399d0dfe93b3dbf507952604831fca75ca3ae7200b2d794613f5dee53d3731edc110b12522621e7e3d394b919bbdf7d66c822f01dfd0fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h804bdef869dfe691af0f151de9658b43e01a8fa452be9045e47204c68994cdcbf1ae87bcad14311a406f40542b9fd9db289eca078ee5fd64392076b076361f4763dfb3957db20aba8351f143eb2c580bb9d882773b8759c89296080970361560eaeb4278c16adff3916e1a6824935749b49b80a06518458837b50d8cda877cec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31b36fe63dc09a2c8893c323c82530e692e6f1d802c46d2ce68de917c8d4b248a0017827a157832f0f9464b0a36a5c69e176790d5060dce53b4bdee80ff254445541b0cf2c80c22c4b57bf62e538f6b2725ae2dad1d97cc7d7402d6fed2c0a22156be60c0edab17029bfcdebfd461ab75fb23bdbed4155f89a0d6a4ed82718c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5474513ae15389cffdab39018bf46e08564bc2b6f889b75802ea15157cef8827b358ec58d15488ce5798970e911b37cdc895e56c7b3cc56a7e1e340d62df99390938bc9b93083d1e4a1560cace5104b056a4630724f5a61261ce12cf3f1e9b4a4ed6aa25e700178edf17b4ace90dfe8ee41a57286819f2037837c9ecac5aba30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb518a3aea43a847355a7517e699a67bed188806794aae90e108968e427e68ceb5589168e83401014d2ca3f875e7b962451a6d4fa03de7dabd39938d1f27fcb56c66b2c1ae85e1eb300d00cd1f21d4430f755355fb4d5b2bd613529d8fa040bfc79d47281bc9cd4033d6be8f90ecfebc95cc03d91bef596079eebbe2d2541ea8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a2aff4e36145a6995e9de76c5bbb6d96d069f6db1157f7a92bb1941e32f6b7354ca508c4ab2e451376a7754f3112d57caeb1ee3719f014dde4f9fd27d4c6acc7c534cbe13c4ada7f3aa7a71db24b3c0f418ffdc2eae5974affcd6834cc53d1bfa11d080d96080ab1f835f01c2f2353846e0486a990cee657ad0a5b53d14ed89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf03f307ff31e18b29a7f7f647aff99583e9c12df392930b893e2e2511c8cdd91c1cea0c1965bff60f05eefbccec6beb58af6bbc069c04ba700b64e074bd759215d5060eb3c4dddd948636d8618949b82ba3cf4791186ec17d8039b7257fd0c17a29520a16cb4c522a9d92f8a369fa9e8136d60eb715f591591673d4a502cd49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8876243b62889f79ea195526b431c9224140bc62953f0e52f9db46be7fb1ab393d39c26397c222f510575fc492cad49f75c3db47ebaa9029075c3bf6fba67b41c14b49d62f451194ca7263c252c48eaa16713069d6a94865339dfb2d3d836127ab15539baac410e0ce96347a2accc69a8903d8d5f8edf865376c03972d4bde3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcedcb41198d7ce1ca769b4e1b3c530a288dcc6a26483b479ce28e4ad8163754099ea73df17706a8ec60c8c55d86bf902f5197b06ca5e8176ed063b5d558c310b019a3f6a6214d14842001c94c10fa4cd12b7f495c2b6342790f650828e4a55c54fb8f94e48040e94bc11f3e20d402e63ec704b54d10ef024c75343d88349b639;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bc7d2f918b63fd354a71b8a33de3fe38d53d178dd9201ae4837452ef95c13837b2fe44b751766860ec6c12c076f36e66ae8ad7ec679fea06ce46c963482bf325d1d94c5acb3c2b26d4784009546a5bc9d4f5ef0ccd16ecd7efa07128525215f2f8bbfd8cf17d07d3033c499f8c3ade48979b9af7ad761901c8f0dc733566d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf047bd102bb1055f48ebd2e945cfd7fe980addd303f9285e4ae15148cc85c9ba698342d14d4fb01f7230e4333b843840d3dfd313b6562d4181896c3965eefd53318ae666c2ba70667da35c18aaba7ac2de12a7779d99eeff78ec904095df2ffcb0e5c0f84bcdc8b774547fd200ed575150f892bd922f6be100123529b319d686;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e50b48776247436c478cbba98f6103a91b308521881b1641ae789bf8e41a8bba4aa009da57c6f279fe4fefb421bd60ebfabef8f69f087ef601ae02b087a80bf76e1bf1c49219ad003ab03dfbadc870f58a6607e0b281fc2929253214aa9877ecc4493e408276bfc5ab60df243517e6883619f18408cd7e76b9ded20a8f6411d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfd8bdc8be35072f6cc628cbc224aaf97cd79bba839af49a89c815bbb272b52e1164ca7fc9063a0c335ba38476bd3fba5ee84e5de9b50537e5b1006a665e6b6e9a220981667712e0e82a16330ad56b3319c2ddc0ee1cb71e01eef08ef6b952df2ecf1678980d957cfc29c87607044ca2fb4532dccf4260b3ebdb23b09691bdf5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2fabc3c15a1fc11c9fc95e6bcc81134f71de8d3c188a9aa2d93902286594947f48114286f1256a056c27a87a2b0dfc2343aaa1e72746f1b60b90de3db2f7de2c9670f8aa7a57883f90ee2d59a68f9edc021d7dd6c8ec29027fa9ccb190816b889650a58b1ba74909274e74788b5945b6ab49ca3e0c94ae183b90e2ed51df462;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a63c6bb05c89b8c583ee9490161ad678dc9272a7c713d663b62f3b639ef2ed3fa2323c582c10da33a94533e2ef2ffad2cd612e7776045aae8072af36dec46ca07a2344667150896ef76417c0e4d0c7e7a13cb57084574532c36ba5e09f6df98ba4d0f370debd16e2809afb8b5574604df57fd5264c858431ae9dead2ddf1e07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h205772f6135fe29edb47559c18d5e6d12a35e80655a6163f56d684143f88894c30e8695214156c3894cb8be749a25512cdf1ff157a40e43a2f07dc2426e5c8929fc4e9425ef0ec01e8280ba65c4fb4a4edd01b2b9e24130fa2749ee9060170ec3715b5f5a429305d9634e1e00ca1e8b2c765ccf85678d31d737d651435c42cb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3143b43e453fcbcc583b63489aa42aa3b9a9bc1f62821532647bdc855fd83e1496f37a33635abe8274048936c8b520bc23cf5493fea5e9a9c15cc6f6a1b1aa04e78a7308a97560742c35da03f1a46f205dac4cd37d2cb768df3739002d43b74c8d9828ca5ddc12549abb6eb8bbee1386ee6568e05f74ac440b8c106b937da925;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4807f964cf99adfa55c6d5edf3a00578cb49badb94e0f130976e88eb1f0f9eb6e7b96b13fe7b364ef5f6a782f544f4657a78850e880bba24881e9eb12bad07664ef5e982b23527194f007d220e50f37b118f6ea52d83f27ef57a00be21df804885071e0a19e6a022ffcf98f79bbe03d8d789432dc38d8614db974e6df211628;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97ac39e86ed390d1994fe341f00f84d27daa664bf5521aceca67fb46b6772f6d3c2baa7c701d5eb19a59762cbee76b7d05ed3e368ae3facb96a125cb207732524c059a532bb0cbed9f56b6e994d1024affd9ff582ce9be8f49e19b523f5fd984b221604a5dee3f020f5f9049c2ef7c47f35b929739ea5f3d884518242baf91f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h793c35ba79cf30e538d459526f208d84c26d8340237e28167aadd159569ffe7082ab3553b746feb3d5b776c5f98bfe2c088b22cf48713537fa239e8d5c99297fce2012abe933c5211b7d8d7c7270bec98f23fee3dedbbe7e9e2f77a93de36805a1e0c08d216552f5850afde66823ff9f5ab502ca46196849ad78039a5dd6eb8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d894f5b65da0df2c1bf1751f74cab3fcec51de831836ff8bb8301d0c419b312f584294497c7a5ad0db1de40b155948e8986959378c52fe80ed388814318a1fa0b585153e600df1953de05a4658f5cce47dec5408ac40d3434dab3ac62b29d7626fcf053da895d9d97225ea056c756e014bf81aebdccadddd8d6b833418dc02b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc3aa5e218da9620d14ed2deac9135203fe6e1f37a2ae88cb03b0f4132524b6f6b1b10f9e94572f016bd1885a7ffc58aa908dfc007a34a9fe9e803d106bdb0fdc3f695a000151102418d1a98005d2ae922c1aa9d62159413830a1bf6b803d1dd134d9853af07d202a9147f28453aa60d85a1dfcc76b9d20e3177ba74cb7e150c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5a3ffd8e158150372d7cf0ea3ea89c8f6dd3d8c62916b9dee773b023a58afb072b363d9f338af4f3ff7323f9b24480af0602e51628ad4973d1604fe2fd6a76780e2d751b55d4afb8077b341a55a0833d647e59193e2702c681990f9836ece6fcd02438f3e012806a11e92c1e89bb52ab91fe5583d5347f8fdbc807c1ff3394;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9172b9625d173ab692e51ff3767f57a8e32ce1bd4fab15e45d6b3761e5d4d13c7d4fa60d913c051fe075190c9266534c7d610f51f5b11205f05a195424fa44cd35eb4ebea6451a72194f6f23a3ef891e6466f83f83778dd48ca6c7fd76d7eea9bc9f1c8724d3299b3b1ec09cbff04e5267c787e5fda92af606c90f7f22411156;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ad989eec5fb9bd55a8a3280e3938c7bb396287b4109f572cc1b7591c37bd468f5a860968a0689d464d735b643c9b00c316549f53d92edc62c13b33dc052eb70112aebbcd72d84fa2ff2252373a386bf4f9cce85d39470386e43397d88ae9e9c9f036782d34f5c1775f5e5f10146d7dd62eaf7a696af6a0041be30686c2f98b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed4ee9e0a7a4ed3f07f8cef01eff57d60e7684e928fe3f9ff33d21286ec96ba01a99abc9abc18402c9713624e615c62a3c99faff6dec74da901e8669782aac37a90272e2f345471fbc887739c47de2d507410293245c31302e84344aee50cfdcf71c21c31ff0f5828a7ae08a406bd87523526d8655d0d5f4fcdb014f4780b202;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h226273d0fd50aa6bd07dc75d344fdcb451ab2ce59610cb135fcfec5fad1ca8023e6e27680ab55088ed17cea795de72a03eb4090e2231f0026b9ff9dccb633a302b2c11ffea4c9566ca48a56291e8e1dc2a5722c8b7222eb56cf5d6d2589afe91c5dbf5bfad8368e3f02e4bac00ce1299d3a40218d998efa250b2544897e6d51a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6933f6c211c4d53da4f1de04d4f149ad30ca475299043f32bfb255e226ff0c8d64a5fb92829c5026e2f28883e329888b9d60c143e692c2471c4a750c6aab96918ade36ec288284a9d0ba4cf849d2d6b2959da4b5afcd42dcfebb317b8d68ed9fb67ddb13cef4e3814f18645e4975c4207b9d65e994e3febe8ae79dbbe1d2f72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac38d3e093c3eaa27ef5de630534bb23615da5cef3b6fffd8d467433f385951f32c95cfc505c866a12fff307d1fc6db14d50c1938ff2d13bbc9f8779051b32daf81740068d9ac4741784d060392dac81e3d99260884a46aa686be412f211bda525311df9577a13d03cd1a1cc5ce57467cf71e57fd0b9a1df948771e2c509a8f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe6050d674f0b117046af33c77b3040e229023ac3c51c6bed3c19348317cf62af2f7b3195181e19f920a12970addd4fec7e1ffbe2230f31a9748dea8bfd4aa2b59203f1c881426a4c92590974645bc144d0768842080b82db0da15d6b5f9f5e345252cde61ef621dfb5b8d0f22d28a893057ff20379f1c617ca9124a9d99c2ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc710a7acacad9b8fc4d9a3a3dbac0ee03fe1bf14484e63dbc258cb804ed6104e494806fbcf2d694b1d68cf2e28ab24abd9877585d5a922c4e7935ba9456bef0b20a100beac44404c7ff8f2a16be8f86fbf6ead3062c6ce58e4bbac8ac22a1b456db81d8b9c6c38bda229e2eb5e9583749eaf5c7355cb287db3de3e1a1c3e4f98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd388ad04863b32ee5a6341d6097ab09de5507286c7c43b8923b0c8268d4821bcef835eb80069e91a22b5dd8b6133743b41b9861b4dfcced7e838ca11ed8666d90acf58afe93b59619f013d0352c24b41a1dd124fb4dbead0469dd6b551fdb57768e41d6618dbd621abf7dc2bcf4f1a0ee95a62657e8c12915e4efdf646bf9089;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h345d1cf3547c352fc8ec51426bcb1c781d5c026daba8b0183736ade489464e136a1eb1b58d37029e87ba004e2f1990a47adb4889ecec9f5eeb0b4894d9df88e48fc0f067fbcf9b8d0be78d74acaa5f1b4929be47fe51bf183118629bde91720e3988178235e193cd2e3d4ca6c239eee9eb529b5b3c231a5cf22af01d35bd6e8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7137ff9cd474692c2bb3de77bae1d5c7122809b640435625b163b88fc450ad6149be4db6f392d8703096d0c61a1213d554bcf1f2ed50a1af12df272d52ba03f16aae2a120ac55b43595c1f1c4f0e57af41c21f6cc6ffcfaa72dfebc8a0edada336bcf9b75f3f30d4a0882c1a37e5d02321faf99a3659a339da88069f3673323b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3900c109c5f9b86e3d6eff998c1982b8e7992c6cdeddab91b3f89bbaf2c4e7480c72fbf5ceec82c9420ccfdceb9c938f35f6bf62fea463b7ce532a3fd8757e5627483e738741f0b4a8a4e949ef4202bf3e0394bc4a48adc4fc83125aa57b24e63db1c69f7219c6faf1de150f0e7f91a062c9297ec4b57c4a87f03093ca62b2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdc94b591689765177627aafdcca474ab3c7f27c029a6d9725548151b7a0ca6cca4870f8d2fefbef64a044b571a6c0495bb351bb6891604e23e1560d0e12c0faf714b5f7bf37b4fb3f249dd848f1d8dfcbf3301190712ed02ee6e449dbce2c8d18456782c531d08baeace370a02d85167ee1a9fcd9f779f0b947ec3fa8bfb438;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c791436cc71cfe983184f5a7b85705dd5b28fab9432c90a8cbff5d879f1db13d59ff8b657a1590b8deb02c3c9041782c2246c297efd268002643f04a385aac664449d4980fd954c3bfb44916b6c06dcf0ed2f4fc0be64d32033a20c733294f5e6644446d78dd7c42b644f0692366cf0709daa15b73c3c5e933abd981d32e7ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafb122143b38bd2693b89fc7f892525e4fbf6a3fc27af97a567be1aa00cb5dea4961ea1cb0c0d743e94bef25cccdcda87169189f747506745158a996e9cc84c028742b7072b194cd14f914be02ee638ffb85f50ebcb99195897c658cf573b8dd79c86197a62879fd55090df7614ab60d0ceb37fb615e906a6544d7698135de01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1200ebf76305df89e29c39014081d213048767b09e7779a463526b17e8e35efbc54af99a2d5b5d176d8d06e220701e64eea8e22a5d0bc97129f6d99f8b20c2a3274d334629d05a876c6937da9ede26d61b45e5bc73b714f7116a0e4c003867b0651b9836cd2c2ae240968c9259ad8c980c48018a361341a38990933437499448;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1fb1ee228bebc0eedc36542d319b04e2cd8ee10f06151106389450073e4b9b9a7429999fbc039d3a95a792ebc33d17be0d82b207086e5e29590999fbb9861753448225b44658eed23607bf641f325642c87ebd2c26801330aa65d3dde9b7da572679e51b5b15b425a0779df8e24265fb9af1039c5b8a07f52c5c2b77edefe73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf9d0c78feeb6393ed4d2f31222a3b4e18024aca923600d0d9f5b01d0545deea69c74ac4e5128df4723980fa868e7c2a81a8125af17517971d385b7e36b66b6e2e54b8868f3e7894c2928dcecbeb5abf97aaaf092b14ae55e37e1fb403866020bebb5853bc55b024b03068fcdd119e14baf1e1b5f11961c34e8d10f3fe1a007e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0458148db5e5902542b006281a43468b526f3aff77f9224c56761390c69fe76f3165080ea9e3021e31a8be128b7e79598ec19e579d01ae13c656babe9b124583eac29cf78883d5d7aad4317201235c52b50173b523f1b2dbff2728d2ef63333ed2648ec86c4bbccdd2acb00673d409f6046a22112769848bdb4ff8c0e5b5e6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7ca6265e311403ebed3384892ceb336b8efa217a9b889c911bacf4ec913bc59aecf924f2e7292fa145272a02a71d3ede83298a167f3e5c5149b88491e6bc29ab29c2110498e7ad0c4bd73e84bc104229f2d6578b0ede6a5ecab39d11b6a9f9b983da0e027aa3fa605cc1eeb14e9beb803f051fc8570f807565fcb883861a851;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he57cabef575e449005934eedffa757b35aaeeea1f09d469e91c2d2a54a8fdd1c49c2f0f44ef0aba1f9c7675800ba7b57ac171f1101bf3f3568b962c0cebc8d4c09c1806a573a65d5f2082de98be547c3a55ef178872cf3dc74818a26b2a88c8fd52a09e382807f5d6b50aa6007c49b6c5e361c98fbdfac9ac88034089f355f61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf61ac43291ea235cddd091536cd1ab7a899ea892c1f672e400eb1fefd98956a6257a4561a4a3ab2be263d988a0ff8dcf845bd568dcffb52f8c291bb942803b63affde7998c9a951fe0ba47d8df0f9adfa1400f113850357a96dafa7e9f4692e8b8c5940e8a2de7293b8aa98867eb331fcf8ef30b460c225b349764ed5bfbae8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84667c5b1bb93171ff814483460e456ff0d1a80e84bed2da0bca7558b44d72f85ca9b130456a936c1f6f3406d64fa061ddb080218174b7176a1c4abc5e1fe9c5210711ef2e90bafbc2afda12c2906b117aa2d263de2c6cf87e82cd134723707ff7a45505f1d37d8f0795431d4c3abef590cc9afb151356e63aff77c0637ab247;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b8b331c55321030b1a8479f7b87b0f5f3d897f3a762b7f9ffec320225f6fa210f2b0aa49bf0f7b5f63b12c0f0d8834ef3d870c7623129257904edc56e0e6bfc0c2eca3dca9246c1937aa7466a09904c1fd7d0055b80ffd673962ffa1170e790b326e3be4851ebd9158b509effef174df2d288b62f3aecc8e75fca9c54b1f005;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2db681dbcb4a0f961baf9715bba8755a396135a64a2509b65db0149b753a0d55fbcbe8d82b835f67ac4a360f0eed1425628cf494bd42c5d50e60c7ea280b6dcf67a369b0c5e68447c726566bd5fe939c3a419e946607bdcb670250433e0de8ee923b1bcaad570ae979cebd4612ea96e7a5caa4071fa4f500849fd4af49af7503;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cdaa483efa4ad17ab39285002e218c6129344fe30f262e1de6d301593ae29343e17db894c6dfe1e22534f015ed75162ffa140201bdcbd971b88ef5c3c99d6b0490fab86c4d0bf3c9c7075c5f019e3469afdd82bdb302061ae155dc4c359d7f487b699e66dfa797f9145ed9b38e6f74c0f12a97d03a2cd8f5bd5cef6cf0d1271;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5b9b37694169742194ef9d7fb758995835762da5c315c44647e71b38228add02f1c5282016aceb9cb8465a7aa091bf9de99ec84807f77c7a9e831be5bed8e85d97db3483179f06914d7f030380415276c6e48b829c3236ad5aae72bd68215fb85f81ef901e8c5fb8a41a725d4db0e394dc903fe6492f0e486e00da816ea8e6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55284d1cb97c76cb25ba09da339c327c5fb6b6891e7179813385416c8f44364e49adedbf2611aedc42434f7ff749a6336d123f1e54263f23d9a7dac31e38fc88dae962fcaf69288735805d72e510ec8196fec40f30106bd21b9938df7dc778b163bbd65573543c7919ff8cc40b1c2d97239a8a7dd61f5a346290ef261de895fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5d3221c9413ef46c54957d85d8b7bc663ec077e1888b0fa4b00c52fb53c9bcbbe2f3386d540fd64422aa11bffe8bb4e4d939b27c5dd7b5e8a401617c1734d51618658905d5ae526d437d7f80261ed5b11af55577e998a339cebd78b58f6e40330545313db028a326ae4292d849e49fd6b07490ea77241cc1998c54831e8203c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20b8243055827ce73aeffb018c18bbb7f6ec9348a8c4efd2fc487a741dd9a2a356704323c1ebac8097282c3d6252b656e7de9da89ae768ad28ff4bd946bdecb5f771570cf883b56c7a9d0048e232c2bbe351bc58f889e947a34ca976ecf8b45536757bf12f39be622b7217e8872ae6c8bd5671e03b711a4cbbee2c00cbd79e61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b0d93ddfc8d06ce34b3f66a11e6992c2480906b01fb5d165924742c113b41c9e828d90b6baa845500ef9371ea33f7e33d07b79c4afbe3e5a566e128d6a013d74fe0e49cff25c000daa201edd9bffd5463dd51adf59fbb495268784699f427910fa85309cbd1be84bbfcd793d7b3cf5c7e648fdaee0a524ad12bdb72faba2983;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h256a202f4cfd537d0e045ddc432810c50ed0978d08ced0160d792e5f5cf0afb1833669e18e715f23268d555dd3d00ae1abef14ddce549dfc69fd2c7f99a8d4825ee865ef298801993ed2d4e228333d1f1b0f2ec2ff9ae5e406e59b55218f7272c58a6a9ac48f12f8cf4d9f9322e6f7b38613b45db591ac9332abec64ed04ee7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59e3c0abe3adc028cb3627b41d5d6e30f2afdfbf0e9adbcf516ee211e5edd82b96624beaf2ec5ab57475a849697aed8f45c29a13c8c3805bb6c72484f7c8e3a2028a7cee17e628c63b115d190d2a8f858b57e8c1fbc7d07c98a7c6988c8c490f5e1c5bae07b673bdf2289f0eb757a3bc33e418f5610832c846b82590d2ad73f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1729394cc82065fadcf624506c9cd35c1052099945ddb7f78b30882ccceabc7a53c72faac376532b1de2b759cb9e463b800642570b286078d0d3f066049b55023a48c9e7df2c39c84b18ac83921ad245854372f13ce6fa85bfca41aab4f0f268000926df685441e9b135de01c9dbcd76d2309ae76c7ae24f5655462ed2ba0ab8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16d409f0443016167a0834660ccadedd2ee9ae52bd69bf013012cbfb66a5d28fabe3f59721b70d643c1230dd35d3e0864e02088548a0e983e70e1444199f197a7e81118d5ee13877fb47943c2ca5355bda8c9a3592c55d64552c03bbf5c895d7309019a23574e4c27bf363fe2baafaa5fcf5e3d871215b723ed2830f836422a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbafc536f970cdecd838966c30167b2e91477be1e2f6619ff41772b6170468bd3e9374f45f18a026c087eaa47a748a564e0d485958e4a810ac0eb61a2e8cc636ff6feab857ee8171d2a3e60f32e911d87fb09a11db3b9ccd4d5267f2bdd32f86c3a4029c517897c9d935dadc2b8e149059af31aa7b3e959bd72442086f3f90ff1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h323137bab96ae592a76fe8ec09dfc33353ece7c40a3ce56dfe3901b9c2d76bdf351b87d96231615ea32919faf0678eab0f103748e5653e3453629e7528c871248a7965ec0abe3d98beb33649d3ca28656e980995338f0b0c0ef418ad615766bd2cc1e18666cfcee46bfd13ba1290f85337595043b4538810ca8583f83dff2abb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8641a9055ffa824b94a2697ef47b3be0d912c068377f4d6cef72ddaa1877fde29e9d7470f3e8d2384d8606142d21742ad20e434dd08262b655d06bcfe36aa3741c971de571e316a47a2fbae41b5e1861209293d127aa6a60d93961f703cbf53a577f5f96d33db1c643092a2b4dfdf775e35ce8fe51435b3c60579876eb0f691;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6050dc597b229fe98abd8a15a4d92ab715255114dc0e2f53976b5681d066bdba50022cbb479857391d85f1bacf3c450b534d1954f04eb4e607c70f576e9d81346f2f2246081a14b6250066e2b72f9b495c0d7c5abda5e33c39f43e2043ba78d534d542dfcf0d04da1726dad9e148b8b9d60808b4164aa3b0f667f30f5f1394aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2e26b6222a4961a5f10f11eb89dcf8bbc29ba657b817402c8e7208abe1e148ad6f7f0283f4dd030df813bcf007850ed9bb9b78be6d624c3f72546b0a71b832b643cf20c3f0912b73a77728369d6caf259c009c7bfa75865c6a40e3701e91d327e5173f868d5995d9e66d49b113e533219e8e9ce30aaa7978b86ac8aa79df2c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1884957cba58e32f6a1b51f4cd385a97b8b93e2eb355966530b3ed43bdcfac71ef831ecf15f4b5cba51926a6b5482110c066b29438d8748ea2816d5a7f14c3036ca37075323b28c9e056bc396d06d5e36742b0b6b5a504341e8d368c6a73b5b4e1d420bb78e2b7e019ce9caa23c251f15f0f5c463907101724412ec1c78be8a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb3db99b2b1a759789949be82f2e79ee103fa165c8dcf4fd98b3553f582b15f3a3d6308617f666202251953a98bd194f07f7f9fc11be6b7abb174c69df02864680b0a54d591f6be82513ca6a76fffa7254cd4dd0e1bb4e4b36046b8c0286efef5b4e5448cb6a1156042b0892c1d2b222ca8b339971713cfe3b952e4919eaf59e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57d59282e94edf65e85849ce8cd19a2f4bdb5727eb6106063f3149ab5310e6944691abc341760d05429b8a1b6dbeda401463a8c19999250c1a27b6f7d0dd43da689088c9894704a6e2ea504ad595cb8738c866785075c693f4551591def79f7af4b758ad55f861f03b4e5993be6cf665054932bdabb84ac8af611ea5b2944682;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3faad42e4ed5c4f2d8c5ab8b3868dd2bbb4424475bc69ca2eb4a37a4c3971ac07e8c91e1687f2d8ddcd960040e7cfba2dfbc6e1c4ff27c4d073ea146410bec9253f73ac4953019e3a9e8e166c82e939ad86348e2028bfbdb0eca09064020163de91f25e49a5fea62994fd840c792e73a232d514fe7fe8f646ac58a0201fe1a98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b153de729b26fefd4fe62f8a40825acafd197f0e4a231a4878953f4c0279fd3b9874d3fd08b779dcf40b4185cbd694e5571c4683a2c41a049d7446e27393203144eed5ee38c2768ab90d170101b582c9114ec0b72987d0100cea8e5c2f9200c16d7cc27046f3cc475e8d40eae99e5cc246f09a4e13281a9f6b4706a109a9313;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h627a58a7d3ee10dbc3a87298572b6a0e5f4547ec668112b4a595bccb984d2944822d5eaec0910c478982f7ca5e300958fa173401a5097a2334eb6365b5c445aca5161990883e0e69cd19ead6251ed34f9b9e33d7a5d7fb67658b99b218f0b3b3b16221df5e6de3bd10f9a4af95b5c165a431e97c5d814c5024fd798543ac1433;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83720e48a7ba77f4a0fea4047133d02c40c8f7eca75e28451a49d7ccf1f3a1331167ad7f995040c463e7bedb20cb54962b673ac6cf7c24eceed123b0c8278acd1ee4d012e943f38712afae30fc1b3c75e114d533fabfda96779c2ccac7a5bb31793dc6ba4d5369b18c6066c8f34afec4feb396c5ef647bcc527e86bd16ef3b74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8903af20a703c9b98e8122996f339d7cf6dd7ec1b70195c75d01e6dfaa609ee43f69de9e536317a64b65921a8f52519b305e35b40d4c873e8827cac5a04cbdcb390601e8c6d2ec2208230d920581ea5ea4029d9a17c9817c9e6eefab01842c9a187a6a28b502a9dde6754b926da90ea88e4a774b13097963e87bfdbdb8384e22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa5d53f064f772a2560effad18be46aa5f7b04813658d42f5da0adc799f04d71f74d27c9789fd852c9e46aba52b417eb8a5599642a28004643142ac24218d17971d2d1f3d3a93eb18b64371cae5b5f8b95bd1d756610c7f334fb8bff1dcef3f3c496e5f9e1223930e96c97e527e3a4aaaafd2d04a968f4f951434a0056c67c45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4822ed95c7fad94d7469e2279289313b289228cf88c5b62519c61eeacb192c9707e16bae9dc1ebb292e5165217b312e2fffe64affd5c0d517193430a8234e32ad49c33dc150ddf68cb050c65253acd32e2a5e2b736af7f0dc4bb50bd687c222f06d1821e6008bb62ef2701428179ca34812032d72973842ee704bb532fe79d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27a353e1936064d2bf7502414504ce36f94cdd192e1602292d1479bf3351c2f50a5f87dd736b3558b5efd534d90725925a2bdb44e57235baf62e371c878f5c67c2ad9d7f3a722fc0b364aeda713b8b4332264fc77889c0622cea9a4eb2580368227d6448eb48146bdd092ed7f88629282541cbe794562bdb67ee8f09f697f65c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5728de6f655365749e8f99627d42fd1c7d67803de5a6a172fec611e52945a622e0eaf3c88e9cbf53ca12512507813ef148545eba49f7dade9830d0941f80821661ccb3225eb86581bda115b63afc54bcb5825df06d15d5152daaa56ea797c986c7e1ee69da47b8c44ec1c7f6c83e974ded9ce751c945ef3c9f2455504666021;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b8df2dc7ddf6d89686d509e29226fa37a3207a843b43bfabb9604afdc15f678b1ace201618380a078c7c2d7b2ab3820adee4081e57daeb90cbf2c23ec147982a18969ecd12e06e625ba4bdae7900e065b02f7a536cd346c111bf10560d9bf12af8780e0429415591933b914e75a530823574077c7802e267a308f003915f811;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72d7c5bf6dff847c498a9b5b5ec99b32ccd0f84092b909f6d3f9f2f67195f2e9344a2da0465c38cefa488b4c75abfefdbec581dd20a3b6a7c08e6d1a0b66d4b0e0dece32694b53e8626cc32337e5b86eedfe866f015fefb5f992008fb9687e0bbe9420895e5602549b988df18f2515e5ce4de2ac9d6fb03097d6ab2580e73eb0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h597ffa0e14edc414b5dc31add40ddeb9cf8399a60a6b0a96a25417e0656bd66e1302292333de3ce396f062435742b2bf950211fd20d37134a9658139c9321e4bbd549bb19d7f23023646326aa08dd24d4a4ae544c23df5d5a1b4fcb0dd3283ea76ea7cc3952aa49632b0c86abba0bd8dbe8407698013fe2b16009d9c276f9b5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b7a1899a8c5e6302135f5c6e9dffe944368fe197a0e204586101e214a711da0ba12c6a8cd58d49930bb7eb315d3eb0259d2dbd2bed67e65f57eadb16f5d6ab39c12f6b27a696a8961bcd55f0dce5b6f2b7cff1eb0313cfa602d9d73e4db51797229cf4f2ac478513a6183715eba92cecb9260b7a444ee73343aa4a12d8de379;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1b139e8b12a1e2e0695aac4e218c48e7c88bfa2fbd9c53b058b43506c321c2a17b6b0743568704767e8f2c108f0cd74c6ee1c899594c79902211613146b52c8f3a9fd98efb05b0082522b3e0fa12688eb2ecf7d80611ed74fd68ab37b075c2f705746d8eeb635b3f8b886a7b91e3201782791d740b11075e192db36cc9c435a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaa1b8f7bcf1360c4fe9c0889a6ea00eeac65f47aa9d6a6f548c9ce15f0a0b6044ed70f345d4760aae3af5dac997ec382ed238890c2216fb8f84872107663be2d8b4f71910ea748cb8169ced7a29678fff1563fdb895c8e03284fe18363a9f31baac7d5856f7a9f99de8f012660996bbcf20307158cf3a544e77468a67694e6e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h910732d484edc76d5b6d794d2149945809ffe878d38b2fa1b4f48f48fa4e25ac361632391aafacf6e887a1bda80fc6de2f0a1fbc9a4597abec9fc9b09c003c327406ac5126fd32e74cadf4b6c47fe6ec38b28cbd3b68bf691680720b6f7204f6ee1f7c0d6cf7e8ee7ce6cad7e208f1cad2ad358cc539f239ec39d0c02177eb2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e8f1c0064a800eb250346e5e35f8960f5026b5b2147d968ab3f5a8af52ab2c3ac38b4c4cfc59302c7120620307a49d757a54214c42a78b75240f7524983e35c0c254da039818ebbf4bfdfe7417ca8b461291ce64819c9a8c7508922dcfb25cd59d66e7fb478fd7eb0db9b9cb250d11a548b9ac61573d928896495902537c310;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26ba573616084d86818d6f84f6d33e5f42557ba3d92a5da974dabad0f81d7db5770fee2409d7ce79b5466dbf03bcda1c093686e2642b347dc755ab5edc0b26f39c585f4161b9a06a79555a5acce6d5d1ad1f1e931a090c03e6c306cd34b42c3d373f001ffc433bb56b1f310cf25c189029582e740f9ce0158fe7fb6c9efc1c9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb3e98fe705b2830e6fb07901e3788100900870e4c84d4136ff011aaf640d29bc0787e9b08d2a0ed525cfd89f91c10486e5fa56a91948d3ef8c5e3bc15dc83fcfbd47a922404c80149c769b6c8227df1f1e4bd4561640860e5cbc2324588aa0a296caa78bc5a8ac7e73b4607129afaaa2872b2144bb519146cd093bc65f68991;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bd34e73f00d42b7dd2d836c4fdea21a7626cff54eaa8e94c70eda64d036ef8fd707f3012ecaaac00da1a3c19992e15a970b10f4649645b69925131702403ad54c23d8c19dcddcbd050be14ffaf0ef03451f4be00bb792205a582d4df85b30c5009ed83074180f8701a2e7b62e2956a266afd461d3984e316673f0d3af8503c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15bbaa7523971586d83cb71b083e40b3f6a56fa64bf621d671e97db26adc5a15a47c7f5abe84e2bdff3005cdc7fd9d35a9332e6597b0bbe828483451b3eee7bdeafdb48b0acd7cb4342f2e9548e7d2a938ead02271be15851a2e7b549b9eaef9e3a8bfc56bfe0f1bc7fda218b327862208d01d7b3acf8fe2a727b34cffeb6212;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda6b9b5191e22056e0cd289797555ca119be9af367e6528dc9f8bbf902bd4102436f1231b0c3e28ed4dce80a15abc64ba3ec9c410d0c8a4e6da04c73f592be8be8045d71f9a0203be073b66b159e9b62f0487261ffb19cff50c6c55cb4d41016837794d3ba2d5730db8197b9c6fb5c59e206ab1fa804fd2e34d0cfe6d03069ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h648b199a0c5ca95cb735688336fd64eb1d098bff0ee1de43e923db2cbe13fe7bf22321fc6a0f6c8561fd4dd696a343dbb422bba9bc2bac690d0d96217e99690241c76086ab4de2ee840da869551c3a957392bf4a5a5d7d4b4623862b48f00f6eaae983f768e5f1f1cd703b9f114ec8d21782f7f6522ece4d9ca65233a21d29b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24169d51792727d3bf7ac9847adc3af0f98a5613762f9bd76e7266779436b5850c370b75416e609174ca627e740606d9b398417759b34ded09ef0ed22bc6f7e71b6e340dcce5545c940a8ce233b5f99dff88c2cbec039a8dc983a966565cc28efe54f299b08d598efa7dd33c18a59c964565ff3bc3a08ee6373a9e920845605;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e2793aa52964caac80ac6ef0b88a08d5cad0e2d1b867bd83c7179ce2e519b482595dbce9ba66c25bc9b211f669f017e79b1d53307b17c6a61b7f4e37248a52293d7916f17d79f4804ed3fe16381c3c817896ebee523e15a26241d4564cd9a6550ccc3cff2a9819be55dbe9a1751f1503d59cdb87cc280114d41169979255449;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2aa351dd2d246314de467ab515b221ea9ccb3cc3fef6e58dcbb2de3ed1b97a888b91a972a259c0ce1d0abe33c10f8457b237ab83ecd7ff370d0b8a679c0f79e1752fc6e0d774b8c9f0eb815567beac9f3250a93d787a7715d37b36f608d194de30d1f825a11b9301a6990ede95ed18960ced7f814c374e7734a48fd811fba42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h672131d825018fc7b41a45936dbb9e6a418f33339f066c7212d9cad67c00077cd860a9fee0693591b7bab9d972777c07fb90e489a3dd49305edebd9f6af00d3b71516caab1452bb12736d8e16bd728f0ec9f2f5a60efb3a017be34b8cd1a4059564092a7c7ca28cd321a0caaf504fe9e9ecea479f4833757552a522904b99e4c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40baa368d493e9d101d3a118985202e5a3965b3093959d6744f3ca5cc312e818db1103f4febee934e03b2df06ecf95dad089b514379d7764c0f5e16086237d3fb2e8262bb56322b9aa3cdb9616c97ee148ae62a25cb7a7637f6f4fa59dc4a60daebe44cf6b8de2db41a1e112e9c35f1ce01d9ba6bf17fd5bb653ce160ac5176b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61cf12d5ab2eabfd0e6cb335a0ce7e9ed95509e7ca0075ff8b3150abe005db097814448cefaad789b9d04af7413590fdeb74c3d53fb2436316442670aebf45e8cf21bb0e7f1142e8f128da49cb445e7c84b77f0ce87147769c61e46d8f8a54b71a395c5fb7cd782afcb55e50d2474a7c0ec935ccbc5ead188f06739b2915f41b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10418a3d13584a401c109e1bd1b34c7579609d2b4ad1088a2a8f9dd609f04cfa267252e4832134d9a7e139b7ba13b5330746c147270a2e33079cb51570966b5b8213d58a79bd4ec77ca8c72ead33251930c9d7284f41e4521443dcd967eb03996bb1a8d284433e3e0cba49c65b1a624b4ed5d3f4d40f1cb37f517dbddbf19e23;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61f30a27d0f4826250b233f95a203ae57a1167a0890528b86567a986467a7d3e5cba7874d00317d7a2f39f56ef719b11c661ef0ee71b142dbb6061a249ec70738a420999ac90fb65dc0a8e819417af58d01cd0d1e834f0cd0c2dad792605d71a048f4c3c5238b9ed90e74d9b9d3c636519ba8db4690b516221467a233879edb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b04c24d04a12edaa987794b2c821984f2fe4f3fc93c11effdb55ceeedaa2059f74baf973f7b4fe6caf25ecf92cc5f28e737e17efff956d9fb8007cdf11f6c30ddf80f12b784117aa720c5f7b6c2ebe0b9a871ad5ab79d5ed5baa2e37c360cc0c463515add7c950c79a6b3ebedd6ffdf661ff093fac406823605691412f02c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7583d991a1c279da42e3965cda2d1260ae4fce849d34106897bc1a3e6955eff9c9249dc5b7dd5a94f24799df74f3b06f8337ea6f27e000ba00f2efb614f71b49311941e638cfbca5b197fbee5a54f5696f425233d35191ef3f7c8ddb1f84164bb609234f7f51fd2e1dcf9a8ebc00f6e86c668a71bfa59cd1a2a92741f955e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4609bd2e9ca1ccf5b8e5a3c7d7bc5213c4b40de2ebfec025a4b921287023d40c04b065b093fa8b5a7856d6e8ed9e077195c8354cbea50fac389b6f4d5e13f44621966a61aebc359a592598384a9254221fa08e6109ccba1b16c7787dd07c8c554947fa2316a848bc68a78f36a9ea3202ec758a114bca7450ce846647c690d21e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d079593c97df60c1d4cd8e4e1e2fd17d7240aef93ee579d6cc4505f61253ead9485be68a1bbdb8c4162d2b9a736569e254a6827aad56098f60aa78667f8c2aef677728432e4b7567d8d46218c7cf3be62e05dd66d405c79a8efb5ce3ce142841fc7fd1631fca137f74b3bd80030fe567cc7f80d4a849c10885867fc05609f84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0116dfdefd532427f29d4daebf976b2ddb6b0cbb495ae4f07225277d546d7c37153e0e21bbe1dc42756fd34ada8601994c00be414d80eb9fdd5d8ec18f0964869b7f952162bef4bde74f29146ff4a14634aa2b4d14589a27dbd92c5be3f2b1dc27ad3f8f038da42ad15bf037835d4b283b47448b524cbff1cfc353ae715409e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha417a3870d0a9548e223b9ec0777fa226cd48db7b225fd846744ddf3b9326f55db58df4c9b673dc24062a1823fc4b066b152d3187e1505c975c02ead671c4d9d811ef3deddfe0fa2394d250e234bac033a39f85407026ee79dc99ba6828da128a5e92191a3d8db75a6960a5c66df7a2c882f1776f83e3ac84f4dcd15c2d494b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b5d8de0afb1ff476c7e7bae055cb2a14000f9ed9a680fc451c87dcf03c0e48e05fff8183e1c490da4efde0d7eb313dfff4cb87541ac79ca99e95c158e498b49b423694022a51cc60a5e3ee87395606dca5bd56d1d26e28cbe0f8064a0e8d6fe5fe5fc4790750d780052c5fa37a33ca4d612f3ad7f0de6c3f42ba1037d35331a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c87e73eb3e57b4be96b5ff1834820293e9a37c519af02c7724ea65493b89ffda5fd88c992472ccde8643c1cdd7c6449f0fc38c4bd897ab85d51047d26b17bce4e4801c2b565d418ef4840b2596c00cc537c02036327c0d7c21f7303f86e5aa63593305201275b8fdba027b871e8834bbecfa0b42f7dc676d9d5ba8444ad7da2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc48f50d0f02098b819d863956eb441245682dfac610b2b339fef9f9e98f2f9b0beb696f4546548cf7c48f40fb82901c5fa71bf210e0ecf259d42ba7b9b7ec591edbdae7ef6880404dd826dcacc332e1ad3ce388589657d944f8ba95bbaf02b3cbd78b98b734b8ff91a9c99ee1f439b2155655512819dc68326a414c6364db496;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc95c383e38a78502ad92278538d6c1edea327f3e9e154e182f80a11afe16ff55a077c7f17d64e43e5a5768400b543fb43b570ba2f7427e6bb6a786301525387de7d2204c61947c51853455ffac4087d051ec84e5d9a0628d6aa81b5c390c8adae68b6fae7cf8386a8fc8594e6914652d6e69fbe52d544f2765be1d5cc6003379;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a5ab3098d3d3815aad7bf986323becbf1f254c4eb157cd4e8c15627e5be2bc1704b5aec41b9215c0e31df1253b93a06e94f62bba5b11622ba251187c4ccbd353090e9023b914b0b6dfb6841f951284e18a0383867990fc99d225f68d9c4f4682eb332749b4aa81ac56c913a09fe635851cb83ea40c518595e5f1f2076833066;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35858d4c5c960ae71a01ae96e735e96e3756758e0d43e4e9050a5fb8f685a917a63ab08fddf36540a25f37d1b59ccdabd353f2ee7e19f567ef7429c19d187af89fda670f358daafa2e8fc231388d9e5572ff3b7cef6aa96e8ad82bc1229386c0c2845649cd6860bba69a9db73a75d4c7fed57332adbba0d39834d9409e275245;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90517bb7110a864bb693e749aea4eaeb2d96ed34984380a1a89fb18e1f52494f89649ae7fc8f3e40ddc6a482745687aa0c312ee2ae59ad9bd21732c359b262d5ffe5fd88a4909d6f5829dcd6853b8acf29367b9a9de0694728825f48e043bf3edc64626247904c92c3c47969c0fbf8962350e266efb3d41f23208586029e2cf3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a6db77d8d53dd66541b5cc04ab547a03643f8af6e77e55126286b5d4bb246832594963902bbf5974008ea322923fad31795280ea39d381b7beb19110dcbf0d11a61d3395b963155e5bd8fcaa07b4102aa880318b2dd6ad9259086ae377f769550a955798a6c324aacf730644058d82a46d6af00786c8f0de5f939c4a167470d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc51a148bb5311a37894ec871b2cd19ab8e999fd20cdf3d58e536c94d77dcef56349320ad6bea6638ad4e944c70491dbd258988f91b83d08d7abcbebab6d8643ef46341090d626202355543ac6060b8d6c3c8a6812c99788113e127a17a63408b3c62475cdb12b32469ac6aba96faf0ca068e67abde7ab3578d9e5979e2a9af4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54ff98cdf5ed9299da2ebd7c7bce52b9bcef775057d4e7034ccb2f66ca6d3dcd76312eb08307f69f9e27953dc59a7bedffe8f41aff4038e48de35a21d563204be1c331294d6f2e20e22d822bcc9fbf5cccf1befcf2a279349c623f2377de544c224381a7648ce47b29fa6be87a23cdc1e5cec59d98921b0191dbdbf36710623;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4f82814ff6658725cb3443c19d7ef8be5e97aabf7d00e4a6f29c7114725046ef3f9712cf841924e6706b48e7e6e37f72bcc200a0d9b4d6c6d8e312963a5e6cc253f82d7248b56616d2d9178b923f868193861e4cbb1100c14f23d477942c9e761b28a32d37a7d9e2456996ef1c12528b57f51aec30578b49772af01daed71b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf1b40ff4602900e18858cfd2117d279028cf11112829d35b4af053ae3f33b5e0f0fd6e0cc23bc5609c7d93f9e89e661b98c18b86793c21ecb6ceeec146625d3f42494511d60d049fea269c7849f1d242958e5eb7692a6515a8d95dd3916c9aab0e917c489bf1672ce541eca47b3b7c677426a85a3e0c02aba54fc436e5fa75f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572e9f4b1a748bcf42fcf0303a2100294231dd7c0e90998a7aba3ff56bb7e950a5fb0e1a92753e3566a88057f9cc4df36db46d5b0bacaf1394d23001bb669ccf45f76f9deb4154e9a0feccef6cd2546f1ba3cf6c20b5566d023c8de60dc510962d63f0e44c78538ba657a2feb6e135a75abef4ed2bf41cfe8cf096fae9fd5df6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3fe70bf1a7c9be0ff3f6b8cd79cbea47d11643bcbad58f5cc828952a326c3595076eab543ca5e5482b7c6b873f79815ad07b87e1f9c6c1d33a4dc6f485653f8aa85a4fa2b4e32084dd38158afa12609af5b177da35f6ac514f38736d9da5fbc2229a14e36003b102646a8dbf8558c01a50192622477cefc834d9c13e1a1815a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b78b47cfd302ff491084ee9c9b17287f2ad29a402607bb8aa55a47ea925f4c5db8188bc8b3e0c9ab4bb55df03767c2b5fc3199b184da377c1ab9840c50330d9354b2cc851070afa0dbc3738f11dde5ee29667ab98f5ae0cc685c3aa88c5273a66b54499167220896701c14fa65d86bd21799db091ec002748db93b909d04c65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a30c8cdfd7026475fd992d54c2097ee024188b873a0296b73c8bf51cf35d9d0fd745cceacb8b8eaedfd43b33eac2f843a757f28e52b9b2c327f17a1a76da887c9efebd7e786005dafae657f37031b1642fa649e32c7640c5ab190adc31f4c0d1836849bc6ba55cd335cfd1d404188a1349760a6ebb7a882e60f815949d3ad43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1718d8994de062d9361253c7f8a9322f61bfc4056a62961748d69b904b5d0d59aa9bea2928b442ae5b826f92a36b8c65811e31a5cc41fa02231324daf97aa5f6585fc39f7be54580d80b1b55fc62a70d2f80e92324dbbd4304bc9adf05169589b9a038ff7600b0c56a3ad8d976beb2cd83e097d24cd9578536e659e71876e40d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78aeb227648481ca175c208f7da953da318e9a5e2e6835805f8d1a0986abaadc1f24325a0fe64681e55d26b216a56edca8786675cf6556b60af1e2e51fe52122f6d5385ad1b235536a29d03b028db091a1e640d282dc34f21ab251853f3cdc2d8ec3d7598c1ac9868316c8b4d028bbf3cd2263bdb4e6b58c66d7ff3deea93da9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29568f147a6330c1a515e940381286080f40243e3f8f894e6f4020251c600dd5be67aef2eaca142f49a5bf684f6e55b56a19864c99a3f25ef6cc0e2a5790d59f66c2cc93dc1068d2452289b5985ac9a2ba51297baaaff875c87579dc8ba91ad69fbd27e864599a8e2b2d018245f79d3a51dd4321391c83c76ba50a6f9a8028c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ca99292f8d732ae24d4f753f575feb12c9cce7c51757ed6c45aaf824b5d3bbe06bb6cc35f25ee91ff50dfb3980c865f01b3796a75ec4e0231a72134836db39d9f6aa4231288d44c137678096b927d11a88a28b4321f21d3d138b16dd3d13abd6c12b5f6c87197b3cc0801098a8933db2f03e27e9157d60d84475d453ad0ed4f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0c9891a0b117093067099c9d35476f2ad3a9ee5d205e95d49d16ba0f3241319c58a668027c102ef56f33b2e0f99ff84a573cc083198b3f262f69c005c9fb5eaba8c087d443fb0044e3acf5410488040dcb40af299433e6b84d709532712d4717e471425c5045e370a6a9f62083acfc6e697d915fe71ef207e3cd6eaa557003d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ad2b58520e93bd2be3d3520860df2229ebbedded3c6049fa819711db079a69e21cbdaefb1437eae1461924d32d9fb8085a44a8e69b82a32c05349d84f4fad6f6fc9c71026fdfd64f26ab0bff0d4b3c8f04bd11ecce93bb9510e7b0f24ea64ccb8beaee28f0471856e1b3dc51a21b0ffa6c3394709faa92e88d64cd8165494;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d56ee3834cad2f64b5b79c2030e2e126ac5625cc313a8832b5ed211a2af94166e0c759133795ff4a0cb6e1951838b3b68b5c5c7682f3be8272bd7c3b2800a413fab30bf3f0266e67a49be4cca7f260cad20f204acec1ee72646fabe209a362a9488c088201a0d001eb034316be8f97a88d8e1cf2049930bc75fdcb3ca3ac340;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd08157599bac0435c387aa158a2806a19dc498e9b201c62d7814afcb70c1eabda0532d30936b2b979f6a2dbe704024b1cd9ddc17d1bc16ad1b31e5a86b6f40f38f522bc4dd4c2d57d5a384bf23683763c556414140c9c871dea95e21f9ff527335c59972dcf36aa8b436bce2b749b2b74a15199575da52d8155ce23091193c7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63fca658e7863c68afbbbd32d78d3c9107deb09d16133ce268d7fb730b2ebfad450e9c0732f9889e85c0c05e0a21b204cd59c063aab17054cf600cbea0f9343b8f21cd1f09f1c73720685e3f4d62ae6a983e005e91d48b559fe6aed721c5f33b34ffcf9cfc1fec9ebae4021afb16352df762868b97236ed04a2a1022eb5eb534;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2149da5566193df4c4f2193a305ffd0cd93e329b1f805d6d23d000305d458612b28670fcc362d647adeb59d6c9dec57ce1addc57d19bd4f66b33480e1ca116e1dab6dcca58453fbde4ea6416eacebe0749ec9a7f8a2af46b8d64c98f0268bb387e31ed4644b6787cbe897dd5e6375346d14962ef9a3eea8d06459012900e5c05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fb01d06b9986cd85a07501276a5aba74df473112f52d4f2212a90057b384357e99cc922220cb0386501aaa6aa93c1b9689f762b90c2245005e2cbd53959682dbd6f5d4045992317856a51d691907948f95d65ffdcc02905e800c49d181df09a9d16390405aeed33456aa8d5d0433e89cf3290fdf228ac59318f8a30d167eea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42b3a02b01513e65ee459fb9eb4d7cb0f57c5961f80ddcef1319621a5c4681e9e62f883faea872095346faba0145474202b10163d6e54a739519566795b2899b03b1428099f70fc8bbc1e75cb5c14cd835aef1615cf4a45cb15138ac10f778f9dea13a8ff8e081cbf8e550557b0ee5edeb18cc52f3d9c413c4d29267ef645094;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab0d9f2c84be2028563469f58837f67610d385aea0f572f79767b3a00fb5a2f18e627f9f0e34275022a928d8b0d5bc2bf84bfe040c0bd242d07dc4cb6a5cd83e479d4f9e6facd7cc7ae855666ef32299a17644e56b7dbd10057a7955c85c4f3a4dc6f8fadf6270d9d59e0d3ffc57c835c2cf2483b4aeda36d9c79d25e70f9cb4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h651c6754737e91d3637dce6c7a5bc3a9a228309188a54fa43efcabac91b1989029bcbeecff713f7112d6591fce558d0366a6d446eb99dac2106e23175fa32549fce693087835e6a37bff9ae765b83e1dcbf1f1d5fef4a09826423fb354835b6e1e3c1a766e552fde213132e922ed54d46043bb35251be900528ca20c430c57d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7041d0300ae05df6320178fc51e58e44fac54abd4009eba7473a2a73b79f83aa6ea9abd6b5a3885088a83e24cefb02c94fc63ea932403b4d1931ca16e4449951beed813a373ae86cf28b489bd8cde5b0d8a23039f4c365df4728319f9f054039695b4f3d654bdfe7fa4db39229bae4e34c62efce2793c89fb724b887e1fc067b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62bd72226a7ea0d3831c2e0037d21aedbd06c955863a5d3b1892892bd4527e077ae4affba858d880f81c2cb1c1ad74e9d09c47785d6351a204400325e5d352688830b7190993ecd243ea25e86a4acc6e3de17af6746fa6cbadf4e083e896499486ba2f85ee3c977e4d490abd236fd93aeb910b1b60730a63eff54b0079379897;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88dd83ccccd7d72d8b4f8192c4974550e48c3dc03fa0de1f0dbb6291a3262eb9f570ab73b7652f33a176f3cba6453fbd2e6da08975501baac1f4bc25c2fc1a8d212dda0d2c963df9dcd7b7c7953c5dab055de3254ebcde92266d1a34ee3787542a7f498c7b4e350c694aafa5cbf4b51d2f944222f196ba3847dbdd45e1c4a610;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he42763e99671c0ee006c7f2de04cf97aef9f9d1cf6850d2e17aa95afff19f62ad851169f45eefb1cef0d81b247d667250ff927cfc3cb05d78f09f243c25abe064a28cf944496bb2b647c69f2f2ec3e9a37df4708453c4dae5a71532fe6bda2627f61a95c68e59befba289dc2d9a67df3f505566c0795cbbe60c46d96061d087;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5761e3d2cdf4433a3293af3406aff4d6e3ea1a3fe4cf9cbfd2334cbf797d1f5fb07c29eb4207578f447147b6d7dba3cf8cce94acef3542bed5b00c30d0ddee820f271359db9d9015c12473137fecefffa3c268bc1c67d46d26faf7c6ba187433e935044175a4bbe1909078fe614eb2238d289df4e54bc6a228e259a29c4fbf86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf6db02fcc83e4afc37ca6b2780a0beeb971856cccf89d299c22fe9b75faac603ba6a622578490a9c226f94f9ff934be878aab1b7c0f2574b76328aca5806909aadf4d01e387a8bb613919f8354db9dde47acefed4999d4cd48bdac4f380a419d138ad3fe3968165c33cece7616cc4f650c3bc6d6522b23f4bd43c478fcda094;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1861436077ac3e0a836d509bb8525e5724ce23903d41799f05dcd5aa2d238e1c35bfb8347602efdb054ff8a303011cc46a1724dba6e6f42d8486230097693d7c75c66e6d9c88d87da6ea70578b5bb757b1e8e2912a8e206fbe8e801274f2f4e48e9d159acd3e16402375029a725e47bd0c78bdf1c49e72f6a610343a5ad93060;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb566f88421f6996dd331b6beeccaddb54fd004da9e62260d33e28ebf4f9eccb9376e071e066d45113368d378893da1d55e54b612cc60c30623d080730adf548bbfc0d14499c2dd87bbf867c299539d0305def9e4ff80a1ea103a773fde53c33ffaa7f8edef30829f425d1f6036c0cbdb3650fb457a368cefa2921e944f8bf922;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7edc1aa3ff8a52cfc4d47ba9d6a861581a36b481e0a21a9c796dab7f9529d290e3c541615fd374b5682c9b7a26de5cb70556d702412b6356b9009b0e7a3351aba21f814e93911b6f1bc97b7bf998f8474f29bdd33ea8d94b5dd5aba753143b317d12a50bc4877ec41654b9287a7b1fabc2670cd0c2141136ab55d51774782585;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hace1d3bd4846be4531db504232f13b3e447191948b28a79a2be7e8d651ce6ef67f3acec5604fd892d9d87334622f97350d963a8b396850a0d26c08e3842bb06e745f01235558a7d597676e16ff64e1ad1302160fad770bf5416808ca729c20cd0ec76a4c3fbb5ef36beaad176074cace78c4852a0a32f5050eb2d0f4460399b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac4a8f4de4d0ea9856279f334e579e065f4772154e199b28375d48e5dbdebbfb2556bf17445b4259a0f01d613e8c122e31674d35c7777ecb02e03e2d08d689ec3b3a52d81653fb7a57d31ea4835267cdf0ad4789fcdfc4446f8ec196b3b1e39b26c1b3b738ec88e25e055e303dc7170faab827af0675de96238c8055a1f3e15c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ec7a6b64e773be732c579159b141e65d273726006c47c31210a08616c7652564f6929637937b323c39e8bfaf90bded2483ac5c9c7ce600ef77e6c897f96a041fb89d8758043b700b6fabc5587728d536aaa2bca0d347f42fac9a2f7a34378452a7527412aae4f7f9fd6a722ff2bcb69a01fafd11bbbc3d01841731c78e574e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92c09c0c93ee2c38e29c381d34e37719d5c4f24e249f170442c552d7270b35bc7130280a4ede8d00c5215d7d7540df91c65161d9c9700e56f064d275dc2fb9d4a88c5120ec02c6e48d6f1459833b10bb2eec770798b97a94573eddaba3368e8d874745cc88b4ad26ded851e1c2e5b371770a3c5fb29a0273b844dc7058f98a16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h111bf336b0874a079b64578a4616088dc6007b63ff9cff9872a625253f0ed6736101e089216e5445ef41985b3caad54c03d57fc89ce2d76f05d3db2d324e755526ab1a83a6e19db2523495f0f38905039a130755589d7cbfab838fe9277c9f2cc2aa989598c0da2af0e5120fe42d7ca81a36c75bdaa31ecbf576f9ec8f562a97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4e97604272818761f3ccc9f32813b87f37aa15e3db058fd3e38486662a2f40a26d8784bf48ee31860a0bb8558adfdd876e3cd2c177313231e30f4b52255d9f248a0d79eb097ae76d78d556244b109d149f0cf3e5aa13b7b8c3e70270b3bad681bc4d4d9ce69b0702566fe2d3337fdee7e0f807ca9ffc780747b476750fdb240;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9690bd706793270cf063fadcad20d7c9c7f459396f41c313775e92d0fa6c1b0abf2cfc45a523fe2fd56ac9a76d58389210856037ff085f23946bcc94ed101f138b9db917d11f2ae504a3d064dab106a5dd5864311dad9deb42344797a2ccc95c526c597019d526d153dcef6a8575bb35f0af003dfe92fd028772e3a66e60802;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h317ad859aa5157cdfee16d2b52959426b48980b8456c3614d6abc052e7b6463cd6f0596f8269bec7a3d9a1fca67bbd31d52bdbd17df2749182c92827eefa01eb4d29d46d850aa5c9464fcd3d439e054450bd9cd1ae9bc1be91a20334363c7ebc2d135c659de8780ff990ff6eae17babb88004190e0bd4d60fa1cf3d52135c80f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfa9e6c5ea147536d863b8f784447b2f29a77cc0c27600c148ca4e333951d431f0a5b0200c76e06e52c76c8d273d512ba02b5f43ae11896805fc225e19f69d1b6c4d0051e41ada88e6a129253ce3448fd786d5cc2e15103611cf86342c3a0c867ca2e51450feca446d2bcdc6a93e18d477d431e7fbe99bf6f3bb1085a6c7e098;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56de4f5f1c69af42fbf35db0f8821dbc475d7b12240ea247eaeb793e786e662a95f3681a205541c44a193c4437ec42df5c547c50e54625017a31d48b84ef9fc2154c7d737e4a648017bf9937012ded759157b02e2e48b7e03e35af1ecd531f28bf130c9f86a2b33b15a192db73f11be35a16ecb96dba815b527cb6128dfe35b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h209f1f947dfaae79233a31cc8953ed4788e33d4764e15444e5c68e28abd4cd520345d006f017f43adc8527f0d87470daf9604f63bd7b125b001404739eedb37eba33c2613babaf6bd0055aa372b8d1972b5673d123c75249ac696584b502ccc36654cfd744287780b38ab6fa6561e39298b3e12f086ff5292a1941a36101c94a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbebae57dd057c3cdf1d0f92e8b6b00f1f7d0b5f2df21d3ae74fc87b696c1d6f8b5f1395ef1b4a88c2a1eb3ff70dee740bcfe4168cecff3285ddfc9ea2e88bd2c516bc42b473226f90bd79daf81f8f2d2f0f70dd13d78a8f5b2255180424b3681f9406263c584977d437f078a0e376ba9b5db7714acfd91b1fc14822d6bebf221;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h439dce97b230a5eb5b3e3872ddc6d861f3228330c8ac1f89c76ae75a8c44eeb4dd7c1f8d52c947c9f9b58e5b414adb75c8ae6017fab220df9c706fd49049cff357e6bb8c2547005fb1ca50f7a3cefb72b6929d9634aa1ff885200ba565b66232a5ef0d2abeb3bb72c7938cc553e90d93df203713f8540a38f51bd24d76a674e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h215efaa55f46e6cb10d11200a65de433f132832733da74fb3404d99372a680c7a1bf44a4cc78d5db1a6b16988a38259b4fa1a5c1f17b571354a73ffbd185fbcd4d4c4d3b2bbbd0425f28cff56c2cad32f716f375173c7ead10712cf4bac0de851a5fbe87cbce4fbcce1945222ce11e332ecf0ef5e250ce71d4da6ba0c9b12bfb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a6036fcf19dbe7f6ca746cc315bc34274ffd6f6c331b36100e45e9384f73c4ced25ad4767b7697ad53896c72760fe013c67476f93ca5db990624197639ad4ee85487505f29c9c86358276ee6e9effea684020afc84ffae67644557b0bfa86022a9bb7bdc443cecb7c0e84c2dd96b88bc1299e80f85eda1edeef2b6ccb91823d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h154b3b4977f61b0684e358b73ea98c255cd8271c09f56c8f9612422e010554507774f91c55713a8f73eb8f9a2d206a18df2c894bba0a0a3e2482b1bf4e19fe3ad232097af06e5e3e098c79a8b6f8ee3259a623f4bc1ce79babac78bd2338a87cf8c401f8c9e6086a3c82276f1d51389305c3029845197402ce926a73c093b2ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf75c954c5ed007c68175f4025f23b93182d095eb01a3ba9634f17f6b22fb40da74e319301f74c947e424b6135217e25f72bc23d2d5ad68c80e3542e989b1f4f71706d6ba354a4c989e081a957f91b1228627d769ff09ebc1a7dc84f01a51345d3e75547b9885a5459b2a39d6d2851d6e181fef5d51a3adfd4685e9a23fdb188;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a46216769e842cb41742578e16bf855329bc14705d8dc63d291739f90719fd0356c6720c5b1e971e90c847b545562121d1cc8e059a0ee792e1c570c79e771ae3961688370fa97a91a04337d2f0cbec461d50decfd8e68c009f9ba63908497e4bcfc5c815eae80f838ec595072aba4096abbc560f3b8759239f3226758f4600b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd817ee38efe6235032159890a3f02fd5a91f87acd820112cc1cd74bfd12122914ff5a3d9f1a107413d2b23f07d198bc792ba99020f9b6df4d702e0db44ad42090059cc208784ee2a530d1b596901ce8513ef4b4e3eb95a14c2c361eb2aa3a4bfa7257fadece766dae7e7a16e18fcb3aa42c50ab0796aeab266484d61e4b0d90;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c628b6b6752c4a8442752bebd67ee3527ce7c34696aef3cef9e82d31968eefbb478d3009318076f7d0247e83708967c7fc038555bd118efdc4aed4f6fdf9b71ad3dca0424304bbbc3ea30bf35a30f298c67c08b4abe107d655a998c3340d96969cc9139a8a2e8be52e167d8cab15384870076b5e6384d4a87c66a2641ecb391;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b9a1b512b8f86032e1f4251af35efa1feaf16546e01da10cdee68e3db8b2e81f2cc9b8501877878ebdb9e9d2183c95b055199dd648cd1dbf6ba4572755d262fd121e911893f5acf615df0282430fa425bc78752f6431867e708f105bf3d94e30dab140289876b89cead62b79b6354abf598c83a22408c0ba1c48e73b90d4321;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbf23d4f80fca2d1d6aa1a010fcd3aa62321a5820a542c37398433e4d9f0c412be3f9297e0f54df5570949529bd500929b401c39606b7bd499c4f685db4253636fffc2cc6110a928c4a8c436c2eef4f1991a086bf211f21d079bb0a9c1d67c88df6bb94b6a9c87a2f121b4365d6884664f7964f964eceabe540a80f69cc6e8b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97b3e8efafeeaf158a799a0b4b6f933c43d39d4ad4ecb49d21d664dbf3549d206f0c513f43b9f3774bc8367cf33cd4b3b1d58c44f10efb5921ac1941bc3cd8d54d9535144adcb67e2503f0d2b7bb17e090b1a8ff588b23d735790fcb13e653e3076117dea5a9c688c87ac382008c9dfc38b0576e8d5b2f0156e2c3286f2a0edc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31641acde3c1bff546141a6a73e68feb800adb7af105097e92211601fce8e162900eba034e14e9a73d7cd325156d856e76da6da680c5ea0c39b13dafb834ae2808e8d382c08d70cd3209b176e486c16aec0319442bf6350ebcbf884e86b62e945e3717632c4b17b8b34ab775f89db6fda090d85cc25117f8a8cb65fee4e23718;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb328acb3f478a4b8d7a8e752d234ae1349c94518655efd68c6effb4464bf8e4327f75b0c370d031bedc1ada8094405aa1610d378fef4d5cb4e6cd71bf8dc4263283479f5026024089105e1a753379a204c20c83c036dd2ec218a97f67ed11729375f93c7f26c6a5c9996f139c119d5feef011e62fb413acaf31dd3e250d46db1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h467ba653a1a3192f0c53df9f07eb5f2df0d9e284f0be0463b5431cbf9cbb75a0f78fbd1dd25f47efaf25bb192caa4151cf9814858610d8cf30a3559e0f927eb830e1a07e88a957c47a747edbfc1c55151a63af7a353491f202744b2eff31eddd9f135c75e08a3b6bf1fa1e4f5ca632e0a022111e4e65dbf65629e58bdb504cd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h101e8482f8262ec1fcddc66ec8e4dfdeacfd1cf91de4b6eae2b8be2fab68dd3e35a80769f22583487edb0f6eebba0d1f229b5a30c5a79c0d186c77ebda522eb5719ba0f19603de815e37ae7c0c6b95d210fa6654ea5f8710e003ef7dfad031334e62d6a28875ef4a8d2432f1bc29dc494ec0a2b0319c6f2900dee7fbb2127f4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebd4dd4d873c6288ed5593743d1c578802fab5874a7290691cdca6db5dd2c23103dd3c5724546f6abaa7ce229c6907c9e3dacfd7b51bc08d66a0f644a0379ec762f0186837f87871295fd4ca8a7e6241bd976ef640b77cf87e61098abb26de2c2d27186dec121ef50549cc1b8406a7cf5ebb5d899f303a20023a61f3d633714a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88c0ed89bc66af512baabaf66a80f6daff4eae533e04c7853b46d4f1aa64a1b090d0086c1b5a7c8d0ae808ce1177bb10bcaab3f4cd16fe09f42f4eaa3da450ad6f454bc054ec2354429023d0e14da1fbe21cc19a4a242469a6179922a14c297e51140ad989e6b266a9db67e45fea057d0a0da46de41b0dd4afa70f60aa150f02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cba854fd6662b6f72610f32829f1f13a32bbd1e47e5c65a696a7fd6019619215ef3c3d5c10e8964c4101cef1ad258b98fb32ae2b9d5e0e919aa37f31133fd0ac82eafb79da3757a243ba6dd4b90d41ab6a8bcf09d9251146a17878376bf815c21e8ad15d54e43d6d0b707b2f9b3a04c3bb6ae29e0e90c5007bc92ba803869bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6953be95a2490b9b9de17f948cfa49d776813d8089484753385ac4b6b47e5ed11882ede28ccaddc258fdb92da3a6e95e2652c5830dc60fda2e85158d8ae4c0c3ce6dc6cdf5aed4fa2b347b4117fe269dd167d3d4005ac569db7c0145661196b4df29a1704172a1960a11cec125072ff60e8ef90666d8e0428f070d90382d5e4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7863a8bd26551b18e3199919bd4bfdce8a6dba80db9c1df0337b53fd28d2dc1178feefeda9dc6dcfd8faaa655d4e9b877665cad327e451c3f435325b1d47ee8193d92490e8ff42070596eb8bd63051eceefd1ce1f33034810af38c0229c553fac610fe28970226e2c61826c14cb59a83bc349182464f7101025f6c6225839abc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf249f3dae2d151cac62872cdce21395883f5f5be38d6c3b9866018eb1906f4b25758bbb5dc1f34774db54a42dd7976f366d65cd75975a387f78547f0796eeafd5d0263115399f301c80fa68699a7042de65e9dedf2ba5c66e71d37e529c1aca3a8d0bf5c0c17a9054cc192441dd03bb82afff6cf1a9dd7c0aedcd47293277391;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f2b117b24e61564bde60e7505bd3f11add20ff9b2abb540ec711dbb10225442ee6753e1d339dcf77e2954d4fb5da5efccc4153759f6201502bb7c2574988eb3355d3dbd9944543ac570a03ca9cf45056d8702722abd14ecd27f12e8aaf2fb1c44345b8438763b8ae1e58849b75109fd97fdec63a42bba2e6860db89d7d0cb38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab36a424946379cb7ecf71e271333db169ec1e4df4a0f41292f4d069d37a8cc1be3171208920da5af77ba6a8b834130c6a3f4022e5081857d51e2dee96b28f6675c131a74873cb1f56de224951f738ec7d53a5191499b1ff9164b7d2b7b9dab966b3a15b129aa3ff1ca14dd0e212d1dff675e13b64f394756bf677b623c9f504;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h473e975438a0184ef45d2216d08622942a3d056519beead5eb88ae7b4a3bb58b6fa050e8f6563aeaa00232a6809b3d5ab8eb5c372b05ebb897ffa7e7e74517a9b444c98920e3bfcc30599c0fedfa9dbe563d654601791eb9a2e9df0331ed159e99648fb79609458317648a0d8826f763cf25dc3be362a47865c5af0b167eb3aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97d9db0a0a25149763bff4873cf2412eb96170eff80860fb96794330ffa2889f759acad26ea899b5af67f4b1d0582009003832d2444a46e78beecbbb78a082a76a584dd336bbba942f6d33e3039a64bed83be934fbe87d5ae1f48902772fdf90dcd7f4bcb7f656e13951eaa00b153bf3d32069a156d35dd28b62633d2a91293e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2862810201f29ce08db92a9273b143b040c261b23dbea4ca6a202eb2831089720817ec6310db3c932aa026158382319a1732565f677855820d9fa8a4236e3f716762e2b250c960b8e905babf7525d0dc570f0d6125576b4abac1cbaa0745720aaaaa72272884a41d0c79ff21dd984e1332c1726b24612753be7ed62a8540f1c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he01623ab8af517652a95ee0896664495901beb164221eda1127cceb71680471904a79d6762e2c16fe6978acb101a5900d3d85fa26e69ff0c3ba23d7cbc458ff74a032929f5355a98aeadfd2e431f8be1c1e5b75ac842cb029313d34de49f83658af2248342e1bdefecd40a563f747f00985c5a51df28246486cd8cc2efc0896d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d3af8492afa7875f8d59aa262d943363b31817019e30d9aa00ff598c2378216772754129f7d3b33c5d34e72d841bd28129e277b92c8e51048b39c1868c1023d898844ba4f5384f47183976f88f8e6d9313e64c07d6b84cccbfa0c353beff5971931485c4fd71bbec1e59fba6f33a9a9f2c9a3bd6dbc497b4a6933af685362e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h588adf5c935097beb277123bb583bde9d090a5f79932a93d2fe3b974db529a660937178fb6982ddb8a0ba7c05b55f8eadf9c2dff819b547164c53a64a2120b429beb3cf14a67568c3818eccfe7c6fcf23784b5e388711cc1e13f88b5614a117c1360bad45102237e07762a18b3b9cd8e94fb37f314875ad3aea283b7789b6e96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8221f51d3c9870a247a4d0717d789fb5b823b1c0d12c6e004e4148e1b7f4f6c00e12ab84e3b80e54f19c5f236b63769309d39b439d6b5a81488bb68c344fb1d07275cddf5f942935d0bbef5d01aa0f471ae0a126f49a0e61f851e1d115d6460e3e541c8f89cbf8830e53c5adf61dc9690726b2553c45154d63c115c32b3df02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9a75089825f3095331761b6aafd4cab89e29b9ecc3ac25d759941ab70b5d173a56784fc10d32b709fd1def8cdad03da46aad217d21ae9f3f49df45c88d6b18c997d70d6959268f6eded4363c3970b61a9886ded3eaeb347c313839c11a74482d5ffdafff24c48c1fecc512cbc3e64f97d4edb1600d00c9ab5024abbdb528b2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4909dd4b07730d2faf070177972c1ed66d0b06e76e0926fae1b52f2616129a0cf0ea991dbb10d7109465d24d566bcf50fa7ecfafa6367c4d225f5ca9e5362f722fcbccfeb7ca444c2c52ad990405321bcf9fa6b9d3f01ef585b501b1f91fe57c45fdb0bde1569962320a83b8976195191be7a3f7e2764e66afab15215d698b8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f0e9deaa69e1d9981cf5a7b558adaf00c90ded1ed76be41351a1040f41152185f547a506242e8ff9f004320aa4891e15acd606da314dac076b4cf53e0c5662be85105d9e4eee0a2fa83e46540031df1040541cf27797e5536e09379def55470f806c1fc93a1422a28fca7c729d654ba84c0dd0ef4d09cdf36a995b3a0cff11d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82504217170165b57f56b54d6d9b3b966bd943ef392d384bef59a99920621a675b43159180d764ff4327f30e384930858982c2c8c8d59d68a4c0fcf5237fa021fe59dfba520869a2ad2aa9d2d044758e2acc16d686c6b25347fbab4695e38cde6af7741c1d9440f1a056e964667c5672f22fa85088c3be3f59cd365ca611f042;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43b54a1cf482fe310471c8f93d0677708ba71ef335af93b3b6daeaf18e42569a920f0a66a02c023eece9dac00f3893f3ae63cf3bfecf8d0cac2cda569adaa1d19d9616b2d2dfb616e139ff2e45a421b0333fc822cec4fc99cc050cf032c28716080c1dd820d3b5f84cbe01aeef14631e8aae7f1a4fe12ef3a1a7d4b63570604b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29160c9be8e42b69dfe1114960e6f2ddde97cccf213d0995b33fd45a4afb4be8e570be98070f5c96ec132381c50f63d9c1a55827607cd5ccbae2b3af8dab1fe51e9826feed6e94f9f088ae4e37c7efc70e6ddced30e35ecfe1ebc58c587010937eac48cdd0feea005a66142643be014649911c348d07d7a7c7248bb87c063876;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b2b584d696843c4b366ad7a02c59d755d3f3973ef8c98e25e6c9e6f8c66ec7b48fd9d131949eb163f71bd594075589baca88e5d6d56d20c79969ef0389e171c0e5a99e6f430de9ac10d54b3c00ae567f6d8c6b29ca67fb6739f4c5e7cf7de357d2b2c25160a2c4f6ea57d54d61cb4c5302ed1567731e0b5c88d86eb91a32014;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac66646fc06b61faec6fa3cc7ea051751c48ab05042fecd2f745a791171d337fab920ef492eef98434e6c10874b567123ad7e279c5ab76aa3aacc57ec8bef4b82218272d36ee5436193a7b817483c48a7762babc94e241285d7e16f2ac5ca5903b34ec6a32434a0d076199caad8f2444234d1dc837508fc7b915258c9da085b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8469cdbd48931a2db87ef73dead0dffdf1958e9a4019a6866ade7c0555b8e871f8fd24ae336a10c6161371b0392895ade9f10852b0902922555cbcb578232f368742296794550fe7278f244361806060d4731250ed3a1ece47bc9bc2e20aab51b4eb87115cdad522b12ba749d975e10312933f98cdc05fbc11a8115075e91328;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc34ee5b46a2df997e0b3f6e0c2802555d74a9824ee0dc1f3d56bd8120a9aa5703c2298097070cfeaadf68ac504751e37cb437c4ce77e07f4920c7c11037d2109ed08b6995a8ad7b187f9735161d86049b0a18187635025544d6e25462aa8a5867096eec92987cb7704d937520942d708c8e143af0e090d3c6bb2c5837a32a1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1260ae303182708b998d4cfd80fcc5fa12cf6fd082c4b20173027d39ca59af118a2c82afe98c9b164ec35b2ea82bf8d13c712ede0be5170fc7833e37b040bf5b07e5d206b2b4a602be31f4b872fade1609897d1a8bc0841442b0ba434fc6b6fcd9598e35a647ec1c2dc4f17b2f6b1954f54d3719518ceb2cb4577842ea52f0a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9110eaa55d752299a9ef9f30e7d8b9684994732e1920dfe6f776a035472b13dc8eb47b81706101787c8737bf9e29a23094537be623cf603b5de08a5a4a82a36287b787eb3a435079c6a06597e50b44d2c8d3504f5041b48d1432bd4db52da139ebf64089a266190d50acb86ac37e97c20202805925b707d43dba7fbdaf8c3011;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d9a29667ab07a50eb2c905d27adc9d97eff2789baabc8e77e2701e6aa5e4edff30f24a436ceb152466514c8bcf7e9ce7f39048440c358cd380224071236a44625e895d8f4b54b9e1dfffb8168eec52351ca910ed671a22e112bb907baafeecff14e8e788d5bfca8e971775220d91cc457cb51ba4acd7fc92f0986265378c3af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc69e755ff3d20af91cc77e259cff67052cfa3c2c5420cc5d03ac0a2a5d388addd10ae30411154b3a1a453b1b31966528d0856631dd4e4c86caea3aaafecc6d2a679e9d8d4935c7c7096429ac42b4aa847d956911e0180d689f29a0086189e1d23d58c7b3ac223ed631f49777a4073afcd343d27b9296ff247d078eb73479e116;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb07e010e5c54cc452e9ea5605d5f9d327e9bcd16139b18c6d037353b636c7b816132b983b4933f548c0636b2fea36dd9fe9f1401bf6bc3fd7a1103d90e7f1095aedb27b045dac7a32aed483f713ec5bd934c17314819acb9f9d28e9c5388a659a847858e17264076d41070dd179cde148255d43a157892ee3c33a8f4718a6fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2918ff1c299fb5ff0ca78ea40a1e384c0c4a5ca272b9d976054b2ee0d6ee19e047c92c69a8ffc4909f00f7ae1afc60ffbff5c426264a0c4f6a69145af03a7dd97548ebdfc8b29779866485df15d8d32065cb57acfa7589ecc531d1d9684db68c0483ca9ca17254c72a8c1a97c337a615c0ace839d74e2f8157fc5e168661800;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28a49f1d67a57b64e5c2ee4a361676fee2899f229a757c5d5f7c71b6abd8a39545c169638a42e331f1119a8f7a91b1ef50a2eada21710e1e0cfefd8d35760d1ea9ebacf1f0a63707c928424cf46555569a3d33e93afc5dd9d27851d2901a1990d2dcbd8a39ed0aef44d48094aba296751d5d5b528e2f4c82f8467c77f6c07e43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h213bd895e3c2c80beaacd5fe4a6d0886e03c37c47be34ebc7eefa7b22947126ef4a595b10b6fe06f1482704ec131f808fe6df20f36c4fc798f42ca06adb79f349e69ccf44538524b5e25d547603453e97c66aad9cbe03a35354ff50f2c52ef8d42e173dfeefa54a415f6fe120df14d71d1bdf92bd7a898a0f0e864daf28b316c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf37dca757a7a99388e0c622466e4023ff9dbbabf99e8e2160089311f5f1b7adfaa46ca29022b228a4fc6e1dcafb229a24dd9eabc6396ce61c6080b7ca55f4d5a32cfa5815872704ae45e5077aaffb7ec1c41e61e3ea3a20d861eb54f0c2923280d7e1854d1445a1bbbb858caf5e731bc700871f56dbf39ebabc1e7b8bb0bde8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dfed8f09696c6a07c3730af0b31826cc2039f38c332abc24c8830195f8c8b04c8790da8edf6437f6052fe826a717e0bafd1a616413131ba3926d92df619e2364e3dcac10f9be4eb947c9b498957684909585bb806265c1903e0f0fa81ceb3250b5c486e1b65b35cc48f23ead09d00ff118a79c11eb2b4e4f68eddf1eb9d5529;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1552a60a5fdd0e74171a3a106caa184a7972da36154d631ea529bd9bc6c48c905c2d02dc4dfdb41612c83956d8d94b8a4df0f4844dcfc363f8d28ffe33cb36264d948c95faefdaed49baa1029386a204881d430ce4a9acd68be2fad82966c400e813dee3aa8e8f20304f7eb930245b392688b9c749e903a8ab5866b33346e2e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfae5218c5eb24b01253c701f9826688cf6b9890f145523b35802b54186e2475d8c9d2e40f153c269bc72bc0751441a3ea607ab3f72d14aaf2d65cbd1b263b1ae607a14b5de88e37645c92b5cd95b41162b5b209a5e512082e01bec7ceb4dae776de296a56e6961b80f500300b557a57334eded805c8a5d74dafef46a853406bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cad6d1b2d0f9428269504411e7859f5dbe12c5f61d6d9a33ddf33ea2f0f8bf9ae8f364ec4fc0e50a5cf9a81d838f2b333607429f596677d2176a2a6b8c0e8bdb1696665b48fb47da4d339fa2749a5b3245b3238c211ad36240e06085703f2d31bbf691e4abb0d4251faf7328920844bb3b780219d8d5d4250a768c7047e84d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ceb57bbb004d99a6d80e0c39a7861740fbcb55a2b4b02f76de977b3af401e016d940f2afd1fce8da48ee263a9f83a101f867bebd6dd0741618653b13c47562d3398fa33139908d9cf8ab80d4ff60616538779a214862ab4e7ee2f55d086b3fde9ba012e72aadda5273a0fb7bf5f461016e0d60cb67124b18fd3d54e2b8398b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0c3d2b513b80d6cd72d01343f5ebb6ad09c92d861e6fbaaafe9b56a86759c668f1d3c081ec7560a1d5ecefe8034b3b35acdfee3420bb01bd42d2aef82406edc2ea51857ab59e7fa40fef2e9dc0cec8e7a9068b567c29fc658b53985ab1a7b96d59a8324de65e27aab2c02a6663710423c3d82bddebec4caf77547bfbe8e7c69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82b63b9daacf7e786cf420c0243224f7f87142b22b2c67e0864dc98ee5ecfdc3da5a52f549f4b86cec9e6975e27f5155c80759d2364d0a9173789928b77f5b6957aa4365ebef3d95425248bb57b8ecbeff302a7632e645d9eee70c8a41dad979e7e5ab6788d74741516ac4edadb49f154fb6efca473300922b4874353bab9375;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb028585f51c5b93116c684feb281db891fdfbe50ae7457371cae76f107e4e05ecd4047cfa1fd093f4179c6c0047ccb71799962cbdc8dbc4a5a4123b41399cc039dbda78fd1d74276297bc28db095f8a7e0856c490c591d469f9e681c0f300584393e0964efa406ec1786af380469d7b5dfcb2e584cf54d075bd79cb04a6422ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h219b98ea6cf6f5f4676d415cf5d24e5e61acfbf3c618dcdfe04543ab149836a4835216191da24da5c058ba5a3b011cb3a9d9d75d2f6129bf03eaf0d612702a9893a9f0d7dbbb6811679c0d4d1a93a0b74f3db353f0827d7fd8050981036a2b6876f01d10778a3fd2fd0b0216586f21fa6adb5f18f5c2345fded7e65f0d3bd867;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a88a52c649b0084dc266c0d1eb75f89a7ed3e3207807a65218d7e2e20c6ce51a0b77a3d901dec33a883cc514199a5fa8ef232834a7dc737c41c3e886892d50d307f24880715d6352fba68802b26c0e3d4f89ab634fb8f1a81c24a8bade7a1161855f4deb97bf3676492c46109e37537b08d1e5b660325c5347be441e23a9eb4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'head5e2851c7606f9299230a1169461de1d700d64c17652fdde9753d0fec60f2391c3b971ee095b8bd48bb36d6c24fba6eb288072c0a3da5a685be52d7462ff76afe5ecc6ea6ab101368e50dec05e0901f329ddf6f7591e3fb514b97dfc801a4725839730558a06d1f033c471b6b619c91fb39214820828fb672221155e0ba047;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde5bdc4bd8711b715448beb1cbdc8caf84fe9a36796caf46e18393c2cec9180274143eab006cd317572ba1030957223e70e7882c8615c249b03f5cd348dd597b2f1c60bd23f62d0932b5ab64a151dea750cd0ae47e0b0921410b7720458daccb2ad93a7162628488b10470320496a8cbf32a632958d22e05018e3936e0813923;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5cd641e1f526138b86cb62568a53fe6ee41fe67904ee3adba49fadb7a536fcd7412a1c35f2a8dfe09d36c2fd1886b47ebbdb8bc3679fb1864c05f444314ab32eee7625d0c45224ee662048928788084289348f20dc67ebb091011e5ae9293975932dd3345a4179efff28900b07d172f2f532f5e48979849c96559513f80634;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b3595b22763e86ae6a92b66113b4bbb739f50062b7e64d7fccf45488ef4d8b2c3b4784ba9aa169f6e017bf25a346843382699f96a52de9c3910b5a2d46ec498d342ba085652e9aeffb2ffac3230783985c1ccc85dcb939729fb879da223ec7f415a427ec4b06e7539b36d0d4019e56f522c66140ee32af836cc451c62486aca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb570d018992b1a812721c4eb03e733b2dca2f178edb589e82ca9e15d8a560ab61689adcfb629f912a575b8b68bff25781bd7073eefc49a4a677cff8f6634c19dafece247860055a6cfdfd6a8f2b8e54a7f6c338d5b8da28f62cf6f421c1fe4b93ec441a55f66e7a25c3780d26f770af58cdb8f5d6bd1932f1921e3ef7385aa2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ff95f3495998248c3b5c12279d5bb15b33cade091f6195fbe8de5fe6b1c88e53da74954f0195a85ac86c7a944c65d28f2ebe8ec162e2d4a0bce836b9704229879cf5173b622fa5efaa8e53e63b786bb7db7968dfe9fc9c68f4b8e042b350b27e15f06ad92d329eb470cfcccd723b1fc8c557f899161f8cade414f7f13561c18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e7989bcf289202bd8b11be9390dbdfcc969299e5ecaddacbed99ef57f13474729fde4b95ac440ef7059c5c1b73492f0abe2a482373cb3c548d518f94f841faa5e5b7e8b59930a871b6b307f3ea858dd22f28a96b7d3fbee6fbaf66beeb61773a411fdb90178948d1fdc7d3cfe04fbce1ff00d15a8723f730c8f60a721181ac6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a471920c8e2a7312152736a941de8ece45c2cc72a95b70660e090723ef66077ec15ff367378f172358feffbf0ee1a7a23254de2be87706c91f7e758eea855c0ad896f81931137e5c9c62e6ca5024cb061c4c86315b28cab4ba6c210347a96a3440bb84e8ef9bb57e52412088541426e82d4c53488dfac842b0b7c9d800a27e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h379567327ec51839114dfa5c3c5dc3599ca583fbb413f3d83a402634984458c5a982a2532ee52fcb3adc9ed95d83b98bb86313aca68a0a2cf3a5f7cfbc8d1aad5f69b2d0591e0276ed9afcea145bbfb1ca58f3c9a7d9ff2d9860ae727d5fd80a3b1e3ab9de8cdd3f13e5ef33cdbb8cbe00a730b208fa4a786db2371d89f1a57a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17db762ef526b4fd49135a72ae807764ce69e5c289fb4d44f5896f19607b6e211d25abf93a2822cfa5c02ebd3114bbcbeb79ad4d5f84334d942ce0d1270697acd3f4a9f72d09aba9404f2376c6ef13a94335bdea0112a236ded99a850d15348bb0789bcdab4823a92621c36af62c849bad15e38a614247fabbfe5c2c5281d513;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94892dfc9f3b6b6be1b38d317301204ce5f59e622c56a4a3663c7fa0e2ddbe70a506d41ce816ba68effb0ee50c33405796f14c9169e00a1b8f920b58629d9613ceeb99db231302a671da877425dd93bbb7c6d566a35f540ca094b79cd969615a43c55a48f85f34411ffb3c36e9a61700ab91df422a66d87863e02140b0d1627d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a09826423a7090f855e5e34b9bd0ddacdbf3de3aa5918a99b5c55f056e1e1d273505081f9de7a92d0d177b0970e5b55eca3609be63b22963775d9731aa63c751d92d9d5dce7dbda8bfac0aa3c310f3644baec6f8389b9ff95bad1bb5a3bf59cf9679bd998748f141fdcdb170ba65719752ee78704af5704b00038dc78637e77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h646997e152001d398a0488a129355d2a44e510d815b09ebdc1b7a34d65e0fac5d74ffa782e3ee2577b7662cd0ac2b56a8a33a76c1500f741dd880bb5f3f29cf0217bd75bac84bfe25e7ef8cad1f5ecbb46c1129fbcc9499e8af39510c37ebd62ce29bd40ff22e768e5572f0e649321c266bcd98c44d2a044432be7b9e000d06d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22889c04d8e50a2c7a5c3a682652a474189b978c3a34c8d67e447a4e619be1a872887d289bd85c4dd24ce0ba962e7867ad79a2b52a1704c0b8f4c6a74992e9197d2235412dff3d19fd495b4f6ced9f8341c924dbc94c080d3e2fd832986c7de95d2771229ee25e1d03602e1f1447eb0f009d219305dedd35345cbf717ff495dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc55dabcbb8bcdd46c8d7eb3d7d0ee3668176c6764f508c64605f8f8857346d741bb98a0eb721a75e611d0921a1057fb612eb51bfb0acb5730cafcddaca8113615e19b6917f17e4efe263d4abf94dd08423512fa193c49490a746b148e05d41331c91f7e71d79114f5f87e08af8958b8e774cb4bd23e6608250f19dba3d66b059;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b3bd1c11e034359e165ff4d31acdc3efc5e4e6802eb028417fc8972848cddd866d29e633a052fd27f092602d4361a1c8ae504bab0dd28e7e61bc48713219e3bfdfb3a4d65d3a5b3f1be80e7c701c5f3d51fd65d78001453e947fe3500e7e475f545eab8873a628c15e023624aa01472037f15b5d0dcb42e52594e1d083a244d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29cbfb2dcbc222bce3938f2e99df515348b9e8e091a1328f18c97c30869f11f33ae499f698b5dd1074d364847b8f74b315fc55543fa094bb8260c9d275ac6062b2b765f9e8f45c87ca05bae4bd4d96c5eb938ca405927520f6124fb7800f60a7127f1fd7b2bc889b65fdefb512ec3834cddd5556e76d71fcdca608ca8f3bcf71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d16d7f5bd5b5232d140331c9729195d5974c78a9b85aa31fa956c2a45a241f52a6a384ba25f9bc0fa70d5c4d89711a0f6bf54db2bd21aa36fb95a8020513fbdc13e3c52d326d995b69189cf770a16f6cee9aa303f24751c91ef0a4a3bab84e3e8f9adfc3579c54fbb18c6e2f57cac5ad100b3f76a5d925c6974cb9501a52fa6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75316c69a80ca9acc5515ebe49e1510581e589921be951e39f65cc06de125d910c297b68a269b63e5c14e013402ab7b519c01677009bb92c942432d698902cccbaf2a300b78326947f7a9af49dec86ef1ef42fb9f5a1b21a41c71b3828125c4ce522b5c3eac1a9e7db23a900594513ce81cbae03b874873e25f6c1732b28ab98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h777514f0b2d47fdc7279d3bb58828b64c637b04f44e9fb2575397cec4c32620085faf1ed5fd0464fff37a0f3d836384f757bf7e16aaed236bdd32d185a927727971cbdb5e53d16d2af8d5fa01cb66c4354a0efcb813f3db796364c094471c5f128dfdd3f34ea88d382fec0b93d128b3740c8065cb1bdfed8c1730f23793143ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e7a6be64903b4fb80302b6f91d41d2faf3ae6036ac253592fafd5aebcd84e0cd2cdd41aed361ce6ee0fe1cae4ebf694eec3937dec409f1bcc5a36f54e6e92dbd1ab6056e187deb9db8a6a3d22f9f1200b68066e6ee69a94ff6319d0fc84e14e4f2cc50377c471a60b0275e3d09c51ef252eab2c8737e723e307451d9f72dc38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee1536dcd541660993e0a7d2fbcbc30c32edc0e35b2bd23b644a025c3dfb2f0846eab0a16f88fb9470bc3d6bd8a4e3282e2262b790723feaeb1c924444788d753c0894ebb2477a27303ecb34a0c495980b512b82101a02e0884da5e6d5bc6e520e265b33dd402364a43713321e3ab2b81e6ff4726a1c11fb4041b0e6d2ee9a21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha987951c49c57572b89b8fba6a38f55d4e1bf3d845cbcd97445fa25c3128e48208f5cd5b17a312cdf4037243a8ed9f18142a6c17ac9216f38b122e637cb3c59b1675f10b39cffbf6ee212471c43067c46caf62aaca6f92520b4df5065122e8f00040e5bdb6f78dbd73647e01ccd444f62d77b5aa532f97a4240ccb6836ae5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6de5a678ab3253ce427c10cca947808f7926892afba8ab47e9e282c16fc2f0fdf196c10684ca5ded2968918cdcf61d5758e04303a42e1f7380d3990320b9b6c4067df1e9e08f84e1f4de35cea4de2df825515e8da9003e8c56e41e992b10de311f0b2302e359b6abe09a8ebe796d1073c45c86c97bc1586d2270970d55fc3e99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5afedb360530cb629766f6e772521544300099e4a150c7e858e756c8055d49955651046f0202b9eaebfacb0527613dc5728b8c2ff2c244beb44fece524dfb8de093a3d54873e57dc9efac063495fd6589e81b547c7f22e5fd10b52cbc9c941cb00f95a31f5b8021727a706628cd6c82fb4a4bbda10c1c05ee823a668bf85a45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd200cac932f3f105f6ccf4172d88a036b959b278ba292e6f6634f59f1b86d4b5878fb453ee771f294f708b6826530ef01786d8ec8b59b826a44dfd8d4da6647402393b3c94c6cf536df0edc2936b3dcc16c09e938097a373d5d3b5ae8a649ed173a43f985222c15567323cf414ac34315d068a7bcb08d20d3a8cec06f89e8c7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34abb610605162975bb0f33960a46abbfb34c4d26bb94dd00a9b369dfa0c03a935e274e17e6228acfcd901841e0a1893f76ff3d8f6d80fd2398ac7a9ffb046544a1ab080941231f356c8ea11e5181e40f4f9829baac12688824b4b895a8ba100c45d3217001f9d2491fcd07c43fc9620deff095c55caa78c9818f192f982f438;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd377071cf04a5aa2fe0bb5c8fe8e8301049332622b8fc5cdeb644949902b06f767cccbefd38ff8982517f6fa564d496a56ad2baa800b6dfda3de5fc19c737ebe00c2e6ca317c8c4f0a74256a0cf0b9264e540dba55a56608959b53db67a51eb6b722cf1cde5612b0136121831145e6cb272e4bf6da14c9d9cbb946b2f9ded2fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ec95dcf1e29636d1c121ffc10fbe75e9bb74fc816fd9334586095876ecc5af5821724cd82a0e3ede6d6035c6a127ea720de45eb883af68430c5198554d07377e4008dfb6d39899a7366188e4b9524913bc9eecb8abd5421f2aa8fdab8b8aa7a258458dadd785d1f8688c60587ec39e5d52065ed7807ad27c97f0f48e9bcea3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc91d69a1cb1080d70c7acd6f3bf6eff8db1ea017f2805d3a552838174675b8fb559fb2bac561a089b1da2aeecf542afeebf1892ac3ce1c50b15ca2e3ff0320c5b71a0f5b7eeca243dcaa22443b0c58f0f979e1725cda4f71ddc7e979e1ba99fa238c58a838685a98c28f6dbf5e46c816ee71c4246f899093748af95099ec6617;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c639a54147cc548c3a0e2106e851a8f4cadac8ac41e439371e5e390ed59953adc8c4109454989a0727e888b0a822fc09e332fed56d2119bafa62b5085da207869defdb7a4e052100ff59419a9c26ebc896b7ecb9cc33e34660a397d02f31270e780934783e062b0a5ad62dd111a88c01c9197e80902230806ff4a58b3acb872;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5aaccbe7d869cc89ae24e042038132cf4dc2eca89079b6cd141c36bc72ac5458302f169605cab8de41094f65b849d486c25e448dbfca1910fba21356a641d7ee54fc2742b5b35ec138cfcad3e7393d7bd826e84b9acbc5ed3d1fde59954d049cdd50200906f7eaccd3503bd408c418b66237571dd64c4de14bfa66c61bc6d58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefa254d13a87ca0288b0dd58b746efb092f56c51c71db6c1b84825d3bf2d6cdb548ac58950deaadc0acdb8486cef5ce03cf64778f21dc25f85d2e26bea9af5d8b52d45cc45b204e257315b1f744ed6881a13d4d3339298cd1631ef7371a328b2985d41b16bb1fab977d65e006dc347de154688bd6f54f9a5345e44412a5f3e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca705bac69774907ec1b35c3ebe2e48c919c448379613160a561266bd067ee16172b2c5968e117375919b927e274f5e7ab1c85fbf1db4f7587df4680d628ee49dc3395bdf7db10ff2f37db74dcff9c7bca82a4caa45efd8459f5be1aa238b03d25a11363a760f3ee80e63e4179d980358a8dbd0c9020bbdc72ac65d01fc084af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d48455d76c15ddfc7b61c4eedb32bdcfe0cea7a495578b5eb890a0a3912ddb64b947f2c113a3b73225bf17b9c576987136d6d28dd2f29b109713d035baf0c3a24e9949870152618da221e5a33db02fe4d045546cc570537e03226ed19a143d0b8ee572257b0f27249051d326d00a323a4288b3aea313a7e3fecbff65bc58ead;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd320ca63042965609a5e0b681e36dc61fe808d109a6117ad2f18bbe16d4cd592fa1beaeccc3a131106b25157535c9c728bc680c91ada0a763a28176b8cb3a77e504de494a9d999294bd1ffe00aad8ecb5d251d37e7c26b7b7a39b01f84017440bd079ebdd60a339c76e420458b449ae9af8ca22790eb412353207aa460961580;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bb98fa500c26e644f4084d38e5643a4f0d24cb4e8cf9e066acaaee8c4287e9291ddb2e9dcdf466a6fed0a6a3dfe6addeaff3f465eb6e1ef3371a429257a2c315a49b0607557aa04ca008565da45f33c5f25ce8daf237b3bba8c016c55d9912863ceaedd169b2e86f91845f03c7f7fbb142078b745b993bd3a9419ced2828252;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb10c5efa63a8b76472036f28e9582be2b88aff8d0d7076b6b5a64f829ee09c607a7bf78fd1b1eaa3818ad3cff6001f22ec472a0650873814f2bebe962e96bc47eaeed9840b58b0960e4ca645392d0ad221018bdedee003a62c61986b20053da8ae8dafcd81a1ff4df46e5b8fa7359399204999ee34ca4a762a256c30b9d3f33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fb676346c1dfdb32bd745e4a7712d29c6541cf10225ee5227d6209a28431ce4b5691571b9e8e75dd76f597c38b4577ef16c6d44d7cabb2e5094ddd40aefa409ecde86832621aff0cf5fb5cc03d68bea33d7fec72337327f3f01e868c43ac8499ff52705e53867c18a818ec3cf32cd678e102d46c19d4c00457855e72afd171a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67a7d44904085d0fef78bbcff53d807019050f857318ab2e793728325629406b0ebc2d491e0315c1b754960c9cde9f812815eadbbce284c78c51ebb7ba94f37af3e1f3e3c1bead44f1afe60fb67f1c5200aa01ebb744bf83346ff2c259c2a9069de403d56530983c39443797ecc39a34fbebd9ad395f82aec196bb678b8092db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bbe3b630e1b235471e5cdd2e2f31ee6a045e46d8fa7e60e9fff8080dc042bc9078aacb05d66ada05f2072d46688f250185602af5b39a238192c12ee6ca0b112bda0ac36a5fc40b1082e4d24cf5a1558fb0dde8c234196a2ec6ebb1538824db78ded2663d88b295fa37d02a805a8d21e1778d7ed85bada67160544246cce6218;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf96f6c51cc63fee4a7c466df3af55edc924c436af46988e7f9cd0c3f672f07ee09f579a9118039eaa3ea4544ecccb7105770ae3288de6b4476ae73e24e8cb90b5efc014af7a8ed557ebd017815c12abefb185b8184bd5fe25b43d848e96bbdc64d4410f5ed5e0859be9cced0ef2429d09e18b5ad34f8e313e306bb450648d71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd44115668b41f66591f5af56a2d1ec1a2f5eef7cc4b668bc0317c0a7cf4325a31d984451e2805b4befb8e9c386d207d6aad14d944713e10340a9ca2f8895e49ec2d543595e249f99e68ea94de506531513a9a4f28dd44011785676b8d233929ce5dbeed9438064f043eab57a3c23cc1081bc35079f03f97b27d646814323195;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0b5edcede15365d185b4b5261a4f73b6b55d2e57d7adfdbad47cab92107499f85b04af8ecf448a1fd7d3cc7f4b5405a850e36ac2b481db2943347b11cf55905c8d59870ec0b344918f19e9694b0020d8f710dc2768d5a33bb1187c1a2c6103d1618083fbee51e02c5dcb469362cafa164be9b0492aa3835a60a2b63f28cfc0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b4bc52ae8f13e2ce8c4d7bb5d6c368a02d0eb0b6b14da42002c1e3961712cc25d2783147151fe448ad5bad93d79f8f8270d8ef2443a1b9e42e7419130676ea3a1fa7a6417d1458d7da74ddfafd86c76b060be20ff0e7f818e405ce848799a16d3c4adbc2ce6973865b01e69630c9c62f26e97d2a0474c747c0c6f2ad1a43a33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5809e125f7698e522845a453323c003ba9db8ad5676b2a513385c9886e4681d748dd759942dd4e4b2efbc4062c2d06d38ceeabaf480bd01dc602388ab3fae7a158fbe4bb8eb4de2b9a310a13c6f7c5c3e8ce294835fcdd7e94ae082cd4e65006d8a18321dcd9c4d06f0535f492c228609d196ab6b196a4276681f84dc832061e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9682abd7da0b879781955aec42044de56619955dfff8900033df0b7accbd2393b9364816bb6e8e982753e14894487f5593245e4f8f7fc167b65eb80815c06604c97db4783831c2292ca31b71b03c9acda7cd6a073273cc7210bf7aab6dbb42b24c78d0e9f65b8f6c8d00478b313bec8f5cdceafafaf01b7262ec04547d465b7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b02882f84e3b364ccdeedb12b076ade2c4e6815b890025b4f62d524a7941082ba9d37100cb697afd656276e75b9eb03d63d84971fa9300a35ae9703926b56f49f71eaee9fdb04c0f654b32e631f621416ba66d27a290bc0a679cb34fc0757746f2f86aa8c18de0ca73c0e5407d229d2896aa92fb092a72d32eb60a589cefd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e1c75cabe01be332904315c7091c71694e58c354a33e2dffba0e665cf3a8cd2598771a515f835ed8090db2cbc3b07ba4364331493461e7499ff06a36c2853974b85e6bf90647ca6267b6dc752cd1a3bfc0b87c369c72edefad2a40aff63465f2bdc69a906cdcd049869115b21dae66912dd5c1215cc7978dacf7602500ab869;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41d6e42e433ae72a963fc93ce354122fca54865fe2ae00a577f3b04a518b59b80d93ed6b9b231a2405939b49dda2875f740787474b17986bd6a6ab2bd6f853017006df0335b968fef1355c77c2b59cf9a441232e5caa493d71a309741c43becbf5cdd70b1170ae3d6e8c5a1cbdaf704a5a132f33744f65958511d06ded9ca5c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60a988179bbda2d5fe64b2d854644f94b89f9af8d8b9ea2d13ce8edc5c8b46abc783eeef8b80160382a719fd6e9295c97391cbb107cfdb11a79783ea0ced3d4f23b50059cc64b4e874fe01c542efe98a1d78b1b021808ee7a36bfb692d8d1f4327e5a6356d965fbb63430e92030ecea2e7e0fd6588b9ab9020553d1a12d7539a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha58ff659e274287604dd7cae1482daffabda7ea561ef213250263cef70d41183f2926b4d29e21a5e2f362cb4e45f0d3e9e1a5b80e6fab6406f867cdd9449afbe47d825346e81382c86d03b06269ac3b86a0c29e7f4742a35903bdbe37c9e083a9fbb66de43a5b7dfb45e4fdf800050d47e059615650756d3149d2adbfd569e1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf81a2c3fb7a308d9fc821e5b0341ac7c567a5c30c850d1b0f12510d2057271e8e55c54e1ec53bd784d12e9efd74b34b1fdfc08de91861dd0953fe0c80843351734dc86f5123c04ca22ac35c66847c9588b2bca0afd712188766e550d47a5b0321c3960eca55bd6300904e9507ece2736861f00172a774361a987669070587490;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe2e3524afae25bb69f5233fe5c0ce9143f49507367a7ca5773110e442eabcae31b793a656bedb56188bab4596a34acde03a03edc0fa5d6f39794014a8822878dfb649e24b4a492f549a495c345c6be992192416c7b67c1075734c90fa754d3a19d0751f22511bda590033a02e2ced4d829ec3810da8d42a0f9a09230818118;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdc52c1d24da5e30a8288d37409d504d3ba75436f01b835600a619ee08dcc0def03573958e426de1923320e2e7599cd116a2871333b5be1723113df93d558c6d3e6ed2eb9f0b4fc1800c4a2b066faf8a491ac743af3894f3b6fd9833a2d69558b5cb7dea1a3c81f0b39ee3683b9f49398bc0ee304e5eeeb370b38c6598bfd5d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41e1fda28c0555325babf241bcfb665e78aa0e9c872ed8fbd86b654a53176d0c0530afa4690f15263e79c0dcc7cefef8ed4f8e331fbf579df329c3c5c5c3d06e04953e2b8a75c5641e82fd3a7c42ee7e3e42111ddb5fa13a07290cb66114a865d0c85009ab37c7953a260a75a31988af4d229964783c37455b990302bbdf20c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h616bc296f352e535d67089e6a687fcacc7daf2152877414d9d5b593245ae0c713f977fa00a08cd4ee8ed9a975754b36f7cdf5ebd9f3b6aecc45497364460e71098a67d49331e436ca25c3cd893b448298a4fa2a89efe307ca66b91c7b1501d3b62f1b4fe447e197842e7493609c88480e6576597f9c1dac2665e8749b8ec6bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4e82d1bf36a5768ec479bd5afe6db4ee888963e4add8abf1d9e807b0e71974407e4ddd20b2235bb78e847b65b964bac214391e991d2c23b2c10f144309f21d3fa12a0efd983fbf99a887699b3a903c861495c01991b02d9a74383f5a5fbf3ce5a4559a890f98fe7d93ac26b94fa4cbe9aaac7e1894371513485ca3544057331;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h106ad34d40b7c5ed37493827a076c3c1e44242de6207f83a7b704d85f6ca490342741554d2710560e16bf598a979faf52b62b6d111da0ca2ce6f92d689b9d35cc57b7bf643600400f923da880e07ef4f967e3048164b04530ddb45c93dc2ca2dbb9e1fa0fa43e6758a372dbbb4bdbfdcb9aced8738cf11b0157d6d525b7fcbc4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h602efe62061a1efba0ad1fd596be545eb1f57b2dff5c167419a28fc0e3eae3d5c37f17002e4683248fcf9c1f89837d1a0db77365fd04fcb6984927d98ad0069e60ce8df1b7f8edca5b844bea52108c79293cad429eda5ee04a484817277b2791c9557341efb6b003425ea09a851264e529f59b210c60b482f95418eb426a77f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ac69376877ceb22b280a5678feafc6fc4730c869a433d9eae7229487cf474c9d91dc7a8b39146976badb453dee9919f4d5f20374ad8304ea0f5250ace080d9705abba5e472866aa8f0026f3ff1ed6a8b46a21dc2948870d330e9aab65e2ea8382d7257e0b0ae1347e3f740b09f12f375f2e406207b679f68177434ecc8ee2a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2acc1987f7973a9902a71d382602a6c3bf313a787b9ba1bd372e48b9bd9f9dafe170b0ae6a97ac2c49c07ac5bbb217d85e0d97a2148676cf32a8b50217c85867297f31099a68c0fbe4d780e2802b87b4db65c187cd4ac7af87ae405820147508c7c0692a77e934508ca40b5dcff21daecd5f6a533366b6c5b1808a9c93d78d68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9349d5bd9e48e0d38673cf09b08a07958cf34b855c539a52eb75d5648fea907b43e7a285bbc04f5484c7672c5f841ac638a1eb685f89f8d03e7bff9808073f893545c44f2569998b8e02b3735c90c7c4f3f47e19990846fb264e16faf2aecade525112c66e19477026a8a17b79879e188c9e76cc20a333e45c89d79c04e10f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32623af3ffda38ce80d48a955d3ab75057ce9b836b6088693329d517272703f6d5989463b9291c1ffc29b5459b7e197079046e0da5fc632650d39826789f212846051ac64c6e6f7f0a02d7f714f4c61db1d06151ede8c1ba41b6c3b7b9402f79f73801a72e906cd879ebb457e9685b6166d2d696f721d286143f1129a31ce83e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha156e8990f3b85f1aab2d200d815395ed7afd13ee2f6f752a6261942a111218a1ba7e2fa42ca39e1d89e4a50889923e85bc2043b5da6d5792c8a884621601361d9f3413550f731a05b43c5d44b3a47f2b5f397080e0b1918d7ffec4d6e790c74763659cc4a0f403e891293b75643e964d5b9af4734b91a238ef3881664f1bb2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb204452d46db6013569f2b7aa44a05f610bb963ccb7a4f28ef89f69d1a64119bd46e1e4e4cf0ca7786c499f03ee62fd4a1dfa1cf2175c45d19d55763b675d7be041a495363ac7762581fba53f45183a83455078c6ad48f565a0a92f82db9c41ba70b4793f2ba4d25b67ff08041c05e6831c763812b1df44d5cccbfbaea75f64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0458eac91e979c8aaf094e4c51a3c40fc2a3ef190f5dc776e188a2bd5c3589d6d2c323ae1d0ff94ecab340ce674eb3cac3249978d7a010df4ef612e49a56dc3a0c189925b979d72b0e66ce3f913c1da893424a3d606d5434b09144c1b2b7950c81fb7c4dd49114819f4eca8f0130d77d9801a14e954b5e4bfa316a4571ebc09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bedc45f044b908599e1ef001ee112bcfc3e7e3c5af4c53e7769b520508c7d32564b0c481b978868bb57d162ac353512e5e62c86b1f136e3bc0b7a986c5c98fa872cf328130bd5810b86d886f14ca27142072cded175849fde9ee7970a6fefb0c26358d853de0b6c956813d53ef657ca3c0935c417ce48374e39b9a4668b88a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb77d5e7afc87950725b998cb83f5dfaca4607eded43e3c99371b50824ffa655c752b3dc9304c67459a30edd072713f3bf0f2a6769c0fcb81de01626a21c7d6a3c1ad7c0405f587c3dbbe3913bb1cbbfb335db010a48ee17277a56b52e6bb9b8af61dfd8708071c11e852f29e5bdc2e8c674936a4f20dc28d576d0fcbe7f9167;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb24a6a97b46c637cb3d4355d22d547b59bd353c7332cbe585a7e7703c5d71b6c6dd3095b564bc0c43054c4eb5e5c1d3d075a4f4775074ed7c44f06d0d4d6a837b186f3c459fd2ec52c1c45b6131d925b1cd511da97289a830630fec188066d30869106b31286ef40ca406096de78c3f885208c882b361f2de41fe5070938f0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54515e3b43b85c59dbae5077ce0358b66782af48d47c55923c0dd54d541b16962a490194cedf2728595646665514402f7ff88c2c4fb58507a15e8fadd5edf2eef5b663f23d5a40013ff0d8b4f3e9bf370a9bb08a4bd505cb9fc345874221b18527f4a4164e8eae4a59dad7961a5b108e65235f6748dd0119c36e4a55287d6410;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2f1def8997e806c133c553fdffe64376d8bf1edd95c74786358a1cdec96c13eaddfdbc727b254b8504b5bf0e5251d046578585d4b5f621f404bc03318f332344898768c121b7d8bfa02b4d4cceca5f50fe24573fdde153d2a3f9216633b4ba27e6a74c8955656588b6c36c2937401f4bec45858ff57bcb34449bbe287414ea2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h740f6f3304069933ae45b48eed2d7a55d55a6d61d4ab45b4a1b04689fc382826439fae65a19d0692c97b778d7b0c5a495e5f28c9a13a4c6c32f91e1a0d9410364e7c18a4933ff450935cb9c173e90d43fa608f3e25d22357b3afe334b44b28d9eb7dc23d7e85b9a053365702e8c2e89a9ca37e08d43f328d0d35a904ab09aec9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd75e1c9d8e50623e18a9615709f17a844abc4dda7f22182d350ee4761b4013994ed5c0d2832104b77e9afcc44e8dc91b34de102d4a01a4a5adc1d977e0d2e91aef76878278da0f87357a27b96e2918b5dbc7fe4215e5b0da109bea4dbcc8b5fb9b3b106b41cd23ac418f01b8e11df30da042af2d4d975bc287c49f67cb12ac3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae9cd36ed0404e5c5105ae1cb4f75eae4fac69b33d9873953fb62e0e2de07dbece8ef21b71968bfc28b8675bcc1f3879f765edbee526b49bcadb6e98255c113a36198516ad33fee7270aa7c44a81b15580df6ce3a71dab337436b7cdfffd3361946fad5e1637f3e6374243440cce03c61ff0953c1cb4d7c84d9754aa4ab0f17a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h756d8f2d44463155baeb01978108ffc3eed39c9667818445caee361d58a2b68d03c90d57d7f449e562a3a91640651f65c577c26d899eca13a8cb662ba48f2940fdeeb294b638384e7ea7d73a84caa1af47e9beb46e5a605c8b85d57ed8ecc76b06bc871eac25a88e8b91ef6d7f7fbfc6266ea5e030ecdb2879290e6a1545364b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb2fbae2c4f0b2f6891ee9496a5ef80042c13b646eb46abce379db0c196651363d63da7e8d57ba374902f408e47bc9c9de712446915d1f07cfdd7372fa48e578537cb2f618c00f48446910acf53241efde8b0accd7ae1cfbedff557e96ae4d2a3f67b619f589961c28c84c0856ae390e4439f4910c840df425b10e68a589695c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30774d58fc27824352dd12b9b80d396cda8dcc5243cd539c5d09c653b1500b705e44afb7e81cbb62c13ef665236af3d483dffc368a4e2c8ce26fa9dd3e57a1df7c5c9ecdaddbee06ac801b4050b695d04e1312ff18b5f6f81e963182d698bd8d4565a3fcaedf0b0f4b4b18cb14de9aefd0981a1d415227744186aa30f26b2210;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75eabf8ca077d1a28e79dbf40d9ea00c498ce410085714ed83ba5fc36b9a924b594922b53a4e34542f4cc4c03529dc458643a4f813bfefc3d8109bf7deea28ac8dc6f9717ca8577fab56d002bef8fb96af5b29738b41255d5846678f903787905e9352e649aaefa7b6e94f4ec3479488d0208e9e9fcbea2133a6c69009d3fa9d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha116a8eca80bdc4a6f2d081b5a18c70de73e37730fb2a73003a4f35f8d5ca88bab0bb1dc4ab4de0d7fe89cf0c072fef7a36cc21f6e06689c002f9ca1f5ccf0fb61ddcde7a8211a4a0e95671596f140b47e53163f5ea2708b6bb18e805d3cf12879c88192ea908e1730809e36abd3e349aaa26832d6d20661b1f6f43f8f84b40d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6272c4f85cca728b0ce160589a27eba5decb7525a3374246ab13f78ace4411e3f14c7872179054ef03ed5462ca4e0277b687c6a29e202bf3d827de4b93f72123ddfcd2dd3a0b9930414b5995b942ac364c7aa5190a0930e399b76af8a11308e09c05abc476ddadac32bd85a8300bb8571fe0faafed4fa28f639b8f4cf6131c45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd29a9ee49fd7eb5d7c94c9ecdd717f2975c98ea6bdb00152e0fd65fe3c1c8c1ca4a92b4c12891d7d7052b1f646feddba1019ed2545d69f6b0f935b085c249079669f154f2cda291224d908ab3b9a22a84389cc07225ea6740746d03245b5b03d4a40d34f5ea49f805f79a5869307fd46116baa0b4e502fdbd112956dac2860f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7263e9f7c122ae864c6193ddf8a82f7f3a8a9e563a2584479fb6242bc6a5b632b22d90d8f68f767f4d26f3c2819a99b2fc213df825c04b4c6e4c386dd023c9ee1bab800067829c96a6088b6d835fc950183da7ebb03e221f98f66008ef3e3a04fe28043347e00a00af0c30761024f6ed3978f94853fa3647f0d00d57d30b82b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd99b46130a7153a48019f22b2ddf875c08682d138bae9e8e226c7b370afe1e2a20dcd9f3033ccc7507e5f2f270192931beeb21f6941bccc5e6d4ccbe9331d1e3a0217c9879881df3e4becdb4e18714e1a6635b72a586ed3f3533953751d256ec8a51ab54674acb50cdfe1e72506c603c8e09928828186a809907a28bfd51b2e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5790967085cad3c26677fbdafdcdfe283273da6f091cb81a93fc1961a63143f1239778e5c9ea7893ea4a8d559009ea2c0eba059a50458ba014bad00bd850a5ac6aa6de25a7061d06d62ecb4cec973169fa4508ee8b154116f313ecec335c2f29429d64e60d465d87ac7579146c30ccc5cb7637417ccd142005cff65ad282b249;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ff4c06794325599dcd25e9c7b2181ce1e862e3dd71e38fbad7e902e1380b3f9bc8642bf957de530cea7c9e14ce1161cb6e9649ce30b9eeb37d4d25bcd38631b9b6c5f4907be7004784312d09a82a507fe8791daaaed136451f959aff1d89a4427a2baf0633de710bba0e1b0ef8d82286313be061be968680f29e52922ce9010;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89cd4d5efdff3446c1c484ae296ac5286a1da3fb9ce2c2a7f04c511a6ddcd9cb084f9778929e0af72276ebbe194d09562e153f5c8b85dec40f8e669361f3220e479397045675d875006d17e74daa37d47e4592663808696e2d1adcb32ca2b29e5eee7c7a5502dcaa51fbb38fea19169ed2e23a7db2d842fc19f8c51f94b9360d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d3f94c52193d3bb943046b7dd976ce4cc9c08d28fba1fca22294d5e05d41350fdcd87a45f7022a5ff9b501a77f48efa0fc151fd502c88708baaf626c82a61eee8da786e45b4f2dc0174bd314c9ac3add4f2b9fe8923443d2ce361f8c2fbad854a1c12953e8b3c5f9fd3611e26ad2dbace64ea13d56e3b1812dec231cde8e94a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc400551919f2ae449df5cd7eba8245a446b4c2a478d51f54d25acae3b6bdd5296ef32f724a7ee0dfdf269f03d3f1efcece736e8130c4a7cc09b68b986f200950e0a240a79ee7b856ca260392114b42916699691b2bda1de04bc25bfca719a7ef2f47dc3313a411ca71f42dec39832acd5d6d27d7d086ca8e17d03e24e30a166d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e15bc62666a80c5b4a35fa26c0fb35afe3a453c2b1f817745b3cc6428065a692a2698d5ec33ede0c1d4ed9417321e6cd8124e8562c63940e34a1097a716bad4ec9b29c6c49b36ad14c82356531916c0de9fa523eea67c29aad0dfa6817d021c686bd7600c54d3b3e9412617d48c140359f15614f189d9738064c8d4ff72f028;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde8ac34f6f7030c7b192af291778058bab8118b4f11c6d43c97e7c05e4465b3eab63ba57bbd8070a7f98f541681ed60f3e781b2e0b56537cc6f4f692fb49584eb29dec8810e35cba6fdfb3b29711ac33ca7cc30a2ab5b596edcae0e6f23bb39224ef3f082c837faa77d6e2a1dadc225c9bf5d1205ec3fe6703f55a1dfd8472d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c4e193d0f2fc0923350a72c5a8ef5a67709a1cd0426143dd19fcc053299d191b84d221f6c1c4d8387ca23d07ed6abf316e6ccd5556f41da7e52f85890c050ac9eeaa07e6d49cbee633d5e4ffdccca9b651b33226a05c4f230efb3f22b93a5176be02c33954c6c1fc91c797580c1f553f1c2710029018b08ae0f4d3f3b2ee8e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5944fda0b3fb5cea52e970fa6bf0d4eabc62499b57ace04401339d9ad30188453c7f1d36fc06a9828ae8e5bd3094b13708b6252af8db7a861d1f8603ada15666bad165257e3592df7336b028fba63b081befef1c1c230d386b28c7888d6047c15328e65331f4a62bd82fb49b5614986399f90e8b134aedb54aed475e2744c27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a3923d3a9315700a72befe41bbba48e1aea4cedd4d507eacaa60bd9bd5a47564e5f7568be23321700ad33d4e1cb7b4a0466e42015e1924175abb58281df4cf698824bd85c545b36d0b328bc36348bd664570a70643a09a6aa694856684078ed2d088b4c2cfc1e44784f01a65fd5a0a3b7b311cf931c39c5a01c054f70b9b810;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa028fb3307ad4b030ef4c99192e5f3d6f52be3677d2c0413a60cae96d8ce43484a5218720597d5726f7edbf3b756f5cdca80e5a82a5df7c17bfb4259d70cc3109eae5904e3941870e0a412f8103374dc464e254a8f703ac3440ad249b1fe919b4d47dd00dcbe60bb6611dfafb0d8742fa2483f1ffca7936d5e79778554fdf8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5bd342a00c6c716adee2e1563905c2bb19692b45fcc59005c470d8d7736f4a416762b295ad4112d739023b724b5684efd8457aa07d727b14d7f610dbf7602be0534302509b0b7d51cd23e068a6977432c3bbec295987a51f53fef6f894e653c9740759aec133ac4ec75439122aa77d422479a8fde05dc4a45d494b1ff2256ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2be2f1032a23c469e81853450e3f17d909dcfe3e472f25431fc10bdeaa9f93bd59a9a25150c3605dd49c8a9ba51fe62459134ac4215e7a29fe07ed3301560404c184e0586cf57d194b16532451d8079a1f8084331f9496e9eef0a66aaec6bc3f842dcf4d80939f3cf3cb7786c8f95c01aa1fc05f9aa88200630d420bf84bdf03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2bf653d57d8427ce59fa7fcd5e4ce1fa33efb839b40242a056e357e1241d47bb3a2a488d342f41bd6918718866189214c576afecd9a13d2ea1181edae8e6fe80d8c704c2829dd6f5f2515aabb928419d8f07c248f16947bb268460037f602a01fdfa835b2182781412ec031552a96af7d2721d1def6cc8dd4b8ac172a270220;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1718f78ebf80b56c506681269bfefbfddcfe7c1069d0e08ccad527e9cc71836c19d623a451cd0fb7a1f0f4f46ff80a65af2824da68cc1e7b236b57ce282baffd09c6a6795b0199141ee2831b58d8419d6e0c9a6853957eec6e70d7d18826cde41bfc303bb7205fd8f844dc149898370238117a492b577e237d521fa4529882f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab5d709e137eb434d47c4ae7aff087323137ea6916205219cb27002c5414061aa2cd8ce076bd0d2986e23fc306b493e6d278ede8b0fce73fc3160d95dc043e8d0e5c12e9c2d1630e85ca6e5fa0ab0c70a3a22a92804ac7470067f2ae0ca546d7bd905fb79779aa33f360f6b2c7a424fcbcf029196e64540cbe4581951145d6e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fb3d9c2a96c380cb720c528628ef5e9e9fc734567ebc318145be54a16fe6a43bf7af185e12a913b0762266ec016ec46efa5a5276bbafcb6c6b7a71d4906aa62ec815081963def94d35415c773a9c0c9953486979f618ee923d52135069746cef23c4cb8d0ea1ac85f9d0b4ddbd53647b6b6344f02d97d91d8be8f32f7ff34e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h938935610c0cf10df6ef5c8012b31705d5cf7eb695f01dd683731411307df5e13d497421c64693b07ee8609a958881cffdb79e4ba4bc18cb19eb6a7a085e58ca65aa62cd851a107434da9a84dde7882f409dd0aa68b908da5563b41bae529408537e2943c1343990f9e7db9ac76eb5db9f954d9635aa78157b0d8e849131886b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc43f669d58dc27ba8fab472a5bd9fa0f353d83650e11d7610dddbc1ae3aa6dca3ebaa01478f72f2c99d1ce13db603e06003e937e294459edc085ab491779631cb8012b383ac464c9e6ea4a4940a7309948fb19c9f75bff056ea0b1e23c740b295ded22f205b5e629a7443f08da56fb4512b716e5d727197756d02941549dab1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb205f3f0d0e5c07667d3b06ecc00e3dd218b62328eaf32547f5cffb1e162905c77f17779607143e168a03ba9bc8f6a9a0a21be76cfe4a0b90b46602186f253ed88ea81d49b857c4cd4a475bb5e69556838df5f5131776b8f3eeaa7f4141efa8bbf666525cf4960f3c2da81559b7176c069fae1679737dec0de00458f8ae4561;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b3a453d2ab0431820fe70ead87972d8ec378a54e31718b05de3e051652f11f7e44ef5461e56739e9e3b4b1310bd1d5bc879ead38291fac2a2f6110e58a9a1a823bd4468eb2e8e28428e50dfce08e3b13b6914d18e522c23037667e6f924259c6bb100703e9f387a7cf565d968edcdaa8054b4bdf2383d9f8687be33bcbf73f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a6f06ebc572192d19f8b983cdb48688655dc6b45aa7a033ca54ffd1da44a050ee746f37196c048b9a95ff7ba344ed7c93cbb25c8a89c7a3d13955eaf90712298acece5e8d36edcaff0390ebb4016b62727fa5d3fc043d4f56b011dbc618ee705dede0a21cf801d7781376465759c4f0c68c2c24f79d4320bd83242c1c2ce3b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h933eb0449b80623a67fd9211141063f6bd3ba55853965bcca10365cf81c355e44d3f654821028b45f66423ec1b00065e73bb735f06016b893095c3e30308dca1b8efae42a2e9e450c97f2c3d183834a89d6a65399b7735845cd15ca4ab3e521cf2d80624fe00f08906168b1faad632ca2d60be9d645e912b2b7f196c82a05ab3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h510153247a32a33a23d188902eab2e880ebb0c4c0883d9f7272a0f94ce8c15c9483a4b5a6ce81f97bbce7884198f0c61d3243e15e892b1918b62578f0e984084327016de7c9120e31ff400330545fdfb3f1cee8ec07f9256a65479b938b747c8d184fc259f6d901da21089be538e1da43a295091b0dbba083c3bd6d201cc3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4db400b1061b354478b438b5ad0bd3c5e7f06b790eb11bb49e7357e04c918b7417328498f4e2a9a8dda9d7b1fa45542d66f43a225d39f3d4895005eab7fa40b23bbdf659615520766ee97b0c88107fda3a4f0581243eae3090a42f5ae3ac43e7628e9a3b329f6c14285fa637c5e0c086f87d9d55a32d9d9ee2d9ee94683453f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb3aeae79db23e3a02e32f046ba00345e8157ccb4ea4706467b8255ad4a3ee45d7641fada6af66d3c44049aee1117dbcbf79c01fb3bedb92c96a6c193ed089b1a35a7e5b6874318d24a6200a4396910fafc4f66368d2c18c0cbd3be34dddb3b28eed2c99a3b92edf63ce91eacc9602b7c54b1824a8ef5323aa87a8fffc49a715;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22a4a88c9ce626664386f24211ce5af3098affcd96530d08bd3383fdbd1567b64810010ccbefe9e786f366d40f4067359cefc2dd1f40ad7ece01b6f8310f9599bfb6d69d12f8a9da02b725e1e5d86a2e5a3311b83076721dfe59be2c79bb9a9452244edf2bb78cf01955cfeab229afa63e1f1f773d8cfd62b715f71d009b59cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h609a1dd4b26fa54b8b836c9fa7a57a3f6f8f4012f7fb9cc05d3ba763843f6b2660d2b0a3219d7ff76e49ebdc38592f40572872772452e10efe9939c989f0e46c62bf0a0b237dc9c5f2ca84ed6cc313babe415750f759c0a87618e6afdd81ec13265a1f3984b680f831dd26d6770c6cf93832a03d9520db4ddf9de672f9b07511;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc090d4cee96ed03bbf2858233fd15474c133acf9d9c33954fdeb1ce001404aa8baeba16f92ff99b69ad2b1589b19dad364275936912b692e6d8c56d6f09110fbf4b0ad619e2244c099e9837ec967b07b880016b75d20f5074249725cf0434125c4a5a0b477ec9c0d45417e47258fe25b12ed304332d264256d75e4ace326daca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe04b265b52cf369d6579e3a0d78248e34ca92c1e3fbd699864718ccfc49644cfd8d2cd6edc6d30f8ef0a952842a008f534bdfa9bb29c4ab0b52af11b448b70bd90a1fd1a385693a1533bf2e06b53d2b746cb469cd17a4d47ab9b1b6f86930dae0a21d74eddc72584e1cf28a3ff12adb7dcaa04b5a50c5cb67d378a24b1d8e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he86fc87c64a4d3823fba7741dfcdfd7b87f34b378618e18ccd4b540791f8e44b07bf23bbf972e7511e622461a517ca3264c53785a0764548d77ca3d6669f3c02af0fb15886fee85fc10c6635e76391c00f85638f852aa2e1091087256134815789382202919f9302df6793ada7a37f7843b5ae0cad5c442c211373de0af10947;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12b5935abeb580985b3125bd894f35d4fefa7375117b1730f477594ddc755f6dea77239e79cb2fbbd5fc42a227645fd771acf585b8c908ba81d7aabf6bc22fd18bddc1969703e89c14b48dd5c35524a706799cebc6b31b5d63aa68840ea715eb3265ff0d95b924be36c5a6029048ade43debe39959e0bda35e977acc7df5e509;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a76644606f0e6aed13af45c3008c8c89acd4bc9bd2d6982ace37c0020a9527d050f2c26817380f027a05de7c30264033802246eeb24cd3118b2e1438224c84b4c6b9a0e779ba304049c5d86adce6c94118461b5266d64fa798d344406ef449fd6b68ac3f952696a9a7d0e983a4483e0fe04f0dc38c0c34421a15999828bdf32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67d94ec31b21cf88eede955cd0f0a9197a91c4520e2fc942a12ea3ecdf1723bb1c37bf6b60b4b8f89e1d7c63cc1f9ae070702ffcc0e58d8109a9e68ff6b6403fff3ee8b708a0b194a227559cb6467d88a93b1b55b73a5d48b3c6e29a602a5529c97dec37260c8c3625cf306d1eed71d793a4c28549608f927f8d0e282d1ffdd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b379d1e9a3be85fab19543ac15a584a5021735f5391ae5e342234e3f57edc4134a0b0dafeef0c143fd717a55787326b3d3819abde82edf4829dd9b4a93383f34d749f1abf78eab5557b4143dc91e211166ad9925c1a42128f3fbee4a772bfb5ecdfb692f47b11c9d5c178fa111ad46b8500007bfd2f55afcf61428d9328c351;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4038a557c8335ec42bd1b0ce4805918a63e3c858e520a88fc2cc45dbb11eab4fe696f0f608bffa2c1a6372daf895697cf778e2467b3a32aa1f3bb1a6e243b2a486e4b86b78d06105c5900d1587a729e522b4885dc3b049670dbb6745ab4b32b467f014929ce67270cda350bc024e5d7a73e8bc1ab75080b1fd7547d056d4f16e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdab48b85b0efed871c55f3253ae6c06da6d9faa5f5dd350f8d95db1a2bb3aafe9ded3dfb93e30ac222be38cbaf67f57494b78116303443126c93f3170698f94d9faf599054efdc50f159bb949d165447cd677264ec2650b2d67fa8d9ce46732553da862fa9c35d43750adf58cc72034913e7eafb12264ff5ac81e1361ddcf8b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d8a056bb307cd56b87105f9d263e68152e3f57d782178846a7cf57fafe21a7873823abecefde3e8f98b7dadb27498c1c452a26ab2337f200f73e095c828ecd834c159d051ec855bcad14c23385dd1eb29c692ee23f8946beb610535ab236442fa5bd089613462a9f387c9fa93b6a06a87cd2a47bb41c4489b05b895c6256280;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb650d9443706a5d97a36202bfc6d743bf56047a123896240c9397dafffeac87954abd1c61dd36a0a59fcbb2c44fb12a443dadd8bad2a90fc8c5025af01af4f64eb0fdb98bb6dc7df686f756b8ca479f0456a08b7ce17d7e949f8bdd4a0a2c8155fc272c0413c3b42756c09ff4413746bfffa6a2f39cec5aa9c7933f3664ce896;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bfbed7c6dcfaf289d63824741d51aa928e9511a11ac7266c0a0ae0a872159d94322d23ac7e5ebc6b602d2813ba7a2adf2fa05661e62ecb8ebddba528a7e5c27fdf2468ad2a1785ff913ac13a7d55bd8f3aaac697e12135668a8788cf186395843f96541af4777d09b1054560819492b674a8551a1927308114853ab7cf89512;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc772db07ea47d4ee22424c6191cbab18b94f6ff6272465bc134b944ac4455ce0e0990689290a33bf752fd8018815fdb127c9b6ebde682a4727c765703e112f4be0e86b8fb9b9bcc5c8d00fe794f5bd6ce4ae697b8a0ff77b62077860e4e64fe06526499ba155e47a8c5eed533b5b01f49dd48b48d508ccbaa9ab1a9841813799;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74a845983fa6f672b1b7dff55df52f4f31078628265d4db9ccd76aadee3433d91d58e5cbdfbcd8a2f57b0060e506ecd0060efb17a8f22aa180df37343966df4bd96c93be5fb09c0fda7cc18543f1c023476438f429908a488f88c96f1e5f966b83d88fd240aa49b39bd5387bc7cdf9bd47b4831893c0fd3aad9735a46c0da750;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h544bb818f6b13a7eaa0b96a0ec651268a341b6b8719b8414071abdebfa21f42103085a50d44f515056149547cf7aac35e93fc82878e3b45f9456ccd90d5d8ebc1e069ce5dd015048c41acd37aad3a1ef5a4784c81a6a6ceeb3e000285856ca8646b2118544735dbaa31648f41f80d84d2c5c5307e0a16e2bb6f5ea3cf43d823e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf912517495aa8848872a1f1dbd4e21f09000aaf5094a12008073255940e6c333a71e34b83ed4f9cdfda484e7592250d8de02389c7ef052171e03470a1a9a3fc635bd1c995b7edb54f36b405ef40319805dc6f69748edb08d3af7781d4fbd58c11e5a64dc9a7607a7b01dce7497d81b873ce2f25f7d649dab23f8c4db3f5673;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5fa54fa9ddf51e87326f74522a29c763cbaa36fb2992d8333e54014c91e9d369004c4e0f8d842a53d2a3c15461d23cc16b2003436decf9a90f3b0d3fc9332b8f0a86fba64d306bcdfdbad78fc34806000a91fdc21fd7c55ba95bf8b905a6f40b904921729bf939e929b3d6f9eb8b86b0a32f816c79dc2587048291405677a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd67898c66dd5538d2c768bde797c4c7a99d54ee47977cac05baded5753614738029a792d2e5600e32e6037e6b19f0ee2e6126ea5e1ec6b139d529da85b4a84f52deb061bc97c4f723cb4be96af733f8fff656755b79ccecf73a5073376d18b0e355682da64796e4389cfec8697e94a245c234a4a20b42039294e07932ad8ba39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h224c7fd4d011e96bf0b2401df9306b39aea4457edc4bbd1ed58aaa115506bb13124917b3107b045092b7597fa11c3667f7531f4f0578fe80c0c2b1c0c9524ba95507ccb253befcc77ff12ee932d430a2c017289ce403173416e64ae95b88e4b85871499b7b18d8e6a4349afeaad0fb7dda4cbedf7e5e8468486717a52d2cf98c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9344dddd20dfaafb491444c259334d9c923bca2c82c32216b394d8693120884a97ef6d9e3ea73ff6bf238674600190534da3071ad02d13169ac9416e90d9a5d77f8dea9a9a59e444710f9b27e140fb0040750efc7c129250ececffcc814a734191718b3241bb93061ca115a8883c1fc10a4b6f376c235e5b9808592428858c9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72d80fee5d30ecf5988f54b7ac772a9700342d9e371420afa3293969a33fc4d7857bf59f1835ce9360f30c58bd3d2581d1fd7ce56df7091c374b603e2daf188e79661dd7593141439ebaddaff41369e346f0efc1be968e5ede3ca039df1c034d8436e0bfc65f018c4454c02c76d9699fdc7afb79fb1dd0b414dd08abb0bfc39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62f3df7bfdb2ed8c91b28c64158db2f7e0866a10c61c5d868813d30e852f8aca8bd441f1d0ec074c108705b8912180d9d66667f1c52abfdbb50d9c90ea4d63b93e7b888f21ad37951e979698f0928d529b24fca0d2d90f130b619a0b63b7f91fc57c706ffe8d32a9c57f45d3c679bdb9b5af8590c676c75fc57b709adce6a89c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2989eb5adbb07145daa86ccc7a2a60577830d9b96786d93eb43088c5662dbbf3f042b20f38bca9477d07abc39a8d36ecbdb83abe9130377217bd00ff72645967522e6a5782768711665ebed935a0b016f1d4289fa9d9f21b4cf3d0bd23184e11edc196a7d10390b7691aff6461556a854e7091f9dbc5c9f065b5e6d3558c6f8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24be6d01ec5e40f8c809c2ba1d45919ae94a97d3e1479ded26bec1e909c8c0ce4ee4865c1497af6676fffb86d4e3a2bb6fb4c321f6ab303aa812c565e28834af2f9a048d0caf8004eced6a865c927c43decbe428a7719c8981697ba52d4137e51d5bf7452475a323c4e58bac9163071ccd99a27b580ddc9bbdc99a09bb74b4a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86b9eeb4525f1ac70583ef8146ce76724ec8f7f3564e5b02b1f69317d0e955ee8674e856922ea19bf28efb7242d5cf8a36b50d0cdf0fb64d4e4059e144ea7b54d8507dd38bff58a8c8c9b2435d2863637b565c1f1f723b906e8b385a09d43a871c3d294d47bcb03dfd4c650a1d2158cd0b227fe46213ec9d03efb68e8c358fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98187f7f57d2ed35d9b6bcd3c5ed80289c0c7bda995fb23d31e89db36beb03ad9e6be335bd7e4c9304c02038451575359789fb28795ef2bd52a55e8b8c671e3c70e0cd99b35c4bb20962e28cf538e31f8ad15c3693b7c299db1cccf7d097ac3fcc27885edbfecc10fb5f024a0c692cca1e069ae854923e12b7468b27e8eb8625;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72580fbf521633e4b5660783f34009403079fe3513e55d36e879c97ea1fe8305e0c04285aafb8af26b88a5f20855f8f4880ebe2f797036fe3a324d1d5d9c97d1f255f1e327be3dc5692d25854d6c816376a5d339db374666d34e373689922d27eb5c142129d3971b2138a49051bc425387052ccf6f38eb6a76756e19c02fe090;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1096f768caaf92cc58736295f49ebfda1cce2d0f690dcf765f0e507c8960432cb6269b144834f18f3190e90bf0958f23ef874e8ac2d9831673cc328090a0566f0cf8a7e3039817601f8439c386ff9992b9410b11fcb26c4187349ddf106bbb1e5d6cd26b74609a391a60156b3c93e8f52086ccd1bd1c87a550d8e245e25aee3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2446ecddc814c27f6fa52a2a3290a6f987027a1586819454f8da31603e52be95ced0df658be68cd435390c59fe7bf739094b6fb156922e5381b702da427be4ecae9763f6d92f7e5ca00cd716733b4138a510d35c4276f5672974fe943a556e2d5cdf31ba7441c2f01fb004b1acab54ed3347b1818ec717b06527dfee0d6d3bad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habcdd58797209fca0a7c4e4882cd45ff1222e8f8c829cd76426333c4727b328a74be0ad1c4f6eb9d8817ca32c38eb0707f3cee779ce558de88c77592cc13e03041046e4acf6ea0f633444836529e35a7e2a028d0ba0e2994676a45c61f51d0c66a1e8e4a0b9092a4f3d68c3e39f0eb2562c7c0d3ba5cd4563677a430f83a126a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8cab48e11a54d81cb65348aa879cfe1534b4127f4f1a9a38869513356ca36d9c257fcc6bc3221a0f9ab89ef1336ccd5f51a07b71265292cb6a069073f0c3313d92c8f411844df4d68567aad07e4976ee0a23c5cf347c58d20b0b06769ef3d80df29cbfbfa758c199f377be6244e22c4f3e6e872c15664f7dcc9336860cab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7cfdcbecebf5375757e819cfe26d1341ba855037924708282c1f19ba15e09268bd6fa83cf509d471802325a7bca85dd791b457cbdb1e00a3f0bfa3f82d1976e43e9b3f9fda72be5627de71c807ce8cf682abe6a0aec31c2cf2abe854f2cdc20235d5385a374d4f8470b695b8e51ff503ab1f54cf07ab44493a5bcd34959c10c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51b7d04d91649fc05f7ecf5dc3931588f466f620f91212ceebb3c33a6ac378b0e0f9cc78588ce39bf6828f46ba43e63f154547fa2768bb4c85d35fe81b4df74a8d7b797356ea6b63c82b58bb6cc100cf068b51f0b34066c109c34c290eae0bf9d95952f29f76bf3e79b207d49188301a3e07881ff189a6f5c9709544418fd0e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68709ddc43953810c7e865081be6b372340cd157349a696aa110c0cf59202f9781bac43afaaf72d2515379a223804cac8de723bfe47589c3dff02e0a6967a0b18ed99ea4ac838812935c12bb944cd357c3ca5bac0cbef094a2ead5824b6a1d4fd273698cdda1dc5d57f5ac93514c96f9dee15b4c459bfd66b39174fbe3f76526;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98b2996dc54a43616baa0c3c1043812924c50787786d3f9ee3e92cb6e2bbaf1ab99c21e9fb4157ba14a94105abfc8773737a619166f407f82b946b98f98b260dc70789b4c80a9056fb4f85104b593caba0cfa38d4166dbf3e3f1fbdc79215d2968d4ee5b247d8c83a2416aa943aa760eb4f7a5daf37614f3d17c53461b19d37a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2b5bdb4498d010871688da5d87e63333d4a5e4cfff7a2bb4d0f2e2ad1f1f579f2af1696710f6cd20f17f95fe5411a7a2a3d850f84b434aa1142f2b43da96558140ec277accb5f5dfafdf56d4ad811ac08087dbc6593dc50a3b950dd5434685d71ddd9fc1c1c494c388ca1ca5db49b508f68ae3df5cfcda86c4110dead8f3b56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafc944a94dd6db0be45d1ffbdc76ac04febbcc5d3c5d0d44553d1e699ccb00c0b0d28a9ccea1ce02a5ba470c39c287f25355602e92cca75e894b1c1fd9db09416d6e31db1d1220cf4281cfc6ff4184db25a5b9225a4f27bfb0bf1fef493e92f1e1d9a547f8f77c7e7840a7e9b126ceaaaa5e00daeb8679f26723aa6695798558;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd960601806d3b338dba11f81eeeb4373fda95926b0b0eaf45f08612f883ac65b0f0b77197e7495b52824bed5f46893e243f15bea613e33fd68a986cc0e9ffeb4156f351e77ae81c8634a0c0076acbdb17a53036d039b449bd211cca27923f4388dbc55fe8dee6181acdd7eb1c70508aa43b034ab0f223a91c39701778d573b19;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61bb1d3f74effda299c03d219ca991918ed2a79275eb513203529c074499c4c320ad799c3b58182960b2a28c3cb10e33f5ccbb0f5e70f0fa510549b58d668a86bcb8c1d9824c053f82c6a5dc3639849683540d2e90d306cdbd7d03f9843e043077ebdae1d949cb949adf64e28e64b050c8222857a01c818bcdaf2ba21875bfdd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab58286ce7b16c07ecfb6ba15fa5469eea2ee72d9bffc5d7e9dc4dbf22f0df225f4d002bf3cf08c7ff00c9782b01826dc01f35671292dd0521e1b20981e97f9c3135730ffa0a7e4a56b92ef62eab59d48ee3a2bc6153fa786e26b05ad003113b0aee5572b6f90c3fdf77f89cc978325236448229aee8eb5b7b71261fe1b10b2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heea77e456babeeccb52c2d747bdf359aa9c41e0eb1fda0f933effdb3c4048804823085c623ca66c5d0e644fc1ca9db2224c5534977cbba54e3af0b4f436684b04b9927774b3ca3ac07a7727b69858ea47c22cb6eb1af1cd99e716efed2f8c653d50532b41f7e472a9c2902330ebf1b53a9371c1a3ed5d0b5d50f60f46272b948;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e0d454e620c3a929a96c6e1b6ac4ecf37d957e23cce770643887633bca401823276451437c20c72ecda10b245b9824e56bd0a010670eac0678bf9acee8fe2516f50f1be75849086c8e469b0c52d6656243abfc4d51699547bd21e99aae3129a5f3b0e632f793b2fde754c3b8553d3ca11a03c395bea131b3b4949093951659e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d7e9f25b9e33e82e9c0e663d0f1af19ee9d7a99a9eddc6961e104e1b65f614ffd13aab66d747d91b0ac6428154dbc8c42fe7c7ad5c8ee6956ab2f45130238fbd7550da6baa88ba28e966e25cc990ca11c37a8d7f94f9cb09e647de010b2d53a15fb8f9ddd629efe5ec489662391a9df6959d3407274362706e862685ea4242f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ac5e398d2834709c8bda42cfbd6890227a052862108f0adcb34a96052f6f3ba60715a54cff9dd12c84f35b4447063fd59b7c84b3145de9c1c47d1c6478440dbe4b61eddd791287ee5e67b4195ec201d1c329eb9899aeb434eca92c31f6d8e5996c33148a18a0485322ac9e64c3c355bf919524b26e8c70c147ad0f95ea122f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3151f9ed8b76892e5b831bc09c49e656d9c50f8b1b589cf02013ea439f872726849e5dbf17acfe75619f3ad30468f98af730f62922b5b374fb384c71b7fc4d534e338f2c0ec0bc1cde46e075dbb268db46bf50535ff2b21b97d6926e1313d4b99ce01ddd95b262a92dedc4e4eb5c9f67d8e95e9858110f7000d53a17750919ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0ff0c187ea3111ee9e6281a974e41b5f3f93c1dc732b5f2b9487996229a8785bf55025c98de7ff6764ecb7c000e68c2b9e85c2b1c6aab9daad1f917a3be94d78663eab35e274b0ecdade6bea0d92181c2d4a29f157d63649e4cf6ccce04193efdd01dabaf0d0b9b92e0daee85548b72b7805549b994b9bc18b44e5b26e6e79d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h174af8917c6827f6a09b4c5350b37de2a9c90035b6203717ddeb4a874be223efae4d882d6fb9fc775c1c7b8ffbf1d8e7273bae1824718ab397ccb8f6b1a00bccd01eb17ad032e5704032c75b889825bd235a43df774ff03c172d146636a394126bcbf88c20221c8d3904084ecb93258712a696f028c2d15ac58ef90809837c61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc86f08bbe666fd4e74363a89567f58b5cb19dbcc17edadab3e9f32932e98e3d148e120b721757f609461c7323124daad25403dc31de80c74870d61497d5372e775abbb0bf243e204d91477e76c2d80374bda5dbe749d7a0fad5006f02fb7e63e82d1bd09f0bee23e6f48111d5105cc7f5efbd07712c6e129c204a76879c1ca46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7fb48c2a1cfca0cc14eeb6cfafc77d2222715732403f58336f16719794e7a07a02d2fbb18e2eedb39861241c6afb0c7bcc7f54442230b1af8556aeffd1a4fd8b46785f88e267ed75388f37062bea7ad963cd4cc9615bc2ffa68f7aa6a59a79e8f9be50790f26f58210e0d7c71461dfabe80a392e4c61ca0eb6e86248c7e5d77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h290c60221843b39dab94eeffc15c8e65eef5432da146521dea28ea30decb2a907057d440ba9b193075dbd3cc260713152ef29f1cce1be2a99d4f44dbfb84efc91bfe3004d52aa6488d30d8ccc4f84d6145f44f6e80449df05c982d13ee228737ccf0e6b1ec3930ed554ada65725078303e102c9bd6a71a4bb3c3254c021f120c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h721b9fcc2826a619cf32f7ecf4b7549d5a5237442ff06b9f7a040c7980d01b8819d4168b9b9e6539c1dfcc313fc8781ebb1b00d4d97887b66077fded9891b923cb1cc4761b4c44923454b1d89af091764a4cc926bf45189a35afa6c15fe511cfe36af313e9f28432b897ee0877f317c94e819efb9f9697dc103cab0a921c6018;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32693cd49d59c2185fd77b6c88c8afcab824e26871daf007d4574a8330533faa0c0c1afa32b12ab558da9f7453855e6a973a3067fb3084bcb20de3759f46a2167418f0a705cc6ffaeebdacdcd6e391855c47998b3e1a41be87f526f4d809fc0b3489217eff2f1600ea32cfffce3a17f93b9a5cdda281679bdd876639be206e1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8c2bcb364cca0ca8997a79b5cf9a3b53e03731bf6ca0c3cd1924d18d7329695483ba4773b45abe43a84f735b8ee4d9f034812350ce4ac32ed1aa36665ea445497035c4bad9340225883cfebf820f16f8a8afb03a5f1014fb4882d9cbfb02b0874339814a6273f76fb9dca7703c6606f66208bd75c24b412bf04c6e158fe2b67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1548af582b0e9c650af9c073c9c853403282554b0d47a0005648842771829126f2e8aaf625472a40792e0a954d7391e94d3d9cf9e6866525724580bb4c5dfa1570f8e44f6996649c21dbfd558d21aff516aa3e7d80aab97fdf0edbe645ce2d5569bed02fb7688e8d08c12217a8033cab9360cc6f8f975ac90c9a124297bc3f61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15665cae848d63cf3e2a7ccd8433a6576f4cb52da3baa87e08a37e1af738648ac91ea7248526c236f2fa74820afd314c19317a3b716f2116714db4955951fb4b96af290c6657978111a1e1b8a38deb51ea86b5aed2bb7f9e3d0c3e49cab12d8d512ca0d909ac33dcce44c63b5725c3475e32289f3612d66fbbf05008b188d7ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ceb2b34ad3dcd6c51b3fe6649491e0e627b48c90b28456626eac2a8022d63669d4d8a7eee0a17db19007f0570706659198a5255080ef2c4a3058d5ff881f390b361f2b10787ff96cd7ca925d81949d8b0eaffa297f554775fc81d99bb45df3bd730ccf2bc449abd00f1adae939b998f93e68b3b95d647f697f5c4298f583377;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f810e19abb3af7d06f694a3983e8b8038c53a05adc17e0b0f35d632d92c3b4023281e55f2f818e1da75e4795db7bc6696370e19bcb50d9a00ecdd9ba5032ffa392807809939a174e679c4be18c73e43ce1bdb0b6f38e86f4728c91866b90fafd1a16c4a5c8c35c01c11e26a9e0c6a31570a5030a175010444ea9017279dab26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8bf0255b48a491558df4de7eefb65b151e240ff99ba2a4d7d9c0aad3cfbdbfc3a87ed5ef08290960664ec3f6f9f84b2050590011809ce7f60464eb98d41b8e98ed03d931b1c6f94814a595094abe8a1e523e71ba82aad1f383bf61e7d29025ef2a56d26729b5126da5737c519f09f8bfeda75ebb84d17dcf99914def42cf0d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54aff35997e2a1b423d34ca9d33d16d5f85d9b0f21136ed9d859c80265c2edada03695b62bf443c0af25ecabf751d28266d805868a1c973fa6e08fe29eddd7ea969f6c9e133d7d596dcccc8a8eb1262ac0165cffdc0f841c11ddb4e8bbf226e2b98a5b00a64cea3cdaf25e39ba60e97fcb74b4b65a1f15bdae8c5b0e6a044c52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb429fc3a4b135c75efbb0fb31c46b81f79a337bf7617d9ff574c94c7cb8b8d36629c532397732eb03f1f724ee5e4ed72fe616b4cfc3ef9a1ef96977f4180718e3b2dc6b80b3794ca7ec0d043a103b9c0820d97119fcf1400db1492d746843aa46746b0b893ee1e641a1f6f879b4424987b72dba26e7825ebaf43b0c0fd742eb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c87b53bd22b23ef34f0f59aea5915419596e222f7b3fd3503ad42b8f52ae4a8b442c39eda7db99474d5aa154de3f13f315b79a4e2cb29f9ffd50a76a786d0ab92d318adef0a56c91c8955b3d151060dc3401235f70809f57537601cf60006a2773c51406c526ab823ff570b0f106b0b675de491da31a28bd863866bc1134d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50798df781793b963b91190855cb2e84461a2ef2f2b381c872140fa631a938c377109b89004e77469ef34bc4a77242afafc0c6b86c39d45b7d000306ff2edf97219aaedfbfc84058aa04267d68171fc1152d85c9edfa85417c1405866b9027fc63bc016f3e5b60c66f9f67347de0e7aed78ee558d85c4a500cbd164bf896b90;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd30d0aaa4a79511a74ba9dbde402cee49f4e97c3e230a891359aafb5cd0217dfec6c94b52da2d1f108af4483a64995e2082381039b31023b3ba272851d04fc1adcbfc5288a7b0af70b68daef49e1a448fa5c363525b8ce36abf15ee97ab7540690f050aaa681eb3e41af66be8ac26d9418b22872b3d4489e966b941d9a8baec0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661b9396665ec04c70b99e777590ecd1db7ecbf98843b1feb9f33d3a92060d52a2a1dd377551b6c626b1e880ee755eb5064e65e45a3cd413f8c638a15572e653918a7daf4bf2da4b8ab537f3b33ed18356200874cbdc62dcae18cb12377ed89537c53613aaea65bc5e7a9cf7668aaa65c80b1a9c70f608f19386961e5f869b99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbea778a2dcff618834c53a25c9a4f9ce63bdc8187a7dea54d23c3aefbfdc1c705b278f40bc3c831ba520f065b41014064b589d4f3bd8061625bd7d554d2d54eb4ec82858872e1fb19a3f6227428764dc2f04fa52f439200e77bec01a2e2a38bed251a3facda8cd6ad75b35f211b65a0276d711c273fe9b00f84cbbde9394918;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2aef5b75c5a7a9381a4d4fd13548c24d0c0a789abaaffbc83a89e06cde852e0cc4d5f693fc58abdd5daf9449e192206937f86bb940951044ee0e2f92bea36d18b64b8594c4a4849bc5d569f78de577a41fb1cd8cc2389793e84d8a0a0ea4600b85f2ebb2108961f61347a51ece5dc8acbac290f3e91cab25b98df0d6c351f5d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dd980e6d051f905ea51f36743388b1c13e9ee2fad24ee45fdbb65bba9491ff866beebec5b945085d85d23fb06ce43696a95bb848583dc16789488ff2560006dfd8f4ca25806ae6d3749a226e4e6b8f6fe51b9f66183bf14576e7b7e934c125ae95d12baf834c8c5072b2d36b364187b53e511b799a7ed467cd6c2d7a7aa2c97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67c73bb343998d807df0b1448f9326211d21a334ff6e67a4ab54e8fd371ed31af919521bac911ffa621577eb8a03248f62be0da75275f166599a98115f253bd4ad520222dac5926d2607617d3e3cee0575ae6534b1501010ebe1d9b49df199bf87c90a751426fd4fd8b026cdb505fdd49ee454f0596361aef6c227c7d377c582;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68fc375d52f3edf6954f69ac777b0dc959807234f51850da9a57f8d8f43e02e4d739d17ef1ae99d900c43008d7dd1c72533cebe882731fa4b0c6a8f4aa04379dd8a8e72f85065a8197a7fe55bf668c770682de5dd0b18903cf0d1453331ca323cc990d1f30738ec004b956c1982dc8f16f9a47d9e107fe70bb87863d23555869;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1a05a39db8261dd2f1c4bbdb99f9d84b149e7fd61708ecebcf2ab3acbec7b9d66ede3b1f84cb74a0ad20abb0aae29991b8dd658e58b0b944b46175b52442383b250b85d556e2b45263c86f1643f762cc344223dda0e20efa005881883859c55f805886b1a6344c86c7ffb2dff3c6df97f5178e6224313b4000dec3fdedd38e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6ea3b023f868c4a2e2d7e61c1d4323c44cfe4659f07c1c1d09a07438488f03abda340925d503c8ade9d09aa88df9170d7b8b68a4d6a5b275105bcae1508578ad4e5cc1440d48fca46137758c79def6931b37c933c59852ec3eb5341d56b1c0edb7c96bf52aca3c6ceabd53a05fd161f3b743dae969958fdde4db7951befcca4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda197150aec1e80c03af4e5f1612c11390b99f6845e96eba267036dbb3130dbac47d0d836720231432b3dfae2b68a57eabcc1f0e38916a47910b3d757510fe2d3ebc2711a46582e7fda5a78012295d7241529bcf920cfc819dbfca92408dcb4f73c3b19f9b209e8f200403ade527b4536a0cdea3e0ef1ceab1155d4d8b601578;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec66360c8db0e60e3d7d337ab2ecac719d2a97d32e8687a4e8971b995de86ac7147e6c8f0ed3f731b235c306c1f6372e267a6713f54ae3df71491de645c249b1f8382a8216c0054fabf6e2fdfee79731632362c2404a2288aeb1c4995e376780ed7727366378105cfb37936cd7caae0ed78fd1fa786e9cf87f00a69f7db444b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3de11ea9596eb62d64e51f9fca52d119af34bbdd3c43ecdf2e19bad16a4993ccc8a3c9939af7649b66ec01bd18b00b77e388d053532b943b9c2c8b4472571a18eebba908c54fa43fd6f41db5bacec14ac23c94d2720ff72c98f95a3eadcc9149823e29e90c268694550ecd280b7b5372551b2927e0db10da1a287d356b98dedc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he64ff91c0f55e8fcd8b150960fbaed81db34f7e8cc9fa4d8818d24909588413a5fdd5519ebc2146532fbcd113288524bc31721d1d09c013bb0ba7a3c08aceb2104f3a58b7876a3504614137929a034177b71879ffe5678b69c303c612074656f8087cb5571e63db939f8312d03b3c484e81093a5f0f96fe88b1d6cdf99c61ad5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49beffa3d4072597e12ab7e689933f8785ab5232e49ae39db330965a1f30b50fd025ca1ed76e5af3adc0ea2800df4281cbd344996c1de235b750e8d41527146c3c69a7c8d690a72f5ca4ad683cffb96b4a99107e6cc3dec036d9cb27262732bfc20787361110d985c2377e9811574a2937898d781631bb35aa112ce2b3c89780;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h128ec0cf70fca9bffe44651613e350804d88c870bbe7e83a1a27fa707c6ab8adfdbbc8a372fd4fb8f41272e25a8f602a86962c62eb77c711d188fc161d98ab306de103eebe9fc8dc3b6b4a39e284ee439121cd1dde268b2195598359878adf1d21f0e2503eb8d647754b867f4a65ee174ecf627bd78f98bf121db229e7ed089a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf61ecf62fdd0ec5da2dfbd7f0452bd02481abcfed753065dda26ebb22479526cbfb8eb71ad1edeb0f218a3de72afc9a584fe7f4efbb20fb32d293af99f803a21659c447c20b336f9da618b2a0099b9c1dc3243e59f55935597a8f24719fae5e8c7ac95e8d55132ceff83148a43da80df85a8804e193ad019e167e466782b2ce4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c3e34eff8ad40b7b4a849e56ddc5345a5bd5e4e3f47e70df34a91caf599fd3f0f43755989eb9e8f6c09cadf157f0bbb77884dea0b955ea0e77ceae6642a4fa321966f6b34ef2d26be8f84da5785ab2d5976838b73b935a972bf0b15f500742184df9bf0d96fe3dc928c3091b0a5065d0b23e344dd69802c2d55ca24305e1854;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf3d1712b86662f554d6a7456060ebeb26fe7517c84bd5429bc2e8504daff037a445aa50df7d59362931dbd9ad57a97d830b127a4195cac3ae3d2063c2897be242e692488429547a8f5c614bb7ef655b84b14cd17fd6cdf0895a26f7469d157fbdfee7861cb5bf2bcc7911fe558981c6307ed3d0c85c6ec68d383332d3e36fc9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe2fd3074e407f397ef19ad5d75d20e69900dc9d1a2882bf94f8a4116ef24472ab7298082530a25277da5aca7b7e06d87da81dcb162b145b134bcd24bb291f289a754fc741a11195a88da3cad7d9d9c607fbab33c9c3cd870c13076d31b09c373559efccead485d5bc7d76cb01a4445dea402bcd7149e3c5e7adbba6bc001fdb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h814355f31937e7779b908618c03a73682ad1e5c6d6560a5b6e281c8bd6ab75adc6c257bd6518232013b5d3ea8e2f4913320f328f5b7c150e10d3546f642e8402f78d1baa3e07d5387b811a2d2beb42c594d4b2af206bce24fec97e801cc589f19545c5fee23cccb0447786369f6c832f65c6426bcba647a075f81bdee4c54ceb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d955c698959d2645b3715768bd2ca702fbec8888fd86e1e19c128f9b25f6c1c48cb9b35313adcb9cb1c202fd56de574d8e6423e90d7defb9956e94900802c007523a9bb053fe6ca7d863e586703df5b3194930f37c4c4179d928fa4b1f0f56592dc7fbb43ecc57d5e61702f012ae196be24d4a81610d9cdb5f304648709e44d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd02ec69621c56646f0692891f5160c257d73f4368f2937e1feff940014e9137328491d63562c256a943fdcebf3222aa7db0f5edca31dfc4db4998bff2cf49fe159c096a7a6c45d30d6440bae6eb41ed43f80531abda1671080edc4b2e49cce740514cbad832641c6b9fc185776f388b52b977e64f7d9697f8fe1f866c090ce2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6937d23ac19a9bad3d6a3318fcbd6d504ea5ca1cfe2055f406122198bf62efc53cffcac1f96b6795d8ca0a372b284b642e4decd9f4482edf5205bbc7adf690693232508f0f1e666b0ac4c8713525027d9939e0ba43dd423c057f899adbd21e09f4fa9d3f2d4327d5aaa6b07df07ab9f79078b3b1201da3cb566b74b423e0b457;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d29292fdf1ecf15cf1a1c25984b37e9736cb7570382264c96ee4d1f9dc2a05026d28484fc9ae5391b58dd984002406fd63843ae075745d499420efcd942cfc9fdf47c912eb221043d0d8015782f4763dee56e2df998ac6ed40ed568eb8a6b216a500efbdeec60dde754b6f092d9bdb88f5d3d950e3758de5cb56128523aabc4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10cfe02d7b08c2bea3f32722d2fe10c20a531e3b4aaf9f5e3756feb4d3e1d452155f7bac53490aba1f73b73f56c450f29764c4f7ae79197e77f4f6abee28fafac9d7b5b09b73f87bf09031447d89ffbb60a599cc1eb95df8391da5e9e4332fef50265cc5c3313485e7fa48dcba1e9a1a93b6c805581cab1b91fbf44cfe711aa5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fc19431874933c5b8eca0405fb666671d2566969e03bb9e6f6c26962478b0faf380147f9eaa9d58e56e80c1d51c10257394f4109085b8a55fa559a3f1831762594f384b04be996c04db4d2c3535c0b814789007ca46ca83a99dcc5ec40b6625d701bf4fc400572a135e27ee2d500327d90c65b82e0d50871906e6a337ae57c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf6155bc0a4699a8cba3ee5350426f31e012ba1a152b6bbe608358b5b86a331733815c5e618da1f4badf867be5ab52b04b2a910a7f649a92633815fdf7162073a7804a638d9705f31dcd865ac45d3db60106bce6e183451e472052afc607187c58ca74ad173d1fcc5796e9fa1405dfe213b72ec87408c0c0a1eee708e23dd02d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8df249f192aebc65ee4ba48d31c169f0d6b75282b77274fb1e821440d71ec9c4751beeab506800b97c6b64bcb4a83826d0d32c551010a8c1ce817cc4d50dae3eeaddb1f51cb7d696ba67283fa29d568ae52518645469d153e2a1100505f39d71874e0b2751ec40c9f49ca3e05b7d6b836fbe98b1ef425527dcf6877f2fc4c5c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83fe773b90bc08515a615a33762622c67cca8a0ebae56888b27287d0e3d2cd0586b950e6a0b896dc227ceeed32aa278a40770e421d17c1f14f69075f6a282f6c1dfb1e9668fac47cb3b6d07f380d57c5d6318fae2df0a58acfd75bda6d23ae24c50cbd2b5e817a3c9f252a49959fe97cb0ad68db8d935f0d606cf70b89fa8dda;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0b1d0c3b3eb4c94f14417df194b5976eb46f91351035beaa176e7c619e5835799d0b1aa977c9181e4419e642bf1c8689f22a3fd6c9b079468aa91a84733ec650d892b0202a7d699b07f447f90222cd4df3c32bfc7f4fed02ef1f8b08924597977d349e4fd6c9815dc80d52ab3040aec7d80601115f7d66406b33eace2226f6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd15f6d3bdd3f20470976938b502c43e523131b31a8d9028fdb9f5cf33e618740c34dcd68fa6ced94344f61504911b4ce3c24da5c175a71f40f3cd21529ca21dbf226bbd09ad25569ee749139bf9e53cc9c8526be021f488ad3b549b33184c7119757eaf8124c74a60bbdd0817c4fb49efa8c022d2fbd477f171b76036089677;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ca474529fb067b80119e9fc926b0848b3e30fc77a7671d0a7bf00f184cf27024052a3b221183e3ae6778cebcb2e41f375841ca6ea34e08234e488a4fbf1d91f8e0ac213b4730b1dd8619c9a4f3c685ab0612cb8563e8a81f8306fb50da85279718c2d376932a6f545e24d06d6ddce76c7c8ed03b8ad6008835e30c962fe9701;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22ce12ed896a978dde39d596c4a9a41629f9b27ead91956b07d3409481f361a9eae9395d8f2354f2f728c6b626eba2989e1e1de5973b15f9b7d0f195dc9d6d7daf8601cfbeb54e0b5bae9ceb5d9d0053f20e18e9cc23fe77aa97d81eae577700fd57c1735f33dc830beded24533d38af7934d5c71dfb2b404c8c44fbb3b43235;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2079d83ef3f503d6bd0ae0cdcda6433cb8eb527fbdb02f747b7c3b3bfc20bd76ff6aa7b4a40b20e9e4847df6a1afbe83d8333a5e484f39f416daaceb9c81a7611039b639377e6ed9ac5fd601d9c35c4c55c90ac6f91cff058ae840d55a21de1828aaadbff4cf517a0ef6ffe7ac2bc237b7b445b375e84a531258206b868ce2de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37b3b9273c54c04685d0d0da667cbd8651b38f04858b8df01bba4c8b56b7145d40835172277a99c74b47501db26a98df894f6e523c575dee04f3b7ea998dc274a5671fa5780de1598aeb4a4af2e64e47ded51d3e055074018a64edc1c25121e17ee0f67b62b8eb20c297dbdcfc963202ebe83b78210afb432f9e3212ec035e1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41bdeec731f749718f5464f1028a15a23e8abd09f00934a1f4d431e0372a20ab9cc15bf348295c354df204e7530022562488c8b101606a6311a0a2fb076262ae86f20cf01415629487081d0619c375045b1107f6c8165521824237aa3d4f775ab190f400f135ae0740ad9202dd028d5ba9b734a01e27276b24684ba62be92edf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd3d6c7436bc61e37b59bb2f9aa74bf93b6454971d135916d075988ce3e5a6825d568c597b7391ccf4d5c7821d7a677ec06b44cbfb08e9e272fdf2096aafeaf4250816886b7848a5231a3c81be8d31b009235502a0c4e3ce431ff7239fd43adeb17d80698a8dcdc4a75e0725f2b4b8a927abdaa0ae8487856978b4ceb0be482;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61f93aec58efdd2d0a4acadf73675485ffbb28b533fd19f228989a1b02ff3c08e0752330ed96d8850df117e88106814e7f574fa6dfb17bc30c0c9f0a5e23e8653806234568b220d8e71131e56e610b137933d6a5015f08e6daa77d396a684be6c42f2de83e6ded26d94a1da7c8ff04ad71260d923ca9e12ada1e1d548d83205a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31957737ee3ce061ac73d62ca036b1fdf9aa59ace93c6f151ab74d6fb7f35588d40b2e52263f1bd3f7feb47cbe28dfa1597f279a00fd6f0c6e258a8287856f00c2521b8902059c97c65fd965614e56c95f9506723b0653c9d0887fe6a88bb9127420617d6ecc25dc1277039f9a5db43e6eea0027c7f1a2fb9d8f6ce9d7a39d97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9f1da318b9a4d82dc3e9fa6461876bdd5b82e5fec7bcdfed80605ba7a94b66d30ffb13560477726f9b8796ac39056ba37cff65cf869a6e51a59c415fe4bced1eb3a99333923bca233f901bc4f04a6be498dc0523017f13e136fef8146c8c26331a1b838ae21a767ee0ad15bc1e2f124a44f870fe8448a54eeb2b1657c549a20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeff48cbc2342093725b52e89e44485f3fbb197a886b94ebb5079a0ad7a7af7550b60c68731099d3a1f61cf9f19a5e10b96995c1bd551b6db2b83920fe5bd51f343b3c443c2dd14f6ec0ac42d9927977f30284a5c435afe4b9db8c84a024aed41f27e3bfa04bf2c74f43101f00bd6b5cffa0de38c3ffd49b45d0b16b0256dda9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c368e2526250bdee0c878f48ded18101e949740c88f953387357df34f086ca0f5c94bd5a75fb3d87dd277bb37ff2bd5b5be0850457399e64f64c1a9f9d50a14accca0e56346d53badaa9f20b21901ba3b037ca494e25e365afa527c77e0620c5f0f58ec054087c7125e229c2c903cc575c21a449c84ce20254f7fd4f3514162;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf24c23a1bee2b2a8c6d46b1789b2940e02a9a6e5becdf26fe6679bb796f1bef1ef6a0afdb17d113a19570db7df51415321245b2765bd99894d1b1620734d3af026a3bded992cf0dc6410850031c65fa616b96c60ad7fb2221df740a3b8b80a306465df64c1050b3a18dad28f5931e806d1ead59aa94c60b42eae4a616f915cad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5451dbc582722e50f8b28d3152f95d8b66cdc7967258dee261967e31635bdd1b722d2b58f33e94dbe65e45a9daa17e8249a3bd724b93130fb336fcd750f8fbe3f2590f62115a840c4f9a7806e7f4ba0c20690ca7bbe4fc34bea1c0bdc86b78898ae6700bf5f0f879b690fcc1f28d9edc815523e950147aa7da33713c4fa5d15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h405b78e58218a48c0d91002a1a5aa7a26eea06ac8efe405c9f26d55b54634d30557573cd37070e42559a26f7fdfacda8a23cee43711e49f1cf4a3dffc1e361345d3f9e687157509701ce7625567fd52e035af3949cab252c684db623204476d110a29a2e690e8a7d3d7a5abfb114de3910de41446c906695fae9dd89c2d232b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3af89a07e45643cc3eb4c949bd1decff2162135ab6796ebd5f4be86f02c83e9e4c27fe173c047fb1f858e990468564621a6bb1bc32212b9afead1792a8d0c9c2834e5b4b7903444c382b196bdf824468f6aa9fd5361ca18365226f01aeb86eba437d3d745983e14531427b8116940c2d841bbf8bbe00ddbfd711445aa8033e0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89cda83c66f05a0b3d31626c9685c114c7ea638620d83caefaecc1a628207be31e19c6f65b7ee817b77862caf1072dd36cdbc330950c3593c458c39d7c9dd28f87ae20ddb71a69e8ddf8b287e426b41a9b36eabdc6780bfc7f1584ed22fa1471f0cf8a4e4b7813425288c2341e5a316f206be74e77ba42dc88af383d8aef6c97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7ed2329e7375eb466fc7b5747e1ba6134d44717c3de7785afe45afd464f42921e442d456506092f5c5c041def8a18d580accdd49a975cb1438be415975084d2be944a2dde09bb5d905cd2c48db3098d2c968a9e4f11ab49ef212d6ef8bd8a01f47513693a04b863729aa5c7e6bf1a91503633d1081e7987d72ed48c11a1914b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60d530b2d9455aedb717fddb5100d43b163ff54b975a8bcec3920b66108467496424cd72152ce6d96eeb277226a32a50c5fc385b508eddbdf3e1d5194565ca2349a0af73c60cded13662ec1a67849d6f21817882f5896e794f5cf6407af9fee1e7fc4599c01cee172ba29fb41dd3b79a81b30d1ad81b29d4f66d8d864ceb9b69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h346b5d70f35fb5ae22a26f3107ab648130e9ea5f17480c069a21771cdced3360026185abb75a64b9ca82638d94b606bff681a0a67ccfaefc3ff9ecf86071fcf8fd6e1944e217250e571110f8b5fb9b05bff495718c2f191a4b9ca7e0ec1a0cf12843cf8f501f31d5b0df5688eebe72011f23fbb0d7791b6e02d766f73829ca7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5740aa48f28b73d43303e11f828e2ca5230f5e50bda89e34528eac5ae98f7feb4cf82289faf41d79c354e3b31c8f9a5d9d44735f408a51102d5cf495e09ef0a0fda94874f09ff8b2796b2791bb3d2af4d1d82aba2edbe5c97754ae86ee7fd7db76cb7397c96f2d78e212478d9859acec5f7c8bd004cf5b64b912e707e6d789d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d138c19465de064e31c03113c91b4c4d206be6e007c8828bd56bdf94b20a023424d2e68022da898ec4bb15a6d28a3f23a4354184ee2cbae7c64b021053c37fe39a2feef63beffa43309d52c4f7970b320f24529fcef7535bb6ac80fcab10c23ba92749b5d440cbc41ebae5b86edefcf381d209dfc321db195bba2788ea844d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e4dcd5956560da1d70fc435773475ed212157972e9fca8537be42561fca4e5e2aa0707292c4a4e2c9ac98cbae9871ee2db278771e7f783df69588a1b0187f6abe572ca4c65ac73b9b4e3a22b71d4650055676734edd7d075a95d7e5e4e2b8867dd7ad1b51f92a274963c53ccd579ea0df89d4612e47f64afc46fca5a74fc0bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hded1bc5abd6ace938b8ea7b6eb879eb86e52b29af0ec77e76080a81adbb89635b10f0f24140247eafeafe67c27f4eab8179295fe30e2deb6c2003844ab81a0dd7534dc740ab58cccb2c90cf2908346c09c2ec854ba5753eb997788916db8f6ae0bf361d4e69e6b66933cf3d24dbc375217af6d2459ade79d82be7d3efc6ba399;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49a002a3bb423d5d1eb5e0440ca9b5d045e9022926a3c780899201667cbbd2aa5668b73c8dbe6b71ac5b6cccb2ff01c0df0054d1839bd60c9f12d59021dcc1efcd99c3ed6f3d69ca11ac2d8fb078886fa44755efa1cdf1db62bc0a19b09fb9322cd06c8a795e2c7d7f4167bee9bdecc792393ab9b75fefad674f4d2de37d7ac2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a5a14eba47ac1c2f2f05dd42b4e977882ee55cff9a6a17edcd1e6ccab4ee015ed13d311ca2f549c19a57f52a69b628f0f89dbe270bc9ba43eba9f5166c3511d6e9c6cc14c02b43d7282e35270887c8cc45f08fc3d23de1f8d706db8c889220be5ff2e978ffba12279d2e0a722b41baae4402d37927846eb875aaee879d067cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he29af9ce7f6659415710fa0639d83a402da89aa3e485a97049193873f7a2b634c445eacc4d970cda970cc1b9e16138cbdc4f6e327aee8f26c6519e7b5488e34634defda95212f1066e7d14d6accebff27d0c0ae6574039a764348a4606ed6c01ede2d65f984d101a4cf7e709f8f99702a0d6bc5da73ea1e09614a861208585e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4cc6c23f289b3595b0d7ae64cb4d0c8a5b84508c5f0e42c2d4e120fa36e0fccaa474fc6ccd5fd8087cc318b68f9ac6829f3934850a95cd356261e65073e65b283de79650f7646a9e930840e8b8213bc759fcc8394ba92143ea4f9bcb07891c37cd63c8106ec9957a3e2b3297ec7b80ad837271b0b6aa68603141239fc062f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40288ecc9948da517755945444e8aaf609c8494ab0c1ccd61942a71828da09955c45d91d21be9aa7c6d568db87082c1430892800b4c351a861bd23d73e59016f7bd8bb567701936065932d555e7b9e61c48188a31d94e9b86195414eb63c03fb041cf5e0448a4a39271187737992f34874d61494230a5579aa7783b58e8e57c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha932fdd0a9293c4253b81e291f722e8de021a5f5b9774bef32e6128895fa5f0da99739476ed7e3074b9dbf978c11f2e73b56ae8d7522651f0b3bf035de4df76459e17051a51f936b6a94f57843d60d5371744e894c11450a328dc398478a304c3f23c69a6a83a29ecce73ab7085cdf166ad0e016c9ea51314fb2ba8975428d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97a21b976e13cba220612bcaf3be1b4b28bdaf0703e7c1099c3cc95ce95bff68619d201246da47f08be3419e7029c0daca60bc8b619ebf6155c8660ae2a999a282c2bfea03e0507a8afa0a1dc2ee746dee0ac0619c87f953fa98e7ed8a76cebec268b0c7129157b856f685746fc06c53ed23f2b5e104fd06ab506ee6dcc440f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe88bd4688e49222db1dd6c6eaaf682cc790d12286fcde750c0dc718bf87e4cd79576eeb3bdda0ea25dfecc582c2cb59757d7a3a0b3d875d2da78d9992891d31afd99f5495cb5dce47ba12cd8bcc5a4390cc99b65c4ed9061112c0f8f823888016bebf7ba73e00094403d2965b7b64c305300a159cc474f6196169ee8cef5872;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd170cef905bfbd676606348688820f2f74d6d41f43ae7e61ece18feefb8e664ba5294791f5c798e9cef8befc06487dc9845e3f0b180a88b452cab616ef5946d106a501bc88287e0bb88eeec5db75417a09bfff2f910b873b96211fdb5bc80f46d6683ff8e5c9ce0238eb5c0f31e42f58660681018c975fd42423a8398d499b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bd5201caad997b2179975ed758cbe216b5ae1ec21c699c789b0dc610c62a7e8519d952d28cd4e768ee89a719af093f22d096b172c4f11e5e882f7d188388fd8563d6be710f224caeaaf64591c60c2939db2b4030b7f9733eb1ec16815726b5e2ef71b31d11d63d213b5b3cc70d4747a197780fca7e641c222813688ab2e8ab0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f96e94e4fe71d7941f0afad0f1489c6eb440a017c5f3b9ada1b1be769178bed139df002b59021227690fde1b9f0b786daff1e7057d46b6033b9a512f3134dd7c29491599d3af0f4dd44bc4384d45c8db9ccd4a0676ecb1ab2dbf225c04441dceaaa4a24c6e0b2954d9ffaf1da45ccbda0a5efddbf6d9f29e7297285194479b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4199a55ce7d6632ca47a76e69f9a65db9f51110797b7f4d150bc67cfaca1e5d5aecda1fd255060b59ec27736ec8a6683b4a31cb094cc079cb72733ff45e825c7dbe230ef2edcaea9c5abd99041bcc1d1e87d489d85cbd6af4bfb28654b807374bfef73425f5887b56ee27253ddd2f60816fd901c56e438802061ff2aa9ecd662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8beb2fed02b75e5396904a043c4dbfcce360e834b7f90873e8e9b245b496fced86e3ce027657d4d98c4279d5aaa02b7f5f564b71711126f3bf5310aada39d59939fd5c441facdf6ae069aa8ac13a5400d183ff5173f27891599f3de5a01330bec1a61844a3ae11dceb5cdb96b6d4a1b646d580a19d325a111969f61dbc2b16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb70d76f86908a7aeed67009b59f8ccd558e1022a5280452c0839800bac4c8cb99143bdc858380b953b138e4ddb73ecfcc8d4bb4db75359a473f3fd3b4379f26da43cf8d00593d791fc39d447e26659d6ca7b1ef466d5396e8581112a58f6bbccf77cbb117c47a9d02e83ec586adcac932751140e7072b55548a0388fc8f7c948;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d9a91be2b6b859c7dcdfb6fcb421af78513fe40e82938be0dacb56804d5fd8a8a6ea9718d083073871dc99ad79a4fd7537ce7c1c28b1bbd872c7ad21ecda799f1789667f88aa5773b49136730fc36bc4d2d2fee9698da7fcdc718db59fcaadcd9ad6a78802e350f11c7ecb23b481dfdf77b77d16964a78f9164ada2fe924422;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h735e4235b6fc919c705e1a8b53b8b0224f0c441d4de15cdc9edd0f2b6acfa4c1456852f39224fbe0023a2202f3df69034e04406100ea1fa87e9b771fd7dc69a85f95ecf064188628c658253e134c59f0388305f0e28d76d0ff6f45c7d93df2fdd23b8cb10216131b0dd07ab1da836aa8ed2f6659d85095620388c828dbfff4c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcee08eae914a8cb5489288175dbc8504af20176470f2d2a8bafcc7f7ce8e965eb2165736825580be3cb535faf39ef6db178e07d5786ff178c27ef8ead7c68dd8026f7487912f67907a0e65f91eff4943f6c42679f360a1030a1ba5ee1650ad34b03cd1c9b8f7c93a64524c52f0db2198bfeb9a237dbd7e86a0e576ccd39b12c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51992ea8d81703631e0a1b5048b84f258e4a064a125132f036cfb2f125002a443e1b720898a1be574ba74501a65e1265be52500a6ee0aa0e352a78f42180a12b5cd804df4b0b29b73a1b1e9d567b6c11f5c8d67d290133e53efb87e62794f19529ee6f59919fb3db8401d51f7b706c5ef623d8f5ecc4c4bd52d3ec9e56394975;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81e70c21c7bdee346328e3c1c9bd9c1fa8b50b6daabc21627294289f2bc8c32b362f6073b593b1326e5038e134b3d1f81aee6a515c74f2384bb003515c36fd7428a75972d995b511f76fa3dfdabf97ae54aecb1f6aa189a0b6d20c534a05face9a69967429d3583869453cf0f714bcd90538e54c655aca2adac9c88bae422701;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a185d7a7e0f6da8d917f3ab6d0d656d59ddb91a0c9650ec008520de8e6f47a1222bcae0a9196ab623b7bd46e3b7f6a6d39e6789e12290dc2a506dde10a7bc5dde252279927be831974afa5aff8ae747fac0fe1a060d6203f3360d4d81f7570adb46ff309a2708a82a523fd6343aa943dc6696f22e3379c5e9def4e5c105cdb8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64251c91931deb3f37fe0e80e5bbd77325946166bfc0d213c9d8cc75927cfa5e8bc1045b6aea2212b560c97bbf4450692f895ac375c409a56c020f5a17c7242f37b7188060bf831969daa0709301aad9200a2ea9a3c17084efb3295f524ae18018e51bb654386bd2dd0d3b703d7147edca5e6e5ed12f97e59a473bf934ae94d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8663001b5069736bfcdcabc2e03a5e947722bdded09c7d888e925dfb856f5fb94c343bcdf44b90429fab9d65a85268216bdf0aacea72f0aad7f10f75fad1ce9e0e34c4dd177565dedb8ceebf030b857fad460290273a9c885c3e19e1205223cdaf9c1caefcbb053e700f2b2008db7494ffd83a136ecb3d45a8c192094fdb450;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h310113af69b40ab85e0bae89940a4a754b59a72c3058a6f232195dd8151e596dd7192103216f1b646c34fa0923a545957cb5f28683ce2beee89161e9a2d0cd2882440f2ccaa7e6add26aaed514c38f10de4b5606478f076dc3aab30853849a222c7f052e06278bda1a386f8864f7d6ccbc24e36d9a245fbf5e74851b38ceac1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94b4946a287ab1d6bd355382f76a378fe75360f83eff9fedc1e9e6477eabe40f0c2ada867dff81c6609a9a0ca2a2587c6310a44fca439fc843bcf271a8d5bd9e7a42e7c257837da4770ea8fb8520c5bbedd962e6e38920317ba980473919ba19c9f5a9da0094743eea0bf699a7987e30c62e5411bd7735cd0f0b1583160d1390;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5088423dca783560af0811b0021aa700f9b6aaa46b4da1c5de28ed9366c82485198ce5c8fbdb53528f02fbd48e7bb1a9465ba2920d19239d1c95e5c52500d14deec2bc98a13bae27479d6b6b2e21483449eb5c0cd8fb97a5a39ed7779ada0f3e068220d56e8547b79ca8841e5be80d031db3c5092cde258f5820d2465a82f7bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f0e14545800ba0c6f0983eefdccde14b36b69aa8adc73e23cf6ce19589819ce744133219397e210da3ccaf776c016775b95654f6ef1d5d040b215b984d2093017b1c71d28942876cba6b14aef9932d790cec1619f2ee1b5e8f0d0f42da53a4d959668cd905ad074ff83e76cbe5263c31f0b6a0dba7d4433173b0875b1c1ff49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e5705a60c1a7086da0aef736d84ccb9e882ab245fa6e8e0dda9d37570fdc74b70fa0d7edf0abc93002fb6e0e359da6ffe1c6868924b345c275fcf9193ffaa148fbc8a4114fe3b03257f4870a4035bcd0f3873b78a572d1c9aab2ceed8ca6fb423f70022d5ad55084f73ba52f9d9a79ff4691e25a67fa81b25828b1657078611;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37d0cfb7499c7347c4fdcda2de2e829b07b18a1e7196f636790420affaadb2feeffaf5b8072afd97bfc11ba74ec58024c073dcaddde511ff5f02124e48201f0f0adf1b2d3309d0ee45c58e0cfe4eaca8ea4be11e0794ca47b48cb3a69372b8ed7123e0df127f1427b9f590242d872e94f3e206f4ae3623796a974e454746dc7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd788748e0727e809b43568d323ceedc3495286f371ebb81c139a18da024011398eca3c5d8001808d26eeb7a58349de5cf09f63518be358a8ab3117d78a31674136e63a04d00daad8d7f9ba4b7f360966b92731ab0fcb56c523815038bf52ff70ee1c8419b3f3169e13be43718b9f10ffa768f97025e4ec696d73d5ca5ea4771d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6945feefb35b57db0726f0659f4df6abecbcf687594fa9ff52c49f52b847a63a91d78b22f7fc5408acdd53b7d69127ee38a550beeaaf0935cec2fb9e818435fdfd62a2f4138eac275f5367ce4abc868296f84cecc4d0f51c8b2714481b892bdb8a4ee96b59cff70476f5b518c41878a71dfc20c991675e697eaa2969991db9b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51895e69041977e5caf2c698b97ca892a356310cbdffa1e320a558ae618c748e78489f00e8a3ceed89654ebe43414cc2e0a57708f3096fbdba4d41a76edce244f012f6218f2d7cbdbe57e4ec9ef7c244f3a86175b5b3b901b8a1857f0e1a077755c96ec25f39b0203c6bd32238b50e9e9c359e8e554cb0dfb82d1eee903e9e47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb1ebeff1426ea5d3c1fb574c28b25196e0976c81d090c74af1f1a4f99aa7fb0a13f56c3c10a776762476b78a74a96b471cdfc019257ce773c3aca62e175d0c6345c038cb66174c2eb04ffce345925f3067214ad0eceafdc13908e573cd93392528b83d9963290a9978fc36a7a1c51fe44f9e949368372eee8198a85e0997aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha879d8ca0fdc9a334eef3996522b3a0064ad5944ff8330a44d03f298c2499bf336eb46e8a57442e10a0a2af15357a82c574b11682e9bf919f8fc6692dd1b7fb9e6790e93d8fe0b6b4dff536fb79d699c58df0789f6ee7d2d6ad94bc9063ef73dae34475295ec675df3933e1ba31371127b4e03b3f3904133fce8cf3a74283d71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d77313a3bca908e1c009617b5c67bab90e5d1fd2ec28cf7549cf12da4ebcc9ea4de94cf5f494d5ac43747368454b84d0568e575b1c19b17eb7a401e0e9b50a8d9b1b69473a40d25d110a11a3d02dfe9896865917e9f4e77c419c3eba4fed7d62312154039faa753fd70d525c08187e6e152d0b1babfcc4db3a185375ab35676;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h321a1b2b8f828701e46785e3a3d8d1edd0c7fe4be2697653778111a743354e6c98089f09df5bca47909f29d83a1c28c97d7e3c0a873cab8669672882984cf20bbaf50770fb2d212cd125173104aabd8e614e72ae5fb81bfca5f4278c13c7df15a70cc3c3941024a6cf6dc612f822fb7c23347cb30d97dcf619a0113339c211be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63de0ec5199ea4ca60391331abc8cebb23e0f02acf036c3bc4e9d6045be200b09c2dbaaac2ccf170cf0dd499f95723881a5c713c1f79496c9e2199e03e1574f2712a8b9de09d891653b3b720a8a2e2b3a90044c7c7cafc66600fc7c9a9997f32909816c1f0a7a102958aebb6f2b0f9349ab264f1c7ed463a3b4fdad7b984380c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5eb2a00a86e2ea73e050356305ad193877a99fa41c6d110373756b9e28c7638825e2f8a8453d451eb66772e5fafb936daf8838b6090ea4ac720041b359c42ffba84d2bb9be2f2f2cfddf70de59d7ffce42e65de6d0990f19e092c8df930c629ee172bac40725140ea5815bc0df3dad20261701c64d5e3929480222489a93a522;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7023416cd6aad7386e57b4215f7dec391c5ce0c5cbd58f0943e56edf1e2d758d610212de270311428a8141d1a506cd5bdb643a718724a31b90774fdd8269308288baf7953cadbdb532f8d72c07a7159cb40b0a7bd84e1f625e9e4843a8e693da3e7d0605945b71922abdc39f8d23316db16f9a39086da9a11a87e48ed446c1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc73f7110349a27b082bd5ef9f061ac42ffcd310d45ec7012a9917aa74e9ed80eb79f881e018706c52cda2cb0ec10f1be107d428bde0d9f23fbaf5f0d7c3c7bd5c21ebff1b9145e566ff8c2d593a63a4afeae208fdc337a33dad4603975593794a38224dfe6d334c23b914cc4e758f5c26a85f26db775a47f1278c4ace42debff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3743dbd3256b81e515047b8d0257f9b1c6707a3a153e23e12b57a6703c5fff7fd971d7d7cc022023f4d4cda9d743148581a1f772df0d34685220ae026c176968024b27db7a7f6ae0bf935ab5c3aef1f13d39dbbb16a4eaee873e0ba6d0786062f24aa50f4ad260193b19901aa81c20718e6d874f205abe4c722f240416530642;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h335809535bad33275bc83dbb5a9e8af0f5d45384b478841558731f4f41e5156a260732485ad75094663f8bd2d05a5da971f3b42323670b340bd8155bae6911ba49c8eb221c61d6b00c570c32f6f761c4e99d4e649535ffbc09e4c4f4bcf5efce12ff7b5e6b6518012512f309d7c572bb4b4be4ed83af407664b18e8da4c2f274;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64ed9ca7f91087f9217193e73943d2059bfa6fad55fd14ff13835a6dcb5ea548f3aac7c80b8bf687296b7fe19f5c5b1a93f51f12d00e1805e487e67990667eab6858348f857312fe9184042ba447ce6b8b14112ec672a7e7e50ba95b72417a50356c0940ea30b896410d176ef275f326758887bfbd648f9644504b23769a5383;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h142fb1627e1f20d90e729aa459c321ff49cd41b5a517024bc65be901ae7755d6fa752d9734c11c99f8743b3bf73537da2ba63a223acaf6b3a61d76a8f3bdb73307f1193661531ac9a1196856ef27699d69e971617b214dc57781240486de9b58180d6cb03b53c7ac3c19850409d148305f1f8acb6e801633259275a4e52abfa5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c8e14da5a01f74cff8c93028bc6c6fb7a4099d592f5b2bf5050169675427d8d77d9113eb99f8193aeeea5b03b44fcfa6f1ebc2aba83f36fb51d65a958515dd453aa4261410e74bfce490f9f7ccb81be639be94e6b2c6f5d31aca3c1384e8b5fdbddab57fdc717f4a1a4032e113106ddcd797cde503ccd361ec8ec272290fb08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h113d9a69e6d15dc898de8f2df0675a695df4506e8ae44d45d4ba29d31f8b56b15449825e9f7e39f0eae084089ada51fc067106108ee4df106f0087eb4f1d78df3ad9c203afc35d7945185e0f9eeca6de75992190250bdb9040c9d2a96b3931e58a8d7e9e05380c7fd738e87bf702bc8825d4d6dde98a85a2cc2bb6aa53696c2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1be803d6c21b4462a625da6cd39cadc03a5959daad5ecafcf3324f286b8784d0a5d3fd8766153e71e4150cde87b0781eb12184b36b220bc53a99dc300a50a5f71e349a3e36437f06112ac96ffd2ba583ea080a30629e4a94b35b7933cc5761ab6878ca3f6e8f5b5bb8c6214d58908f4eeb493e7af79119ab824f75d412b61893;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had3e54a2f7d136b93e73a6577429d7bfb9387d3d41b41a16fd9a086c11438b3639788d3fc3ba41a598a135de47aa973d580809e077c44779ccd0c4ac2f8e83dd166769f8aa849817ec5326620eba217e77a7ed76efadb0e5aa4485153a1ae4cf9dcaca4fbf328c9ec0146d5ce9ca43baef283435c7a823b1d86ef80083936b5e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h475ea37b85bb6fb14e763a89f9af47fa036daf00d09967f7638805be486da307091a98346b4babb607389774a60174cd09f10ca0d20a2afbfbe5922909f1207e7427bc01ceae347bee39f33ea36d84929c8c028c72dea2d62ccf62eb723fd3605a4e9bc0cd26f11deb80cb7cf77b3b9493b041405fda6a9e7225d9475e925b24;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f9339d4d0f3966b92364b8101b9c5498a55b7a39adc29dc6eac7b4f7b412dcb21c103546863b5413a0204c5d81d846c99e5882d8e931e3f9d22b93dc8d989f9a18a55914b5941d27acd913208447ebdae1a805fce35bd975643b16fb263cc58bcbae33e56cc46f367384d5db82a6fb7e55beee45a19d032e59012013eb61123;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e9653634b35712ede939f45ebc4be8ac87c67f8f6ab9049d17793215df7c49fb330f2c5e215b8e78f9ae0097d837b4ebf3eddcfe73093fb0c8fe0dd47ee835bf7d59574110a31fed842d7fe97001be788640d48d239c5f810c250d8cfcf969b2318c30a9e32f33d46ccfe5cf48ff47f512f41f84777f9b354ab32f1d3dc784d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2820743d7c3b6e56ed2647853d426a1dcc693df182c3b06ab3657f3787c445e93dfe02e34cdff6cd8bd13102b28920173346ff77e35cc374a5d91f22f2801fdcb8a1279fe1c8750307b5344f4374b3b125c18193dcf3ed396187567d5d87dcb3dee9d7a460deab856defef5fd5b8aecec996873a4ff08da698dcbaba23d78e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bbcddfc78cf4cdec322c8a0a94902923aed4664e33446ec46cd7bf95fabada87b0925ba2f12aa972bafac7af0696aa5a62d9da5ed65b67009c2a9334a80f849980961c4a6b68eb618226ee4b48c46f403c1f7676c27b89f469285c599acec548c18f69a663839e4b82e637e69d988f9b9d1da36654684e26fbaa6f131f42826;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1194c549c01048e2b9e694ea693e388bfcae48d0ad6a57dfaf0c83bed653bea115fb88fa737cb072218d4694339985a8c2ddf2f267ca8c4d3e7e522a0046c4f4fc0dc5a609602166acca0e9b032f228584c0e01ddc9153df9cd262d23d0e8d4e2e4120c52637e5745a31a7964b6bf305dbff91e3eb2556c4e535c66a39747323;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b947bb351636738f3d9fb7f7d1f42396a0dd4d79db140ae26fcb8585e5b2ce2d8fe01f27fa5027bf194bde2a5d8d8901867c1d1718fdd0a9ced35d183a738b78d1997906288e32976d89866928cf1cb904fdd8ce365fe23b4ae9b5ddcfcac517adc2b0ccdb702ffd24dd6d3587929ddb91157794d3f05349e62c71670a165bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec15f2c9cf0054ac0702332030cad0d6f9510289b9250c770f005410f25c59151d682717bec43b643e69e3669c5a15eca4a60b17190f011706116cd8d16f2d4793b95166e785387818c50b2f46f7aa9a6d64c73790a7d332e355a91e9cf84542a43e49c841ab69cbf3c06a9940ff2e7e0959fbf580d24e847665e49f4a307361;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a6a3f484382d6c52b30e6248120ea0d1e27755a79744714821d1e312aaa153d26e9fe7180e66541fc01cc7825191c40717fa82b99f617fc2d3f648a4c81ccc555a3a05c319d41d5e5127b3d6af9428d8b2b8356f9e0bcd46524efdbea59e8f933c6305336b33819db7490b032a9cbc3709cf9e55f4afe02833dcb3935bb751c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75e4307dd79217aa9de42179919ea4f201e9476d48574a4e938d01c77fed97f6d5a438944976e36fc9d2bb7176bcbda6ef4ba99c3ae5e298a06a11761d3561919ca06c843c87e187cbe812248fca47877313b9aaed5826c7382df90b17aa946e714543c1ab43cabfa362ee5eced13462f150f9cef9b0ee5ce80da0fdf7ee6bea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd60bc0a96564bf023af4c7783ac70e16847be2558c075a6e3c66651202325f8866b9f8a522ac2ba561de3237209f4475636d18fd1300c95d23a32a9419ee6122a8edb09d4ad36c5009e9bab88c282a11f68e650bb6e7a4d24a3cbb96b30fe65902ba7e2daad5cf99d1584969356e1a5f5efb5b05cad5ac4573b6eb73bbbbcf89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d04ca45ec67c3a9c4a5baa6e823426ac65eb23ddede55589065535e075012f2f69d24835871309312c69c51e409eebc4d0dc7ed18ed8fac0095d94b5250887ef6b9fcc7fa375f183520da7f1c42f02e6d82bad9a643f8c0d7f98caacf3fdd67bde1746a48bf6053a018eea41682fed1b8897bc0e8db9eded2e1b7f461d86942;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e6715edd48aa91c3da6108ff43a68f106952bc3325592201476f0df8d566f538ed34b7224f3b205f904729a8b534a136ca80c51bdb89e50696f4c9dbbbf20bd5b11eba682a5221ba1556ac5ee8fa1c416139c7077ef4c898abc1f778d37b3757df016579641a676e8e763a80419191f658556e2181aa765f56c156314d4952d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6d90792f710357e24eebcce48f7c0e62ef0d3891d5ac210bf21b5c3a17ad4b97aa974330cb8fcd921f926d285b5cdcda3f7005fc52075e79fb77e81f9caabd54e9125545a4fc8a796a70bd7b62ea9f296e6367c6eb346e54a80cd3210bc3f8e76418c1b80cce8d72c66b482dce2bc1b58b840a4e798454549dcf09664363981;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h523bdbe08c34fa224569ca9c0697123cfeb122eb4dd1e43bc5954321899b2bb920dd36c4f02588b7f6fbfe68162ae888a461bed065731a5174d7230b7dbbb23792ddd305777a91e4ba5d5243bce552d9d0c5956392bdebb0c39ae96aa41c3fd15cd94afdff9e644f6a254654d13caffdb9e11023a667945273e980eb911257d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33ab26c427c135cb1962c74cc77b3f3f86dc7aa4ff1445965c22ee07e69cb8fdc0f15b97df552712c8c4251f025473a0f52b0b076a4678cf682e54f566d5c014700858639de994725e946abaa3cc11535c142fa9ace6fd88eb1f79a9d5c262248e391e80308d81524c291706e3c0a3ed71108df04067d4f54a15fe8ca45852da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0b2825c9d48c5261740bf3796a687d0f05163e634914a89cd4b588dfd50f6113b094b667a9103dade170f57f49941fc92c80d2f5f5aa7308f41fb6ff67249581b9299c748cd516969fd69893460f9b55fea97e124d2b7f62549f1ddf19faf65eb39811a198809510e6f20182282079265aee6f3f99618f86653e1c94fe56b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfede2a9fb8ffdca76f732a84b1da97a0dd8a4b423816aecc948739e31865c81167f5684c98d6bba2a1a1a2ca734876be704723e64682c8e525d240c0a6ccbc6f9610a65242a9b0fd43f5a84e2fa649790f21d419fa13d50e982d7119739c0adad274f3ba4933e692ffd9901274acb0427a7b9c1f134d5705886bace5698e4ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c1f1ac1ef9263a804134c4255bded121eba67946302d8ea69b329a9ff3520c91e12702f76506d4e26ae263b6d83a8d5aec0f7d9201873f35096b71c1ef4ff5564deac7b90d3515611d5166f66fc788385cf958e4bf2f413245f5c3a0b18d8abaf6e0a963427bd0a8b8d71546d994265616c29fdddc1b3e0470c697e599b0504;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc96e49c13a61c5547ba1c9cf503337457cb1558389e0667ecd19c3a864363fd334b426f884e17db4d7a13199caef2f4f967f1b05e9867a1665b52d4811cd5b8f1e1b4eda7db9d523bdd98d4aa82c25d72beeba1533cdf3e6b3c9081670fee53c321f9f564929d06d92b89f427b153d264d1d67519878fcc1a267b4c545937c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c7a78c7b4e0151272379e8e2891b4df026d56410b543d74617a60ba75a0b9cff767cc8610ca016f44d5e27c7328b8052cb939890947228c80c30a809f85f3b430a88c9931108176c4ca1e353687b2a5486c96cd1e8621f8eee4100b44b6105cfd228fe1d5ecbaa8ec775efc57510e749d56ecd071e3c2a475f1c8dd3838c8c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h139005eb7a1d3959c4208ae8863945ed852ddd7001841dcc2e3457b1aa5f555b543c3cf07d9fead9c3a25d850f3dd4f8d0916a42538866e4b2148dfb71709a95633fc1b8b2a9dda665f532415af140ffc90af76a35754c73a9bf6f5ef1c137dbbdfbc4ecd236969d77e71e1d89120a80bc870f1514502508b3f00dda1b5e5d11;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6da4c83c5b456066b2cfbc11f9148dec1c138f9f5c75b399ec3be1519b5d6e61ac75a882a3b9b6c6692b793897fc2a752541f92e20d818c73964e03d3231e9b99cd0b892b2e64ac5a57577afaca4a2c1606478f10de3a51005d0754da1fe01d5b8913df4ee8ace7421221adaefb63a67a2d095f3da0a2e61b449196501bb77f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47526e2ccf206eeccef7e60ed2a89f5b0cc5a64b1c4d8681527e01143eef799c92ab3e7aba43e4f74368f4c1897dc8c537639144eeaf58e983332dcccdf30749ba868c62b53464223a27f4572bb5a5d6e94cb37b44e46379e2e616dbf90705a2a62b64374bd2ec7379e8ac29df71cf6c9f529fd0f853d4dc2db1de9b6daaff05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc1d9b575e5b1a2f8627baf522f338b3a015e87113d541e77452bb681c8f1880bdf2b50ace974ed1b7c5fd17829c1c913a19a1f965290e2e7fdbc569a5568d90442e5fbc7630e189945344d5898f4d54fd61b17ea4edf85733093dc012322491951d5aacaaf18f6014e0f04629d3e40f8c14917e8b20195595abdb5bcd866187;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10af08abfd9f0ec7ebaf0fb5f2acba5e9be1750355028bf818213b671b0a374f52321080ac4ceeb70db683550449ed08a6b576c33855888055373edb52e2e7002f047278f2fe466a95022bbd76ec95d626bde2382e731c20eef77677a2e767dffda53d4c18391882ef1ca94dfe0a4c9ed5d4594c2babf471d94486f0e96c109c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h553abd45bab017bd5570f56db026bf2a777435e61d9abbfceb168db145d409de9e229bb96313d57be4f59916dc9e0ffc356effbb7e3d6d0b0669b3dc1e072f4b02afa326324f1097c7daa5124ee3a75e9da7c06a32b049b2518c8260c624e193606aaa4f19f883b4b0c09767999b1da7edc534f37551175f4e3c29ea886f9e51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h789b9840a449fcd3a08a7686e5ca1cc0de5d795c0626a63834a079f55502e94b8bc914188aafeb4a303708212d07c35699093e17d709333399f7e93bfd42ef72dd500da18670d2c0b3e48784481ef5d6deca9726b03a29177a5815abe78da811f009bb7ed496e8630440a0268d9c66b335b36e239793ec1eaf16ef5a857747df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3d4f30600f1e122c30e65793ccd29b908e9ea8e0562ff11c6572863f8f1081bf7c29384a2dd464f95b21f02ce73cbea92662abc3346f002c4f9f49beb45d39de3b53e6f8c78431d35bb8e9517be56d12a5d2baedfe3ba72fdb7f79924e9b673a880417856afd52c3d7e858744383eadf2d683a998b91d0cee5c0114c22c1894;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a4fd2bb69243bd8f57c8f836183a523ec3e6e9ff59199d92e3a98359098aa2f3b2c2343f50582147b705e62f7101598bd897f976703fbbb72004a0887be8602f4a86d5da091ebec00fccdb2b736a68b01b5a61175e9f135c0e3b3caaa4c77975527d4d78985dd44f1e138cd5d30ba761605ea509abb183acf6370a1dde042ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8695b14628df0c7899f84ef7bbc5b7c5c73c2dca8d5c2960427ad55f5deddbe0ac84d1c792e40afcd58c74409fc724f5f9cc1e344f869c48f3afd336d0f25ff5faeaafa04ba858ed3b0eb1ba5128baed8bdf1001562ab008082f4e716dd33473cc92feb334c47471cc40be82dcae2a2439cef8267b4fce11608a5b878ca93d89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e085719b56affe062d1dc7a58701927ef9cfc9bcc40ffb091dcfb2ed54b79dc353a5abf68ba56fa5d3bbea636d5df259fc2c94a88df0313e354c4954190d6b0a889c8ba20465494c0c4cef1dbda97a8d147a7d4a029bf4b801c4b34d7fea9b2a05b90a09de493d778e1620780a8d3bd718803ccbc7da3b42beeff935a2009ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce8518aed6d1b80c9b8f9042ca1be58b139671655990a9900103cced4ec52dd2cbf66e92fbbac43c96c9d2dbb6104f04fdfe787ade628e79f759473bd49cb137c6faa6546e8e521c03f677a7dc07ffda9392af69b867add7fd48a9426dfe57cca9188e5454264902d85e5007d9db499495b55bfbad17df8703c693d94f11fbc1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h143d0cc60ba4a8cbdab5a8220d9acfee532aae7938e9161c30f28d05d2d0824826ab33ec1c61f8f880cf641d13795a08302c0b41c7f94bd91b987efd014b141060b95ceb9042d7860a661656682d4ab4b2fe31f5c07533dac0cafb1b65da6273f8946333a6f1da0271d0af46abed56b1f730b7062b8119a0af73a5952e38e6ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0b04f26a858a34afd5d4694bef95ccb9460a857ad39836f8c955aab684093275b8d4317618fc4cb2d40208afee1585de36e67b2d89dc72750beaf5a78428e1da9684e213fdaa554a335a26b8669b05684d91309814641c42b47b2fc44d571d1120cea4c8ce346288d46b66d525ea617ee4ce29a4809e04f851ffbdb5d43143c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c7480798e314bd65c462009ee4ca81f81a7a752caa9612fabcc5592c65ea79b572e48adf2efc51b4f7f1a99b0d762c9a6158f766d61541be8b2ba422a0fb4c88eb7511338dc7ff9516ae7d00c0995b914bda7d461d8e29ca2d69c1aef837772e1cac84743e737460f841d78440b0397ab72bf1e2a6b256f30b205fa74ef15c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f63dbc8cfb96fe4f0ed9947574ee064aee2c7af56aac817f795e5cd1e73a853f29d1641eec08a475c8b6b0fbc01492a13a4451a2c18b74faa2ccb17e738333568d9b27883e513de9cb9f2e8698a4469070ee3ec6700bd7e11d7c02d680e43b1773038f771c027d86027f02c8f729e284fb18953916bf7648d0399c5c1af9d26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c8e981efe25d64f716362ba4c37b612ac57859e963087feb22a3da7bcc537fa8b4663468e5ebbf0fdd1ddcc0dce257c25ada9c96842998c4509533687928220ff0c4411cee2cd42b50de13e4dc4381cb3ca9200c3f6b961e229cd13a118ab3e81743e68dd7f0947f106d7353a8af1e3548b884c5c3969c254d3587b053853f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaefe0e0c1e59027391f826fd2c1b43fe491ea5e1f07c20a095b9a8b5183a6b1237e05c9c27e37212f97a5f2e2bbd097203f91bccb33a4d55a5dd9af571d8adaf7bf83cfb259c989bb98e0de4185b1fb8d3667b248d81847d83cdf7729b67d7a110e6c43076bb198716e6ae551d70e40ebbdf94788de3be3710a67223a91f04d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5eeb5fbd8f2a24aab91197cbf43c1f09eaaa08dc8d61556fc2384f3c026aff3b62830b5be50ae1aa85e59c11b1996ace3edd2328e211073be5b408397a2b6ef1882ec4b4b95155ee80e009a661a9ae221f23ea5ea3073fde2bc5e43722c3ae7419ed2dca90cd2e604b135bac110769096708b3b8db13e6b470aed84ac91f3e99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ec9daccac3d7abf703d2f32bc4e9d142e2d8e95a3eef52f01f615d0e9cae7667f4c091dcafc4580ae4c5700a636c7fe3d212c783f3a798c419536603df9bcfc319fe634046fe8afd409507a4b1c887cb5e689b0f805d00ed0589936cf8e63458426dd08034673eae7e23cacf1e0331ee0c586f8f002cfc24b0cddac2a377759;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45d5eef1f0e8c6730666410aa03e15241693cfb0107eeace62ba8f278836a0d0967c10c7ccc3f1c96a71a68a5db6434209466308d366191bd9ace53f8fc4ddefc1b5f1646c6772548fb84457bf371a3dcd7463ff5720ab86480ef1aa6cafc63831466110c5240a2f089978e19ab7cd20831d1750db054645bc609d404fed38c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76fbcb0e592bfa4c79d1ddb1496af672472c52e6c6cdd443639a95bfd5dcee87b6821bccc0ebefadafb02403572a943800c85671f69bc721dbf845a8b0c2a72688e280694a1dd5884f51fa23e8a13cf03e3f2f714897be29f8339878e2b75292d0bbde4e6e4a076e063f58d17e29e05ceba80d7f83d577ca1a0280fb27feed9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c15819a2f96afb30d88f95734413fcf9f6d74dc884036ac5aa3a6cfa876c5f0dcf840ba39f75e98161211f2537102330f5419544011f2b71146c4635f53a22806acdc6ff42792a612c259f5a99ae86c1af27630873b08d4fbb06095ee67eae8db83610ca7e78a052945bb4f5cbb4345512d151d64b0f74262dd2edf0f75af69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86ed34c01f51f60a0a8b456f8cf1db1efd58e80b2c046fdf795fc65c092da02789e8e58749f2721f8e5782107fa1a2669a8b4924c546bc7f959154553f6ec18bf29e39c124bbb2330c7a68851238c070f28f2dd07af1c5f8be14089c18c2a5779e82597b3b53a7b2866b5f730746e26522315cae027f883cba24b7876a854bd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25a0a9b0e08cc78bfaa8858ad8f4013838e1a40618f6cc2a79b5474bcee1629e0c2ac7382fa22873067183e3433233de82197ec673953d80fb972843ebf2c56e95736849a91bdc914f3b1ed7e4947c536eb9ce222920307970039bddd25a5465a02b11805dffeef592a770eaef8436edba290854ea48a345c0b291c26d003f8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d16a5456dcbfd7e3c3e145d5e4a305f26116300bec66e6774ca8ef49b5be821762c4373177eebfad22c62eec33de4bce495074327df13b2c1b46440215bf93d24e5fc9bbce20db14a9dccecb2d66a821e65a41e5f020239338a1a6259afe374688074fa8d6def6d58459e2e93de6fb47fa3393c9dc22dcab596fd6c70007a3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a8772a95ae822fcb21250a45f0fb8a8c4797a4cc171cc8b259f78476d00a396562205c0dfce7274a8608c88be784346623a7298bd8a6bb740eefda46764c60de87800dfdb6405bcf2b9bc773a5dc0c8eaab5c54f1cd70817157bb95caa5c1158e7209101895ee7dad8c4ac3cf1138e7fe4848f2e930ff8641ec0dec7fecedb5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9230008ccfa41a1ecd40505e01a6f4eb7de5b93874c73c04da4c9e1e02385057c08cb4a1433c49ca1eb80356fd764c15d031f3ca5ab4e6f275f6d457cf4f17fbfa45098853add296a9df567f529454f2db44a27cbf0716da136b82e1c2fc4b0a785ed82bfbc0e36de5b0d999d5c7f9bc77b1bd1392d61c45dfe67b14b45c769c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce16767a1857b98c1cbce80b2097959c6721eaea445f161643a45d552f6b8f723fbb34e380caae2cb67edff7ecdea1a46f0286af28f8bb2849963295457f16f473adba3e50547261196fa5f3c724748011377f12dac59e51d5b45b07c4ba9b69b4c12dcd3063140ea5a8fa379585826d56f8c6acd6941e6e8350439cc654d0a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb01c8ce74d5650361d0805c043b542710b26c8672929e473d434afbadf2a780ccf921ed5891926f22770c6251dbb7dc2fbfdc02ae6914c604b29aa3c84c749dab085aff9f8d834f228db7b9b995e6084195a8aaa2f3cb18b9223c72deec3ea128e5d61760841eee6e10da10e8ceb9753fc9a58ec7698b1716544cff1ac3f7830;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9701307b86a9c2d73d79fa4e479a6e46bce18f314198d9e494983d4c05ff8824b7b4b7687205e69d0f0a09b1b801014cc63cce5d14a60fe790ff557260f3fb4d4dc284c36e55479c7100b6dbf6581a4f1e1c2d6081d3fe1ac431bc6e83f507da06c44535285fbf2a2df82f7f7d59c79d9567d648886585fd27569778e738e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h816b1a7778073c7978c8d84650231c27a1768f0d53110248887c3bd4cc9d33112971dc91951b5769f8ec7df781775c3a0ce211460864ed95ff4c123d11a68181aa1e5b70b583407fb1d8788b08eadde53eb55004b29c48cce04e11f16baeb6919dde393fa2ba6613c9e35b82223963ed8d0231b599982809ebd3773217428498;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h124cd7a0819cc1c7271472f95547d6e4ac5122360de915c722a4bff4f0662725cb17391458961d71da8709ad478cd28f562cc552211fc164e44249f47dc1fd099ee5f9d2e6da7028536889a5c3419a530fd07d93c83cc4304eb7bd0777dc25eaab4e1e06cdd4968ab81ed4e75920b94473af61f63071b6abd9a1ec11ae7fcc9d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82533fd3245461a89485ba8db78d539f954d89f270b9d5e04c190044bfcda43760a1098dcbc4f36dd5533821c34fc9e7f54c2b1c288871fbe68826e5ea676579743954f645b1c150831025c91b7189cdb6c00abf0da4fc8776f4ed5955710f916c37917630d3a6455b45624bd6369e4b794ade9f6ea4b691a05dbb418f1beeaf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h923ce8d620de379449dd1ababe7df14e5772e3fc1c0eabd183b553a2bae6bc1808f5c3af49890b851088ec4dda73677c4e89227f52c318b8105e0e4f0d5c38203f5d17ec85261604b22873ca35d14731d1a59dbb4dadc7b60041b278cfaf217ce9f8136615ce7dd14edb824cf3123e4f29177350737e2bccb4c669b931b573f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6a06b2095b01d8898e2cb544cb6a093ba41e2c002eaafad163c315d1b21fa76f0f78583f9e9fa508fae23ac0c22cb08ec07063b372a7714acd12c3304fcc21f6e44dfacd92cd6d0351f2138c6a7c769ba980462cd61e6894b13373430245960d4b14bb5e0dfe0fe6fc79096173689d4e8feda9348f8d1b01c6cc9d5d81f41be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a1ab91a34be2b6833191d6a7e4df8ceb593febd4655d94d570a8d13d54fde01f0d6f45019677d5be7853b2244e3e3eaec0b815d51abf0877d7b5d283fa32ea24a9ecfacbbe33bd69b3114b3954ce722aab9bf487372700337ac9e9dc38ade9c2947826b2ee88f301830bf3eda270ae53878ee48dc7009949e22081a5ccf26f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h770c16f90c3d86db9f234b69f9d0c278abef56a6677cf89633d9e76230087da61810010d29e14d016aea99655931ed062c6cd2adab08856fcaacad8c6bf69c381cd4d32ac4b30a0ecdfe0a287c76ebc90a4b17899d8d70dc16788ef25f0f5a201d8af50651b28f01597207d47a674d99dce5ff2eb02561ce8ba23e8b33c8e328;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfccf91d7c40daa7c53c838edfd2418f3a9d70fe6075d5faa0d196da5747092af60ae40f97ee1d97aa18296fa9b16c04475425897bc05c9dfe70dd056358da3c11a89912a48a2b7a1f42e17623a358bc434c2b4af88aef1e5e25f25b783ad41e49073608792daf3ce67c2722ee4ff17627261112ec0d35b4e8a997db71d9bfb54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13acbf0af86fb0761fcb9d886a5d34b97caa69c1b2861e9462da23815727b3d5bab73b85dca55f2728c0db66745dba209403a565d51765d469e15cdfbb56d6a81dad8893f823ce0b13df3ffba62203909d59a06ec1b919dbf31517652941dd5ba3e3c15fe68ad64766e2bad91bfad60178f5605e36b0769d004ca10b62f68c18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42df0616ec1f7c45b8e4260b604532ca7caa771e4cf3d166cadc9d22e8c14a8a8f565d88ffd12b941b031fa970c787b6af3ec49cc38d1805649619a18f427d5ec4eea0b999216381a103ea987ea8a623202d5f95eeb09e40ea0fae0459595a078e5d8bc5ef022904c9df50a4403e42b00a049da3eae838d5422d496710377587;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h280da7d1a8a894f833ded258f6634537ca500d2d3faf12c298fc50383c0a99fd6c6291f21b2cbf30db0a5fa47192e3d33fe1927e5ee5b1a5f279f62df4d708b83b5e2060d18de73925c01db7a3417310e9d7ab4c0ff838c6b64916fc54941ac9b81c2c9167878dc3d1b0c8e842f2318961ddac6f638a74410a7a2604fb1a250e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ff26f819c18a814de825e4d08de4a6106c5ae7ec02651cd0d802022800fa79705258b15febc5b39281ba197566985816c5dfbf2a958b9609eb61b964d72c4423be9ceff945b246ee504992c9fe21bfb89b04d831571ea0bc8f3b8c430f6d21e749e0dde32488cb01715cccbdebfa40b8207912ba8f622697a47461341a95587;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h282d9b37b0abfe7b53ae9da792495e9483a76ebe700e184ef11e06064557905481a3b86532afe341b510113654cd97379b54ec7f2441a88a681c491cfc3f72790a7c2dad5f401dd88e8c12d9ba0f7baa7848490c08641ab677be9309bd6e580aa251bdd2048e82af5d1af7d7d8517f52964d6c10c3e944dd4fbd4881df8487ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ca3ebc3c43ab6066d5dd9de67a408f5305d5a5c3f8085fabe7d5477e782872e39d711432496ecb0e63334f67be861e850900d71d11f153274da7f784e6f928592e0cf66c669e9d77bfb43db98b40a68d20cfc30634dec9038a0edb9837c3c3445310d455dd4cd69eab105ea847c770bb45cba0fa7e5b69bed5391eacf1b8778;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had7c6596867133f7682fd7e7b97d6e3b6b3d0cf837d28db7a104294022a102232ea0e27a10a1ddf7e080f1a2ab36fdd50957e457be22bd6ad00c4d7fb3ce9b4a4d3d0b8f2c60489a7ec485906051e419f1bdf18438a987ec60c2892c39fd8f65e8bacefde32f02f1d77db0a2c98bf95f689636d2a96bbd653b9f00857a0777eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27bfe20fdf8eb9918e561ba9ad136c4e284ea0147fda7dd8588a79e8ea38ea9c02374d9a043842748c7f63a69a29ac923f1a8f22559f296cbd0f68fc94d6d431e39b54268699939a891a159e3eabbd0dccb762920299182a7101004e35ba3fea4ae65ca89e6df21ab41b65707c6e6c44470bf7405ac877cb668b6c15c12e0e2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf16b79ce458e8c14b361d5948c60a56ea297065c0f670a63bb935d355c69a1864d3efb50c9ea1b12eb4411cc2f960aa886764af759416e0a0af9d255dead93c55b553eae572a9cd1f20d63205a10b8409ab4f0a78b586bab2fef9eea6eff3c673a1e4c08df0676b43c0d5f4bf7587ea554a325857d950624a364ecb07fc9122;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc1e8f0996c4c0c82ecce3feb8f88662db1303d977088d377c83d8c14d410dd8f6477bdc779019030dd40618cd3fdf9519a951391f718c120568cc678045b14bda7bd526d47846277f4816bba4b7f6e99bfc1e30cf8d3c3326e7f939a129916570aa8f1e2def250ee1b24fda0d15f6d178b45cff1d1bd269ac6eb9ceb2197f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1f1157159d57715fbc84217e1e791df2c0726c9cfe7e576ae1b6d42f5b1650921648d6a7c46b4d43f8fd01be8aec1412c11975fbffcc69cfe56d0b23b0b969a97b42160b3982fdb3e2b8821b6ae3d050604da566cff83688fb370760d032ae37189a7248dd108768945cabc7375d7913395f29f3d4edeed9864b0e158b69f6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5179ba12c2ff5a3402c3ed89c3bc90c7a1c78f9633ad4826d05e536a94fc058767d7200b546c9e55f4a4194bfe4668f6ffaed7e187e9cddaa5e2830927501a4649af8914239c1e15f7167e6f98abb03ce10ca5a5976ac39de917dffa65449553947a9fbe0e7db9942c350caf74888a674dce866a62438761bddee596aa4124a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17f64533b7808842ab2509ca9d76b6a90fd1e85e98edb2bf4c5a95fa39925746fac8cb2acd57718be4b33c66f5b943d319e546eb314663215c81e24fe111568b8cfff52a9903d163aa13169cbc85c0e8ae5e9413a286531182c29c184b1d7f30fbc8500038be8da3bbbbca31b09d6cdc7b35204d89bdc994599b3a52b5b4b759;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56db4a2dc1f6cfd62983c9e0375038d40e39fefa5fa161e803e5e3bbca8d649439bf359bedba4eac5f6ab83229a16488afb00e2776cf5ae40d22825b4bde2e98c97492e1f6ed5d2e6a92e118b3362d0c68764d066d5db3ea423dea412313c9309c12b2212410455ec7580b7c043a61737a9fe6c6cb7e9b5aa048a9d0dfc56652;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8303196e9244a4881e0f30ce9bc72e445e754f7240aacbe49eb1dcd2662a4c69ae9af462c49e72eed83bc5c024747d6df41b31bdc9487b210763fe12ac50dca25a53094e0507bdd06975eef0445a8c8418dbd149c0d0162abfc81d5d6dc89d7ac093b47889e6f36f1665c3327765bf2a477e585dcd6b22b52366616a7b84809d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde032b1397fc293cd4598f6f52b95399dd1dd63761a993db9a6ec86870e7b11e69a66d5a9eec23dc16a7e225c7cf17be20221f56d17b7e59b60aaad005fc9f3319520e295fc405e8056d39777d8e8d41973fb2aacd4c5d658fad19024e07c0b83da451fb7f4a9401c0ed521533fb45f2c6b5555e892a135998a50e8089c91e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47ddb6f0022bdba5d7b188a83bb8dd39efc31bc864faf261f125b3feb99dc25e872e84c2b294383c0ef7143a1fdf42c8278850c593b09dd4a525827ac2ad61ae2e647af5c30381da11460199f2d95b567c127cabfa12b030e1502102457349fdffa087cf8ca75e17b80162660ef0cf7a6bfe87b221fb06d70a1f8e5bea8cfefa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95501b367d02d5fad3f5fc37dabdc455edeafd1655058085c330c09df82a3e8aab335a4c15cb3c020d61a9610ed6bd12dfa705e7bcd647f70b6a638537a383ba6b26cbed77279cf644d6b2f6eaf9d0d62adaf4e0c0750e95835680d18c2c27b22fc26b60243afeca2de95404e8e89d6a4864d6daddd118e38997ec6002251223;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63c2bb084ff3c798b5e6339d3448009f4aa406259a3bc9e1fa180e4b6773767b0a7f3be971868630bed5620b263c0ff486c3b931d4f3e14833a866d941828ab14c6949abb4f8374e89a61896e34b6e60003c80f8236d2da72f298499173cd1009c59fe596152a1bd07e61d1ceac20e8ee868379a64746feedf7961a55853aed1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0630006ec5a029c7266214e0bd06add683d0a0c98bc10f39fb07e62e69a2857d5ff758828b56456c02c26ce9068cdc5ff6ad50e180a8c3946215b0f01020959900599a6a989805c57fda824058309414318ccf900c018178bf87928f7ec589aa8392ed2d2abd124c05937b115c5b1169c433c0849e1c85a8484feeea112f729;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f8133618a3de319018ef66195d753bb831e4b44982c07da44cc4bba8a6c291aa41379de4bec2a1f906c25dd7c78dde925c0c8180f851e45985f95814a24b4bc1e2c7458349f2c1d7f312cbf82ccf3eaf0ccd844d2f50dad4cc4dc7776117c95d39522b244ed9a7c95bc8e37e3edfc3479692e4b6c8c70f34e9aeed2a880fb9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19f2fac4ebe8f5f7531f011ef3b82aed48d8253300588d82605829a60fa3cf087cb35ce32f4d3e06567e92c69dde51856813b1a6f5ecb65e9d35fe5b228c6758c65049c4bd9b7ddaeec2e23004c49d304935373f2598cea037294cbdedb2793172b8acac8aa804091cc92ea70c71b8b03f67fe8c308af083b1951d3b32d3a673;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3c4a69fb3380ae624b47d06bcc1568ebe51676152d2f7c5fb3874a3ef77b999021862f9aff37f93e00d7ca62def374e221fd10bd92433308b6d95d8f1ceb578a073f2b88651238b2d529067cd215b27a4ce0edc6824603a52603eb9c77837cc50cbdb889accdad14b74516950af8857cc7e1ccb53934ae950afe85201c5ec78;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75fcf8bb456352f0548981420eb5d6e02f532c8c02338b53d03ca91b0a035b9ec1d178b4de16e81227446a8278a9c8ebeb1b8a71101155be1abaf8520d1ea415d3c3f00a68f4f3000dbef566804606110b4facf1bd08361411e59c1adda771b01cc67ab236c284281f38e20caa9f8cb4cf3dbc2fb5f15ae153e8871b4b19ce7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd7b7d46f1280fb2d5cefd698d3bcbaf0a49ab33a9a57f19b84caba0cd33c2ed1b65826e37975e4fda7912fe0abe41b720004ac47ce66254170cc77c3f4e967ff9e90da58fdf471101b1a773facc931f736123d7917c0e2d4a2f54da3423c903e9dfc54e2dcda1049e571c139a41a9bdff653181f713ed91fc757a06831a2b82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd252686ea7f93a2fc4bc12e3479149dc02a719dc918f62eeb1947783a5442d5d12d702c6fd471287edb571ddc5b69928093962891cf7995c0f49eaeca8496312ac9a445f10c57796dc98ad19d4e283ce48e63bf4a170d2c86b8b47fd6e4a8bc1434eb2621366d41ce7f1e38107241261e2539fa75d0b6ebec80201d6f42e8894;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35ccd6e0af314f7f76341a43e87e34b422994d0f0b6f78fe9be1ef4edabecefa0f9a053802a93b71f76f21499d0123e8fecbf60c88fcb12d3e6007ed051614cec51aeb0548f8befbb77caa0f55e68a357dc30d3dae2e377b388d7d544b8a527a25f35cd880e3604768b2d836a019e211a09ac35765c66cade4f4f084e08e65ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29e40a235901a1662c7b523b5798e635db77ef55ec16800a381c33cab0c9164fadb5474cad69769b0c8da219488b14a68319a8aebc634f84ba886803f4d5be59ec944cb3f8e741b29f1dcc8ae40c44ccaaff2fac26ec81de6e068cae47e5f0a756a64e56c19008fc59d3ad2577936f09c83b9f616797a649d9aeae305fd4891a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c89834f5f84cf595c0cb46ad87f6ae4f4c713a959831881439767a45415e4f16c196cf07c9dbb81086285d50872f6405e26066625c74939fb3b988dc9ee1caf95bbfac88995c17d01d9e30046b6b01d9454782ff12129dad6fff09c9724539f0a925af2c375328bcb5030e819ee4a2f517e0980341dee8dcd965dad0747d662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71a7293e140bb1d09da529780e5b55f8dd392172c7b98b3399684ebd72e48d9cc97e56a2317bb1f4982730a8eea56b1d9d4249d1785bb83dd08a64b039d5871f5d9ce283d20cc33f97b5bd194e563a59664434b230f1724dd020241a15b91fc8b9054453cedc39b9ab87fadc34bcd78cf4f8fda8af6dbd101923c36f5cb7e776;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a22fa912948bfe7b3d4f7a4c6384cb2185f4d81f69eccebd54e80b01b7c0a45379c322bfa5bb69dd77bd5aaee3125536ad4cf9e11d762ed7675827e8152b2cf8f9aaec81a90ef16b3b41bc8e47e6d1cb9df7ff068dc9eac58410a75fab30357b741eae73ee81e0b7ec454f660d283c5b6c27ce576bfbaa9e55d27ab05ba36d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had47e31cf0fd960ee2c42c5cfec6e9c1e36d6636499dbe5518f698840900f5859d6047eae1d38e83198327dba0441707016bb5cdb751e3e27db21544387c6e88779d1849c272fbb5824edd73c157423553b17261ec92e060c4dd2e6a14d7f50da6eeb3d64cb08a9066bb6698ca8a013cb692284f8a8c7c8a094cf5d868fc6ea5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he72dbe9e9b02c1eeab90f50f624ca3cd30194914a7342daa32bc623377c372e7751797e96c7f577ad8958592fced1e8efb1640eab0c785871f844e39db6e03e3fbf49557593c22db9d591b5b3f7676283c92e3a684025d4f0287fb5320bccb7c1f3001e16e016c48d62c67b8e4d7341f1adb2a31b4da1a8ab4c8d4053138ad72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha10963683e282c2cfd600a40d519df0950dc65f9e86f24b4cfd208c0eb073eae24e8ee01cb372195d4780765f9ec86059ff0e6f6281cd3310f1eb1589771a5a7ab571e8dd19109b969b40c931173129b2dd3c1ea24c6f8c028b3fffc7014070bf385a11dc36aa6103d4fddb891d5778802e7de76f52cd55f052f632098a3b0b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc39da12af3088a277bca74679e20cfa83d1680664c87352e98e1fadbd7a12ae9658147280787a1bf97ae144fa64fdc823d3135a0a6efd04ad91222e2259b5755aaa392814daf270fada8bd8aeef1b870391c71ac07e0d1a41e5e859e1c55619558b700c11a447fb435444c619bdb4f28bf9c6a30308fd1573296ad5f7e34d369;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0a6affea72f6762ec2e509ead2050c3188aebc3bc8f4914faa1966d88656eb11d8e7335f5a498bd41de8f06b8b0422c06ca78c2b650aaf274c0e95b831940073d6e0fe7d88cce093df2b5f77b2a4c4a78ca1b656b346b1c32e5f1279759c6da3f709dcee841266e87fb41ee32da5393da5f12275fb69629411d8218ede4c4a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26237b2abb217a58422c5bf3c8a9a8ac8b958cb9c4ee688c92645c5c1391b02f0465ae9f969760d9f0940eabcc3b157395b84c6461d248759b4beae5dfc26958cc2311313d427ea6e73c9c24eb0545fc0493f76f3e4b7c24abfb211bea2e5dd85dea439e4bab5cdd1113ee84fa4a2cc4f968fba523b5e2da71812bde61b4d58c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf826772cc8b3e87592b226074ec5f7c621b5fd716b35d08ba26e4f3e1c74383bb374edc5ea039903fc6129506f6d16ef0a90118398328f7f76edfd6df182d6baf1fbdd52b9de9b6d92b471cadc8ec0b59e8eed95fb51996870d921497ddb9a62cdbbd3556281835e2379217ee2ab017b2b5036a30efc844a5dae6d43d5e9c8c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3edf6415d5b7ec7a9c9dbd749902ee918957402ba7b7f4e67b0ad2220d085ee2e21a6f5b46f6c44da686e6796860a089976f1009e4ff27fe9cee80f197f28a00c55ca3d6ac062a639ec94a623808002821a6cf0ac0a294232185bc3973a2228124132745e43a9122d65de9c08d3b751b34c9a261961516b6c1dcbbd7a2cf7016;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd167f191667c8ca4a30ca54ca0dca3c837b45dc4f7e9190cf0eb463417b0c0e59db8f1c0157f1f174f5b55daa1454267ed51fb4ca80174fefb8c935aea24b8930a003111e3735463c0660faf5b4f051f4f1b20ed4e2ed8ead5052747471328669db7becfb63255ebb33b59d9e34d2e35268cba3922b249c5528c293261a3d180;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9974dfa723a2f4bafca365530103711ac391298d4a850a2bd9e1f8722f514974e7e2d9e6a0c3cbd01196b4b8ae2be3285981b99e3b4b9cddebfe14c47e855d731b9a1794ca750ca221957f828e7851802c42306219d8ab35d8e0c4c4ab79d789090ff43fb1ec1803bb75719908fb905e367663fd274603fecacf9a39394c263a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd77735a73a3e9906621ac0af4db038c915fd0e03d2134d5f91346c4ffba55da70ae0373cae194f33d61ef4fad3bc35d7c4a848d27f715a94302cb41700b8b1ddfc0f03488f41768699e3dbcd9d090bc48d60706eef99e1ac8cdc83246abc1b52f71a3094657b19ce0caadba2a4c9de53169cb324db08d0c2d9c8d87afb458940;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3a3aea4a6b1f41cd3f0328a904fe73a7a1312ba3401b1a6e192638a36ae083583ceebe1497d1b5487ae6a3a63795ccbb61e79d3b5ac8c57ac6012a6e95470f258f6966620495482cf03656048bec761bbf4a3bd04ba628c4b0dd37c86a424bafc590130e2f1122e14829f39cb650ea83d9e771f50c4f9116e631df9e1c9a7e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1d7cf3f9ce5c4395a2b0cc0bfa68a00dccda8d6e383b8c7193a35743ebba28db0c8e6fe973a7552d9793d0cf6ae1905b8fe1af41621cd04c4ecb38979ea17595f0acd088f76ebb94a60ce05725fdb633803c594ed78944014460904daee67e53393ddecac516b6be671aa2b3a196e5c1f94b3c82ef9d81bca0162c541defe4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9ec1f88921a2ad3e9a63e660e6bedcaad0ab6808bf27e5142c3a60b13087227eeaaae8b11a19d848c31d296cb2f4d7b8ea3098c3664fb79a16714c7492abd3e2c8fcfde8abcdf6376211bf093d47ccc756636fbed747f1c52d607b69afd062d99cd3888883167546f37dc1376ec28609301a3fc824b8a36ab222c9cf997031f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa1407db93a34dbcd53d2ffd7c698e48a0334cc843f3c8098865aceb5771a4243ee25be4a1631618d93bbcd3f0557589017315c97af0b109c3ffd0f7809e113ff216fdd50cbdb3295a35998a1fc6cf293a29b55ad0eb45ba5b682228f18bc32f6e5b9d7a86251b6d7276ee2986f65ddaecff13e7b74dba91663c266556aae74f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf0be9392b3b6efbf2dc69a86d34bb3b05537fe3801924c6e9d59261225ad9a28d6e9136327bbacaecba54efef5ff2e0a0512b7c9bcd3de3e6d9a85f0e4dce744d1835a2b620a769156fb9c1b619cee44c6502eedd3d965f72e78a687ddb4c110fd93b782e499bfc094506c1f13a8f017b7182dfec8f08595858fc1d7ff0bee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98d772cdfc61e4df6e148aa2c89e641cfad0716f8d38bab1175fe87015314561cd98346b0044be8e581e452098f722a49598b6e126581607dcd1ff7def141c3a49abd8d7dc57e0e53e57855a91c2b74c6e5df9c8e3677a3b84f960ced8eee685b991fd646b7def285543dc5c89b1e523f2266a2de748545cb4f246f836dc77d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h108b4d539a99f63bef8e285ecc9f0698ea386006f8155b1f2aa83c78e7282fc642725c391d7665d4ff9f502a6d47c7637696dcff30de4c1ec80fc296a1cf8de27eb1c9a29151e485492c31728ec96c39359fd94b8c5b8b940791f4c2e15ea31ba0ebc30798712c2b53afff955db087bab9db351e641f6b33b494bf032ed23d4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1315ce12e1611ea19d19102ce387b890d3a3bc70167d356b78252fd438fcdbb25435ac5170f1fe1cd02102312e3766833f891bd6e38ce9221b6bac2d9f0bde4e536e7ae56f840692d90f57c71cb48d2f3a2f9650d2643e3e6bac852f08411bc8f23b2d2352dc798d6c1a24f7aa5893307a7d16450d41b4b189d14af37a2149cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h643f3916f171f798bae0fe15cabe3075683cd0108693346643ecdc0b245067eed4c391edc4092d5a742b58ee335ecc7dffca7f43efcaf49dba1c94f1961a1cf5fa31d143d0a92a10e83f51627c9a8d8936118c066074551d1d311455b35fe09d4c54831a74e3f6476ce7d4536ec649b406dc141fca4f872322457e0295f918cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef485060a90198141f1123e78787175ce1e880e43aee994b5c2f5939ac6577b0a263052ea8570898cdc45e9d7bc987be8e56589c1a394f655ea6b10d64c72fc6cfa0de258123536ef586d97cad07e1780e41086a1f3c0e27700a4cdf6c00440e0bfdf47ecb4687b0b88eac88d3da251bdc5776f68490078cae39b1a3a33dd6eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h219f27cf857315e11600dd90ee435eedfc9665ee05dd49c015ece29b1abe49a0a874793bd77154e6f6eea5286e7c4feb5f89529adc1b2eba5f57a9d214397c38961afb869a00bc18e9571a99099fca1f29aa83a3fce5abb1f24ae0a00e6c6a93c64766a7816ae0fb2900bf8ca8b9acb253aa3906911e4b93d97df1679f77bbb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ec41b82bc0ac4ab750d79d5907b1f170c554fa9c780b748416e4f2aec30c5b25a1e1c10eb9f4648c0a27e4be212cf5d732d0fdd29eeb76446c2228cef60b0db3c0286ed48794208e151c7f4075d48964f2f4b32072b01ff5accb35f50dadafd34de2445677e4205aa621fe64493b4af7e094d5f5931fc3c82e3b4c915f06073;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3090c96530f6c0f479a18f97125a05eb126c502c16be2b05d670f3b610502209df18f7712928a3bfec83704c8df6b0e381b32ca8ce86b665778cbeaf92924ccbd75223f5aec05af28ba35a6e5e1f0eebe278ba503df7804d8256cffcec82ba897a16292b0c46d78d5c8056a94385fa254a412531e7bdc612c09531640d42c46e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1216ff5d6621086e7835438a0c01ab782de4380cd7335fe6c8c3c789d473e52ab6fd2b2e8da94d1beefcbe5bc8dc0a789fe3032de07fc995b48296e30845cdf50b05ac6e329c1af82e46c6c09e65a24d14bb88a419a264cc041c737b7aaec0e26ebd72bdf6bd0bb45d75d20fe0a9db5e891c6a71de6e9f9652e643d2a7e695af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63cefeb996339ffc4860bb4e95170dd4c2e58cc6f1a0c34f80005174747156a6461b8db23cf5ebc57117fe05e8f4f03b78b85094833ab3b6b2ae7c0802ccd49ee14162227fbdca1a2fcc94c83cd96ac9f88ee5445b96d15c215ec579966832109c130f6ef0a9a9ea30f139dc7b315c6036e867c367c256fd8a51b9a4d7e1b547;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hded82c3eb7c380d2b0a29e7a3b688cd339f2ce8edc0ac39f2ac149525bca57b2990ac9ae97552542625e8213dc4c16bd8d2c241d00646e994226ab9e54c9bf70a6fa6be425d7b98e7622349f2f0fbe40200e209cbae5fe8ed9db2e2b6a9255e7ccda13cc34e40845435533117ef8d04fc05c6a8b818cd83cbe8f74e6e7d0ee44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69647a5efce45ee90eb25fb32f0f503faf5cf5ed6d2a50d991f1bace8ee1a2f156a3c6919930e91c40f4282a02832e59835f7aa141765275b767ca28188b1c23402ab3c53ca1c6023ef87cc6eb4368f269658e696b087ee4d7fffc256ac20face8f5ba5376f3738bc9d97ee8ec27c8e5a0018084f08d7025a0417bb360411b7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h405fc7b3e33087331679fb5c8c08f69c5f39fbd92c41a6eab1f51ffa3669c078ef68496699c15a1b13afe4894de1342590f2d9177b2594d6efaa99420744b28e1169d6a11e8f6cf77d3257a6579a5c153d7e5e7f40e929032409f87d2c6e906538acb62fddac2fb9e44fcde7d40e9b510a84ac86a6e8657d4556145ed0f4432e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41f4372c3b9f68cba7ae3fe591a4b20570d039d77ee124ff58b409a95dc666d0e2e4dc87b8aa301998da6ab741c4a549873a1f09d09a8e1288728410eac96b3329f0d98fc1afd50dfdd142837b4c2e3d6002d61d5082088d9452a3268b00a348f62da381d70e8f4f8173f175b16eb71642d370c5673b1dad548548091af663f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e9e5f57307dd848c4c0d8ccd097cc065ea952e6367d2e0b37bdccb8402d9bf8c068c534170c812bef9849513b0370f1ba289b8d3e8ba07028a81f2be31b64f5a05dce044f61d6595b620902ff0b9777d3c9a454275401b03b8393b2ccf33f89f0cc6afa91f557c92e6d7ab0f83c230f0da37f94ac955c01852784fabfefc3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75411878e292e14d9518558d842341fbdaea224d434eb35782240197238174ae8ad78bf2f5e288689ecb452bfff999ffba1765a0b7ffed6cd2978fd540287c5f0e1b43cfea44b8ef5d4305f068ed3da301a2a72536e63c853591160104f62a35e17c67abcdbbc7b6a8d6979256a615d558e0c66aa818730c56ed1fdd79724b8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b9c7981a9a174bd78619b71448b41fa3196634c433331228acc91d8028cb4799b0c962d8dd1f1805af5fc4b8b834aeb436e6c916b91364d588c4f4acfbe6de5fb2995ca5daa5f7c624e82703a42786eb5571f4a303776ada9f413dcbdddfc858e09b6645afeea5da8ecb763a0e5e426dd35a3b401449274e0d42c239464b0f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h470e18d2351b4f7421ba1a891c03da1699f21ca4632a0b3d63c7e89e20ea2a8d1edad424967ec1b45aa126c114158a6eb94e3c6e670ab8a561400045a14ede56d13744488426b4bbda287f9b4639b35f0d8b01cde433f1eb7b58cfc9328854bd3ba420a0fc2f4b74ad38a6bfede044608adc212c428090737f9828d23d346a52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33c9c6db5094825cfb5d4ae4a57e60ce5b425a87ee494c7384bd6d6853252cdfe90a6bf5a83746e223ff995920e558a0620733adaefddc52a4344342088dd58b62fe46d3a08a4006fc57c96e3195eb44080ec79c8d2a12318e92a3b7cfefdc2dfa0653de00a09a8d2be72c79867c2b50cf348f9cee159f7417a6164259b582d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb12fce4bd9db5c027916693dc6ac344c7108538f5fa7e14ebeab7648576621980aeab1384ffb60b01b8a928d257595507f9bf388f509e42e49e4ead6e63be63b835692633ac713fea99d6cd22110f7cfbf15aa360df31b013584ae6db7fe1f30cfadb2f1787f2f2bab3fc61c7ce57ff8bad9672ba09db1a7d2d776bb27375631;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h978ff50cd827da8486b0119a0b4dbd62dd63176c05b4631e20244d7683e711b614e1fc70200e1b3f30947bdac9209beef2be82e38c2a0aab495266663b980e7bde9fffe62226042f8e8033190da2c6a29b5f72f44fec1c27637746e90c48a856dcd2602974fc3cff7b35904c50a0e5c56898a0250d5fe16efcc2cdd759847809;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb08533d21741b916936b516ffe31d48aaf3d9c652a95047db8d11fa41772d440bdda2cb296db840798da4c7d12684a72d57edd2339efd3d6beb797d9c7f8a37260dcbf33f913eda5e8b8bdc6782440aae9dc5437bdc685aff400aa1fad867af3b4a214615c565f24e1421f2248ed13be9382b6787a50565f5827538cfcbae98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d2bfa213c28e6954524423b5a31ca9e5fba66a9a3660606725779624742d376de522b73912dcef92dbb8fc6e52fa9dcd49850c4a13826a70213fcf7dccdea0f2373225316f286ee640df504fcf6a9e0347e62d907320eaf1fe31ef3073f728827e38e0e7fa88e54f9e00197247bb774b41285a8513ef626352709daeb3f1baf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3cadccfae139a8c1a11560830a2901356efb1e6fd5309d3675fc494156fed0960804c0875ebd8efb1f83d2a9e7455a2ee595f5dfa97ac6fcc2514d7ff96c755f8e4176e9f212315171ca80876f70075f9aa91936a905cb60ad4fbb0e5053aa6d89784a499fc6cd0577ed46b7b759f84dde10b9f2ea74cfff29d272dd3be647f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc57f546e45c77a8957a8546a84768b5fe035c1b2a4aecb056c5fb641573bfb4be877cefa8fbbaa08c00b2f404b403c3cbbe19addeb78fd0eff5c7e5b0b3f8c9141b05a9e0035fd9a89f72624dd0bedfeca63b154835da99b4b6babb2b870644d5478c03d7eaf964a79397ccffe61eb7548ea27be413d8fac3d9c41e728eda496;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h198eb0c043ad74846658ccadf9b019708c23b9b6ef8564318bb5dc5522cad5b6bc8752379d0b520ac02eac6d9434eb353969a19f58d70b744b4055837842ad0cf4df062080bf36fec9da1b40d099d63e392ea0803343c9aad0cfca741e68f150ad1ab4ff203fd7764be91a8b46062352d89b1009bead395752f033ad605d666a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8931603e899c2bdadeed0930a386e74aafeb6a1e622d66ac0ab48b58520604e3d79b467bd220af45cb8c734cf4258a8efc791cda04af852e2dc5efea7f169e252dd2667290a63841bf6d0a4a528095fe01cc12e44e0dec2ab5fa026fed9cf908eb103071208fe753c85e17c38cc5891ef8430db4c817073c7ebb34abec749cfb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2b38f6654e8f8c772f523bad9458d59909bdc06b6fa3e832af3cce9d2abc819ce1e517802d800c87f4255708e2d871b70f02d0f589ca94c03deb0f024ad0251ce465e85a16fcd6e4b7c31e6a74f87fe86083ee36860f69e2bd360c66b8a49b319708eaa3346fbf7f1fe74fa08a256edd253c57af238e77acf3d413b77208836;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfde9f869850caf5af98ed61dc6548559afcf49397d254d018c3101d15048d1eec38654763b7f076707892fd71321a6ce003d52b24be8c97ee3b275f41e425bfb14ce5d4ca9e97351b31ec0a2b3065b1c9c3c405c6cefa18fbc16b8f3ea3e11075ebafc0ddb433b09a5eaa577b0d97fb03296cae04154bff11c8659c26c269eb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85f13005719a838d0a58dbc875b203a24293eb8109588d4b87858c66f2f31a68bd7af1ff74679e90652b0ff0d57a197b431fe3e424077f545565f412ec4b05427c8233693512e0caa1d7cb4e84aa7011d9d20df3299bfeece11bb73f2e9c1b468496be7de8700cd08d1e9bac140b027ab55f4fa2f0b9b189be385c55576fe9c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dfd76c898b7d19b66067e6658c9692d757331493dc12a9134830765990610acc6fb631e81344f2b249bc51dcd4e74a74abd52531e9621030da27ee9f59f2e97e14443852009d389149048f3932af7a31a68e2c9bf56ea7d4120c8116452f77b2f366630078224a18460286f6d37ec8f2ce6cc7242705ff7751070fca62f05fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ae93e63d3c4d9bd64e7f8ad0ad5c2b4f81b72433d4e74fe5396b882b74b0cdc63107fcb5b049b7331cc9b86039b6ee19bb8effc76b747fd98f10f9bf428dca473ac70f05226a8a1c78a1250e71aa408a1d890b8fa181368c9ba069688cbf86ecf919b49c5d0ba8f22afbede625d155cffba1ecd1c66c1c3d18dcabf10dcc4fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7794c964bb055fa12f9843d696b97af3f341f8058c4f7127f48f92c87fa31cd56a25c6f7c9f9c81f6f2872b1b8f84b79b3d51d0fff6030bef626e1928f3f3a7f0e8684a3baf5c34e7d3e338ee94bf1ef11871883229f590d59c54e4b3b27fee7d0fd15fcd398bf44af8e371f47df5778f67886c9d19e3d8fca0662160e7f9ce9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94d9d87a2cee7629ee769791be6c8fc0dd4d3c5e9e142487c98a93a2a342353a6c18b72ba9cc3f795920345dd13555590847f2815c8af9b73b9103f60b42fa94f741efbac72b04146ce450fb41644820087e61c5cd6d3199df4864a495ecf7347459ee9d5d4b1e559c5880877cebbbf169b96251f70ed1a7c4f29df7c05ba885;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cc90cdcfcf16b3d0ce303f164e5e4bb2a8be7511fe81c213ed5ff62493df452243652f25bf7f061402b16be856489cafd6e2c71695e18d74f8e6c064583b5d6f621cac733e45dcec839ae02035930e1be742a0925edabd19fb97ae09b223eb1c6564ce27d54514c53b4961adf80b5a26b47a5948bcf93b480e1283593080b00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0ebbd2bf8ff4466b01fdd4fd92aa04eca35f37934d19cfdbd2984660dbf35178e70f42b78f0c23cead226d444836c5bee295d4fbd15483eb017a1978bbb047e56b9e4a0bc9d94f5731968563341bf514e69db5b9656b597cab39653df564db603aa5e96a86622383658087ecb4b39b33ccdfb96230442d65ebb39e142030add;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19177803c832c69fb20aeb3bf7d721d2ed3203eaa9ba7dfab209c2baa1451f0b4ee481370213fd05c1ebf3d63183a6c1cabf8f54cae336ac717727ac5299e9828106f7effb0821d4a0e44df150ab4b0322752c4010ba11e10ddfb6c890cab50ee24a91a7590b84e6286dbb14015cb8a7181e0491bda8e6fb4246fc2d0a6788de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fa31a284b2d57f8e6ff856fc84b810516b9892b870a34e709f9e0eec0c8baf3c68a631c8ffdb157b652bcf4a2bbd13051a3b956494d52bf12ebfe2af846f85d5f233eb98f80b914c2662a92d932cc4aa6ac1c87b3a011e34fadc2dae82bd23a5f2a8766b358fd796b0efb5db6e22d85be94091bc7f15d192a9944eea71f4a50;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32174f87644177b2a9ad3c9f6124be88e10f1c3708628d43852ed07720ff5fdf71458b6b41abe4f97233bc4a983df3fee7ddd818041ac3293c93e584cb46b227384736cdde03e247a7a57b7235cf9feb0b5bd049f70ac27fa92b347466e6ea43c8b252fb684dade6d44a726146c8993c105fe34c2b5e5d1241ac92642bde755b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h816195c1aa7b5f22e9512f6ebfa4c4c15d8da9f935c3308b618ee889eaef3d2d09916656db65f47910fdc7010b4b5b208c1d76f113b99c321dbe47ff01c13dce1b131223a346bbfb0f78004d86137f14fb0a286857d461d280c7f3008d0842b54e30c9646f2eba69ef95d242b0179e72b9a9864ddada2be21a4c3aaa0baac71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h970e1ecb01508472cffff407b7c1bb662df84c3caaf2a54f644519746caf919f3f0286944c33883401844761787a5bec1cb24316903fb4510d6a9e4eb468604f06b13a03daa34490d21d7adc98bb8dd0831c935e5f9e958b925c4bce34c4cec5a975249fddb1c9d59019f3d56a670f6ce7397e5193ad7ac0b9660214291baf20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85d0ffa29fde28cf4f73c8301c93a4fd2f9b15283f44268ef0112da08097155f13727aae21e593466c994d19e33a903f0dce987d6298d7b3d265ddafcb5507057964d9b94170988f5f01affd5843f333fbb3452d1a62dc021c8ba699664e0f8cc84bea37edf4dcbc05b1212a2f138a29c76bfeeb9fee6ed857bf3f3acaefd33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf11d77b199d8b60ccd8b312937b1e555a633f9e501617cc6096e06d1438f18ff09b6d8d8b224a64dcce042b2a1ef923cd941a4510b82e2b9b78ef9cd16c8332d9cef7f9c2a634f85855b668dd513e2910c1f25d5e3caa57e80ef8df870ae8d3faeaa87057a2b36ff3f9532d44643fbc10f039c995927324fd92b30f8f9acbb43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28017998417f52d086f2c52cc46926742241bc6f660ed0d140055e5424b01b7332f2e2da791e48999ed211139d6a501feea666bc738fc785cd1d2a77c33374d991662d4e4c7e29d1e5cac23b720e5e7aadfe06cdd4cb6a2600702c0d0d4ac78efb63cadfe8bbec8dd56ae11b8a47fc69e9004fa2e513f354c64e89c8ec235fc3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35d0af9eb45392a04ca04f473b1142ca0600b20165a00352b8c569170516a2f4aa3f8596a4f30c8fb9ce121b85a32a738acd5d70c15a6cdcc4d73baca913c08aeba93cb7b895ef3c486575cc1643199daa012d0950dc14715ff34a688cea4134f4187c1eb96c4a02c5ffa6f233a9ad8251d12ee97d18e1364b0a7348a1e39388;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h244636c004753751cf7476bcae11680fa75a71f90271d1dfefeedf89a2190f8eeafc9f10108c0a2753ade1e4d8f5a9869e099a44e91b75c6c9d108dfd51c90d8b8bee21003d07aa486b048c73602e5b9682d2c6be378d6f4bce11a7301fd8c575f8a35ac3d1a170fc3f2cc17e0b7b462c00ef6c5cce93aceb2685af43806e350;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ae3e1c8b22fc67a9f052af5154f60f8df9f79725bd4637193ca01cf6f9e94e6c1bd4363598c774cd0d33f5c374f080fc4ff30f540734c5307d79668667b9fb1c657f920dbfeacfab5d54f123e11598b0e909b0c8c67200ae79aa1561921824c30e9e4cdffdce0e9b9a52b833d77cbbdc6136c6032bc3ea9090b8d64e82e8ce9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1e249346d0fd1cd29adb1b683b7aa69cf137448519e83a454736f393e962423761b95386e14208eaa1e4a2d46cd890d8261c52372d613e2b18b66a9c62157b5c4140d0f886182aba8193d2e4934c0ac522d99a39ad74c7ac28624cf899999595ca0b596b3a74f4f698747a28061e319f65f2022d8613e79339952d5fff8916f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36a469c40e929c8dc004d0fb18094692b4fbaa31e55a85669e9d2b56975c12872fad472e67b5a42600a4fd2be5e01a637fa95a9469bb96fefe4532a40b06704628a5f854208c4a81e248d4e34d6bca8554d44935b3911fe481dfec767a3843196aef9b47968c86dc7a0a21c17b542412163a394748f5b2977c3e1499a9dfd15c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2f88c521eef8e0a4e9dc8b62a2305f44114b026b943928e03b3f094e8518c570afdaca59505027e9550572a750690ef479a542954c11334087a019e781048460854aa296be8fa427abcab546912e3fb41041b7ecc290f33234043b59559abe77031df89cb4ccf69d3271bc18fb6ba3aa22135f53f2e2dadf295edcb6a1c0c7f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24df6837532431d7574d63ca45a11fc50a44e5432f2f6e382011d7bae81e3d3498110bc7ffc2ea90a347db0bfe8701fe85aeaf419e994b79a1e660fe5e546596a698f150a1d93507cd5f0e889b30e179da78d6d08c90ac7617be5518289d9e61ea1b9d6b13406899d39224fc4dcb8a4d0c8782f7a757f0e0fdc982917a878ab1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h793385aeb367087a2306acc47013e7180d024bce458afeea0af392d636cfe3cdab54050c0038d0fe5288e73ff1b1cf36cf60907b80ac33994435696fda799ce632f74e9c3dfa041a7b65ce9c2679a4e66dbc7ccef6e7365d667b39398d1c5469635a345f3cb9638d5595c33fa589ca8481764726ed96cb3a8b1a799238adf498;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd431ac560347ea0d71633125851b1a6953b3ac33ce6c4a1c2806f5479f39a55e4ef66d14a9c027f4ff678ef45480f6c48c44908fac9d833dea6c9e5dfe40a1c7f54b0b2d5eb37fa1e855f20cc9956acb1b201bb5b61da81a159ec534b3f4e012595e8eda658ffa71a5e76be92896e2b6df5a660b98b50e75bd72714e0241bfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18007aade8a9103d5389b773dffd0a16229c2cb70aa2455c0303e5a128fe46c950a3dd2615fcfecc8488b2c30237eaec6ce52b572f7cc83b5bb7c96d7a7f29528fe9967d0fa038892ec501e29dda8f6151c03094fcb5a8add8847587adae11acd8b45789a3f0498728ca7bc505003b7e79c6952d5d1e2dd71f084d46cc788adc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce5f61a17b2dd8d4ca8113bbff8d238ee5653020229afe51f8a98a121db127e2ae0393370c199ca8ff8bdfc955e1af318794d09833dcdee2195958828046be9dfbd4ec39e5c5ad9452c3ad53e81c5ff4faaf51774edddc4055250ff65f9ac012fcb86533f7659e4e8916098a78139781f051a710ad84bd4d98daebb62a9f34a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdeab2a80d46993b493c743a1c8ffdb78bbc64cccca980b649ba47aceaa216c3fbacae1a197be7616cc1cd70307ff5652834fb167fa46fd0220de2d2bce74aebef69bc9fca9ee0b3af22c57528d2709a3f0e4d88111152fedeb972e11cf3e0e1906a4af4e62afab674c713d7c9ee3b5628999c349744ff746ab753c416b21a7a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha21b311c237cd8304b9f5d8f0eaade272e0ba1a120c8bd688b9e8912e65dcb7cd8ca2458c3ee184152118d9407944af3a3a7477d2311a12a0e92f88e6174485576aaf719c4ef572af3b55d15477261a20a0eafcb2455c9176385a5f425e2260d613eeb18dc31e554a2506273878abd93cc2d784e9c7bc22c68e455b4fc7e190c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55ddadf831d61978f39b191748fa441ab98196a049ec55546aa0e01288c7e063e3fa33dcf53c4de991fcdd23f44aaf9e2afa9c6491046492f088064e18ac7dada1f66ec7e7b9c35391d7653d663748c25b3c439a8c594ea20566c3939db0ef2978b5cbdfdcffdc4395aa37e08ef7296387a77e62e37895118c74ddd1bfc57268;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he818c9e6430f5d9f5a80cd87bdf021c4a96fe94e339a8d9c091efca33a48b6d4124ac4e8e19353be70530f422c14d7539db08a1429b902fbccab3c664e53317403ce6e78df0d161811741fd20406a4a18a73c7f1025ffd4e3eb9fb46d145a794589cdc9fe2d5ca9d1345032cefc2b8649d463448b50b67b894a66428e122a631;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he513e935b0d0762304e3b158027850b31a196acb1bd3b2d472afa09acf108420f4d948f2217bc5571386f487eacf9fcdfd99c6be2574b80580d5ef3be7106817c36514ef00f71566a14eeecc3d8a962ac2ef75878f0d495ac7ff396e9f5f1731b1e3ba0ab631230e46d0da330bc1d4ea4aaca21cc79dd19c6d2a73381addda52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35e63825c4a818a36be14a3243aec2b2ae1458143136f89922e716f6a5862a7bc70bc2d4d67345c6bf300db5208a67e619fbc6189622027a74018b167453d8f7b4aff2dbc9ffc62fd4ee42c5f06871f24ec99339ba91041bcd2d04601aa8ebcfb634b4ca333569c3570b986b14c738666d921841ef5582c3c7da5e0261249e9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c99e5a23ea8e49ffeb32f0ccd114a6f6254904979005f1df90b710d0e53b27035e0cf49070d18ed2a2b3287ce3113860468be68ac35cb1cf729b0aae48e9d9566e0319a4f9165fe3a61254c9c6db7d084b451237f00ff21b273598392740b97eedb4b3bdf3239307974bda712382d1eda038f5a09068839452f76025ca1880a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73b17d1fe95741350086694ad59e2871cdb6e334bfd3de4c7fd02a5888ecb5ebd288c455e86840ba4c78171e78611e750f81d20f0d9a5b5dcd9bf6382a9b0b99709278d0ce765a376ff9cbcd37508e996b0982c4ffc4802a638118f558443220e9dc09015586fc757eb1472f1cc6bd1fce0af478fff8fdbd60d375dfb164456;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f1dcd11af6a3ae6ca02f82795e0e76515cc9ac5ccd109583c7f5f1086e6e3182b222d108240f71b6f462cb6d2e8c509de91af8e50e304d4dc776fc26bb3473962773ee62b3de18715fbe58ee9d9c1fa78358b1bad1109c1cf28740e8d0f8301dd6da710b34d636f6b4e15807d162d0a9d5836848755d66454e4d65cd5b9695;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b6486878b7d49699cdd58ccb6153ae659a9b1d0302f2b92bf68357a49dac14fdf9955502154b431a05bd8e2db15ebcbed9fbd46d518cf93ad82eddd09c3b0c1b763987a38fab33fcc5e3993ac65ca77b7a49b9d4562146a9aab8a7ca826786a507ba5e7a820e62e89805259da1b4cbe76ec6e6057ec676d6adf2f4b9aa922d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1be5ce97c05f84d7c174103feba5bc2bcf42e4d37dab8628fa29fbc80f721731f25e590ea65556f22f514a229581e8c865369a15e0d37977c77c02167333be78415f84cfb8951125bb583700d752efd8a585b8db6b358b6de74d2a8d19edef112418a2ffc94c6665f8999417e60b0d0dcbd0272887810893cd0c0e986297e024;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2bb0913736170e5b18be45716ba3113433084fddf0861d40e8504d51528dafcdb546369fcb64885a6422101de3409efb344bc279edf86dddf8ec3c2c5f14cef4ca91f604b168efcea4393b2f7668d63fb8e30caf802d9a544820f4421c814672ceff6f784cb83a36d9578440e42d11651341892a011dbea6d9a70eb7698795;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd462268dba0c0cb09c23c0e0ecd1957366b6190cbfc61a2f33ad29fc61f0be9c1b0b8a20e2b086faf30015fe70e2ddb6612508bcc3d1ef3f3cce1be64d0824387ef19b8d905f0c113bed240991ac724df87f87d72229c7eff8796859d30539e9676a5ece43d8f47d9f44b43f46dac983c4310c34c9e7e6791093fceb8efff0f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4098807a25883a2a223901173d43f608cf9ab45ef5abd76c4c3d42711a98e7d458a36bd1c94f07b921cc8a85f18fb0b6203c6cb7094041af39f8819079196cff4a0e2664b49102cf107cc662039090a81cca9cc19aeb2c2fba63e7c1d34f54455505b9e4d7e024441061e918aec59595032ff24ab8da7bc3016137014805faf3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h983ce47859f7576f36547ff124dbf9e4b8403bf96e2dc48d4a1dfc5df7de4c6ec0980b453d1cdc52453f85d03e723b91b2690412ad3590b08098487eae358e63fb9fc252a72d5c2183acc25dd70ecb3401489b173dc91525e1bc0454e417ef2789813979aca1b41b3d3e4df4ce168f8d4991faad8484dda9d92360f59410742d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7e761b85ebddd06df70281c8fc642f8b87a553323519a16dbe95469222bdf44e07c85ed928fb4b5d699e0a1192a19190c67b977585d722bba5fd1c08c58628c6ba73012fd4b62211d844d6c864e01aabc219790c9b96005633a68eababd46e2b5654778fddcc2ed6ad843ae441f845d98b503da6875681bf33561e5a0201ec9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83fd4f572a9ba443771d65e6527e6aeadf79d13a64653f631132302e3748f42f7b35e5b4668320e6686ef6e2fe3fc25dcfab7aa6daf49cd0fd74590157f0797bdb06bec316cbdeb62ea286f33c60d9ea8f9f7de20e117217c6e2e95ae83148e2d4990d2960d452e372138ed4382c93129699d5775730c1c67869965e90158135;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4fbf0b995c6a87865cc231c5d81928dfb8101654f466e63c81a29e1f072355e12e2f6cb884f1fd417f0dfad2d9d54bc987edb61c7ac4c4e7b764337205d3ed4ab4619f2ce1bf9e267b1b50af58a9cea0a11aec1ffc412e918076a158cc8383d51f9b16681ef82c2172f2a0f5a64ea82a50740ddac870a8f2dba80ab1671b5d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd050cdbc590c6818d253977182c0cb40a99b4b4ce0d277004abc4c30bfa2ea7a588f0fd9cc5526416fd83b62e7742a2c652a70b6a4aea6b7f7577f7268cfaef3f39124d8af2a3617dc85c401ea14cc4d3674d0e28264635d739675b078445c0e57ca83bac72757485c7cda3cfcf639fa9303f3d2ba7500e54d9feace8c06a44f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h628d8c6dd1582e8e2a558e118da91ed2c6691f7bf81b8d9cc22e03c9f57a06b2ee47b29072bf2cd6aeb759792a13b5507d69d041d3918d1e561314503ea4d4a876b4ad4087ffdde432236a5db62ed37b258a098917f461ed737d9c325935467661e7e2d2b112663b2b3a621bbb81189287ad4d7674e06b067feeabfc0a552951;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8de4a87161cd6a7a700bdfc6c08d976c5b994768d4a4f9378b4cede65e35b2d19643b908b02baf85620b9cffad1b0041bc783a1a147a275b69a2ddf378d8e2c6a8c1441eea6cde4a8b7104f27d4c34169c30d5e8b6b5bf2a9ae7ca9524ba07119ca1d0bc6bec7851c1d95e1040f84aff02b05af40c4bad0dcafae478dede3b08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57e7a2b9a195940706dd4881ff132bc9ef4fca4e3e63a9c35602b8db905f6b00081096a6bdd6cd328a0daff3925fbeb08c21dcc699f9a2c4a834f57606b37716017dae7080b4a169dc5f65456e1239319b2b40c7af2ad7f1d7998c49aa7c970ed04817cd288e2c35543c0d78d1400380b69a7fae18fe3aa9c1effeadf0e0c256;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48000ebb98f9471bab7b9f8241621f687b831f937870bf309a34684f9058386322a15fd3732630f6b496dcfc673c05cd2ba35d6c6a5303a20f23daf998286f3715122f60b867a7cc71a93d8aa774cef7d6e21f6bf0e879aa3144916a269b4ed8b3a0593e107bc4a4bfefed912fb98f2d4d0df1d744d525fb720632b4c94fc2ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4b3e86d888f83426531658432b6c6da60eda952234e004ca88a68a56ad411d6e076d2402b0be973800cd6a679fbd98e5112e338ecc6c90ce486d27cd2496db74e5a3b846150b8236feff8574315149c2cc2e3f2bdb06ddda51d95236c30041151493b3dce551f379ba58b749b588fd1ec3139028bcf66fe2053beb817695c2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b65cd5854f93ec0e138167ea433215a476e113569f104ba08b77b3b4881ce1d23c6ac93e4cbc685512e06dc7981125e3e6682633fa02632eab8bc449ceca4bf97eebbacf1eabeb9025ca1669a542e000c82dc343a04f7aadf6b030e7a0a1d3fb946a58d06b218a2d56b17c1807f77943def29dd084093340f457b2a2d883ad2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bba39be1ba7525dfec863a73ce71a8a1f47cdaf5856db4e44b2a11695c061973432d4d184be09a819f5d4948107f90f598c5ae35e7f307f2bcaadfb9e41119dce56d2266191da191da16d22f0cb0b915d5489c22b9729c9d10c5d4a0c4db2f6051a70c719fdf6b582866cd821252f85161758c7c5f0995829993c353fee69a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3db2c580da3017338bd9a25dfd6e857d5d1bb973a39c016f364824460cc201b6c90b8d9b8a955e69870703453c8feb96d1600e326e8c074d4d7e94cab9f5ea0b1bee5e587756c727edd11988451f2f99962001acb1f298eae7f775d23698cb63977511cc32969435a0d75048de3c686668059dd73e92eebffb8b66ba24466965;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf6869ce1dad58655a55ae49b6099a08fb9a4cc13d14f7727ee7eb3ec2f5022e1c9f9a7c7a92606c7e730bf2148b3bcbea23cc4d27f912526436ea47c023be2200bbc47192e8723830b957ea7e1e0ccb0d2264c17a9d3121db61c485677996612d8b2038b48c91992156a718c40445eae192fcd3f29a53042e1b9763fe867218;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e6d9aa1dc8c8e3375c9c5252e71682f773ab3df82d4db92b112d3989a5409b88c28413a4db8772901a79369038be3711a14374b0223e7ffa57ddcbc829ffb1640b2f598c231a3d668f0a61dea0bf5f9677bfeb61f33bb239a8065891d8d005355879ceb082dfb225f5a579c6323ba4a3875711fdea1fdf2cfdfdd53c4c81488;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c460dc7f480d8d03e55f9ba1617603416c34932d13fec3cfa12e10ab5f2be9c7b1a15e30e2b9a5cedcec31fc97aba422c5bea8d00073095696f84ed3aae2cf1d7a69b2c48d29935947620cbb33df1a3fb9dd1e1b5c386c8a6df67b5e196d57dc8b10a5a7ae0b51fb7607f4f36a2b71bd209fc9b765e0ccca84fee6a1ebcdfa0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a4259624f975e75a0607fe97d2f5e3a00f57a65ec22801d89f13fec051d155fa794d77167f4d9b83c464e7a740b906d1e167317e089bac9aeb2d3de95a9846a284cfc60a2ce39b8529d631b1be78c638907675d65e09d29e845027bd21a515a438fadb6f9d125e1f56d29e35cd76be79308faa0b0918a084957f7f3c8acc1c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd28d52fabff959b32a18b736e0ff2072383203f2c3a288796efba4e9860dc6ec7d515a1a2518ac19046df8003751f88c893c8a1b43e2494a359c86ada1995bc239c914f6c1e9b7e744e1969273312701e50d99c65717d83c0205cce16b5a6e0d9679a3bc95e6e5145e2c72fd8804c270ac3baf1a5db3ff59ec3b83147aa9bedf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeecd267b66b99ddac4005350fbe8aa762e1f41b12a8d9b98b34d287ee46864ba3b5fa7b7acfdd0f2368506c7746525c3e855c85215fe77f15411b084c108deb4057df6f9b460780ca6f2390123acecb73164930ba9868f40a2a138e5ae8f17a7dce9bfbdcd5ae4105b95e27239f4d36aec38ec2aae60ea6c97a777f8b791953;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h589d26b7ead40894bac96d19115de2e92e824b9fdabfc0a71f6418edd4982e98656e3d1e5df228e233edf118a785ad0351dda8ca1521dc7d3c71b881ec3982880c086cfecfa7eda0861bac4d0c8463ef74f49866e1a9a2c9cb125ff21c91c652171eadce3ab0f7c949c71c2d9ea6d039ff6f96cba76a94f651297726fe3eead4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd167d8b74607173b2a74867f69b51b74ead2ae7a9a77b40be25d04f7de3cdfae83c99510046709121220a75380f49a04470f792739a948ef829d661a373442db7e21c92866d48e088a99d946b42eba3919a3418fd78fca8c424433a19e4eb75c931eb1b02b36159997c392ab056b9434c94da13ad9c83467b9d8e7b1957f0ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he078c8da5daef2f75b1e8cdbefd935e42e918a070cf49a87b3a02f6a7e051a8726ce317215af2ae8b273a1ae9734bf6db3131c6e767a0d6ef5b3efa4fb7f3d21fcabb80f20361116cf98805619eba85500cc82e3a5621deef52603ee2901fe04935cc22d8d7a1c4bb93bdb410f7009f1fbb37f59c5e504b2fcf3b1584614bc7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5861894d3d91f99a1b7560f207a20fe083dd256ca01e0303354b5b4a578b853927a2495e18c9bdff260b540de3a8cd785c37904b9f64cce9573702adf2603b83d7493cd9ce30b12822c96bf16ab0e2a3bb7a0665df71f3bf64a43a72cf9ec2d3922d1aaa64fa5f3f55623eb337d112917d385a8489a107c61746c57092411e67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54d0e13e6a2c33b5f44aef8f7996432e4aba2e9ce6b96ff36c664047a5b5a3c759e2d5478de24096031749e75513980d3870f1eec3db1e257fee48844c71db46e0619a23240f9894831a8be8a2ce4881f0f7aba44e61b043e4560ca3ff462bee8a8bb7c172180b178a5eb18815c2dd48993287827460a7eb0a763e1ecafdaa26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca5c23b83d088a3dcf04e067e1dbb83ed9b55ca9f5726a79640d41ea2a5008891736f91b6d4a1ba06418c80a6f6a81988d853a52fbad410ffd4d7b90da77234337f00150f8c287c778cadf7c7f1f69ea94c516fddb71546639d66d29bccc86e6feb35c567a4d2b26acb19571cc1f541485a5ec5a81a3334082f3cc661224b36a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h862b5cdd06fcc04eb7f21ba6808f497fd6285753e7511189500282bebe0209c2dcb2c5c79f627f784ba61b8536aba3333ec60a68dfadcec2510010f2ba25012076ff913bb9196584eaca9f0260316f23cae07f0eec42bf26984d36bad20801d0285ef63a00a72661f5f99f4480c31bec084d40acf24e975263d1081798ae088e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23016825d11493958cfb9a92e478f283bcc84fc903eed3703996fbed5e6555320ce068b794ad465a449d2ced8bc2bf7fe2338c10a83b5aa02212db6d18ae4966c2c891909015ff0c2454ad354ee64f671dbe4ba41109670a6af341bc45abb949286687ac02cd3ca08a32bbe182aa8af4c04af2245d3df6a36415b2071d11de74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d021d478c691bc9f197d65f89d13fa1f6884598ab49c124e0d14858421a447c0bde97e9bd1f41d073377812653f1de9c227a9fcf3310e40f3f42daac3e502c700003472aad7ddd3c5d6d3fa6c8d43f97523f88a41b0e9bebce687805674412b46e161afe2aded18c136814e0d7985c68dfb1df7efd7e4ee70d42976d1d8b3ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d81ac9609b9f9b149554ee8b3e77777bab2e92432cc622f3ca0379577395c6bb397b8b0cf406ebcf3ef0cb70632fcb5bd36ca19a6a8a5869e5c22092172f498e3dec156c2b0f0dc2be3d5175aa380883a2db91a86fdfca06d2d3240ada1092786f365cade696289d84a1ccca7b883db86cc200dea009e8f166f642274648ca2;
        #1
        $finish();
    end
endmodule
