module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [19:0] src21;
    reg [18:0] src22;
    reg [17:0] src23;
    reg [16:0] src24;
    reg [15:0] src25;
    reg [14:0] src26;
    reg [13:0] src27;
    reg [12:0] src28;
    reg [11:0] src29;
    reg [10:0] src30;
    reg [9:0] src31;
    reg [8:0] src32;
    reg [7:0] src33;
    reg [6:0] src34;
    reg [5:0] src35;
    reg [4:0] src36;
    reg [3:0] src37;
    reg [2:0] src38;
    reg [1:0] src39;
    reg [0:0] src40;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [41:0] srcsum;
    wire [41:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3])<<37) + ((src38[0] + src38[1] + src38[2])<<38) + ((src39[0] + src39[1])<<39) + ((src40[0])<<40);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf63c78fbf855848b6fb3bb1cffe20972285885a3c6f16ced2f7614c670f076f32ba8e5732d3970ba63d86e0ec8739fc0cb590e448ea6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b6bca7da5cc59b2f0d387bb069c3356c9e6a0a80ebba5752aaacdb51f2c60b560efd114d1356e6a3dfba792c14ee2503c0d1cfbdb5196;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4a69781f307b08b2f1e0af462ec5dd621fde70f2ea5446deb11a02ad618cafed97c80c6394ee5f2b8faabfd7004bf5630a1b4b7d2617d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a5c0a8c735d6dd8efa5fdb8cee5f00a6a4d9725789097e59a9ff5a5ae14222740f37bb18eefae4bf3b171e465294f2e40681b75da4308;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f90975801c911c80b2906299c7631750a2f5671ebfb67d853e84b4cb53419a14527eac193b93988316c264aeb8a85db3a9964eed5cca78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1edafc32ef876145121f6be5842c5789f09d7539398bc7b831df55c73fe3e6029d4057b6433e25da957c491f540d4af4257a8c27d9c035d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2c46901ba7ba4e9e986d676a68f16795245ec7409732a5858d86f1896d1217cba1f6ac32a6aeb8baa757e21da51f37f667f6967d01c88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6879bdd45c6307a99c8c0530787fce11cd745ebb258c4b24165cd0609b059afaccf13bf63b5445e682319c142106553a5ca6d568b70ce3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89364f1a14e9f837df9646adcb0ab7fdea0bcb376650ac57febc78b848c0ab863748bcb0dc84d63178740b88ec358516e5eaca5305abac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10dd589fe903a0cedf7a2301c781f78e89a4b5923ec7c86c0f49e16b86aaae1af861eaa0ec89cacbf3a132dda735fddec4f007a43a2ae17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h745762f30e35ca5eabd2c1a2c37ccf03d3b1253127d2c879c81f3cc7d52fe294076645a6c49aec7e0881a5676c06e28c02bd0710f2d88f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1846c1f02833b7b1d6b3267b01e6989430466f58fbce13483f08f2c1443b34f0135c0df8607f50c2dc848ac9ec6dfcebb5d423915d55f88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c0e9d5760c3f8db49f1c5912911250d6b052e46538d2026ac3df6df7274e27b023a15dbd2dfdd92efd92a8fdae43913df6d3c8f30a1d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2277f8b808e0d55181d99618279c3f39f33a5652f888a2f295b217e65db4b6be810527536d34842e7362b22b3aa32160657b7cb6c831ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a0013c1c9b87f9570306b58598d711c526046ea0e9b33ebcca72de50c129910356d118d42684dfa499af0e6edff2426b9897497df30a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185952ae53209d0099ff61b0bd680986f93670f555e8a74bd91ed1cfed0235ab6ffae8a551b88310af484da5dfb9f8f1d28dd4c1cd8798a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0d1941f2ec7662ea48b634f195004cb00f871d2e604aab6117b517a12ed5b4906633fc3af9fe1453ea51586ff4714c64b24e0222e1527;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc8d13d70bf56bf6176f316fc019115132f138b0f0e6b21a5138c0437f48b7dcf6957ff22a659a7fdfc5428d76102bc44f58a898901208;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7231aff78272922be244d1b98e84d60c5f7ab7937d69dce1a343cba4e8c9d7344b082bc4ccb539938efaf07dfca468e98cb4f85415b0de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha622066b61cee9e80c1a164a716e5e7f1fc4debc3ed7eecf5921283a8448bf1e9049021e9514d3c15fe3f8e117d410d97eced694fec700;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7bd9afb4f97936052d4dd0aabe5ce7e4de1a69f81e09459b80841d630504a3f75d6a34ddacb1cb0930e51faece23eef6c3964b53b2164;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfe7a35673b5c2ea95aec3ce2dac8e23594c4e5065061d39547fdae7e4a27328b8e2666498aa310529c97f54334552c79199b3462fdf32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33649edbeb4d3ee5d9915770037915b050b80d9d31b0ecefccd5aa962647449ef35135e6d172cf78b51eeb574b1ad34975bf35421ca26f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4acf38f982de9287470aa65f06a8b92d5661f89489a557513da65203c076b7b163eeddeeb3e28ec170115e89a3bc441913bf7dd766c523;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8e24feff97b0c862babfcf449d1babb328b10547746384b9fb0e97707941f3012128b200d408ca0dd3d5c54a432500e423723304344a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a106acc23017b9283e32aa8d1593890642256f0fbc70ec1f8e4aba3914f0e00570ea6b6dc8e57c46ecac66df7aa52eadc27426f7e3152;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcb46680ad539afce84d8aafc1d6736153d605dd038e5e0d029f88affa2c85278e39290d542fa663797c9444d3926b2115bf24ff0d642a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f28cf4760c964f41ebb5d8ade053d0fa801f4fd554b8efa835cb2472b3284b88c2bf5776a985c494fbad2af1da6d94784e28da1df3736;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5a5973d72bd67439a71c768a200488a9b73b2eb69e131a2b549adfd07ff22173fcb3a5eb8b12a2b50ef707725c84f0bc149d38c0c7402;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee3ae8d5f9e7605a8e08eb9173d92e58d95dc4d1b07e47e3cea45c99353ef9c3aed6ee0ac5e67e5bb18a7ed0d60503906ffd65daceace8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142ea102203912cba9994357bee0c5435c923e0dd2cb33be9a96b4dafef0a5eecfe12ebd8c01f8da48eed9a62234693a503a3ef9bda83b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed703c891f46d67c15f9d778fdde670f87246b0c709b33349fa2188ec9f5c8e5e17174e3db13f2414afd3f93a5b5e0b858f9af4a5f6387;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h323428fadbe5d8be28f24a9476404e0735265f1d50c698524e5f98f930d193d9071b238d3e01b1f7b7c5361a8e40ef3f173e48957e0e0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c4bde9aa1ca52ce156dc954702adec7363eaf44fda400962578ef7eb59aa1acd9aa2fe544778eafbc5b52234983f1ded2bac20f9aee28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d07439dc1ae8d7d899643ee283f007dde9a4b711dc6e039c81bbedc0f1c3825acef1280d37fb10e5a1f57ec57e659d68b51217afb9680a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2dd97436eb2aff0ceb5ae6f8ca65b9202bc0c655ff361fa806a0b29956e5a8343252d7b0e2e13453115c6d6cf1dddc629c8bf2a8e805b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9ef199b7f4c922da9ee9c73fc1e75aba69a18b49414b332de0be6ad3e19f1989e271eec828505f30ec7a224a81921d94d1fcf789c8827;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1961234c1f2c1f9ec478e1178300a6b68d51199d419cae79aab71416ce9dcf64e5c40b02be5aba3c7821ec97a91f466ffdb266c87c13b28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9abb2dd0bb50a1a56319e37aa263e0e94fa388986b27f701cf2ad496a678e438e320b525fa7dd48f21f5b0b973ac7790428de3e1e0c41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b41874a8ba1c0bc6c0af59fe768dc012847423c30bf1da69211b679d81f481cabff358dc5516439247b71eccf0e08beb1b03ab0f525fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7170b437158a54637df84d77a4b475917082114a51f54217c4c0da339dde8eff4bcb5af576633bc764ea22678c6a1ad51e5463024fcf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c5bf68a7ee9c08cb0a908f231f76df7e9616fd7ec156e63f9bd2619373659960b04c3e9e76860dc2a748784ef6a6d3971aade2a2982d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19efe48ada8c2babff77e6f12c2b3d3f62534f16ac6f0e372a3489cdf087ad007ac61124c08d4b4a7d957083331fc5c20937b898cd60856;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164b605d264c19f071ee0c07dab07aadd206bf9c79e0ff90bf2e7187a3f08de7c669a4e6350323e35ec26d7b1dab65f484e6af78a0d2fd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae3d9bd952745ff3efba3cf49c48db54ed5ebf1e394fd3586c2bd9999d24fc0cbc3233f5855229377751b93902e45b8e1a22480f3de9cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ed96fc6297fb47dd0428faff16008ef57523294ff91b45da6d6c1fd705fcb8c04cf81415b9ea682989be320d6f0033dc4ca0c0344b569;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43c276e48f82aa185f457b4e9f562e6d17fca9cf1e18081b885d680ef775198b2eab893d66a93f0e467ccf5abef86b61465960bef3b6e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24eecfb353f5c7eff2f094fb466877247980ac07c96c7a34f0c4392fd4ba2d5de928acd26d85f86019879e616ec097563ae3298252f62a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4cbae9c6bb8de84dc12a4ecb59a284ef4f98b3b80f89fd3db568225f6e135b4f1a2961cb01e98a589658d96017d4764c1dae4bdfcacfba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f87d6c2331d157a18c29b27cadc4e06ef9c47188bb29081e11ca743120c6036a4d6a7cd55a9c8e2f4f07add3dfa14a3541dae91325889d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he58869317fe44d47d176745b299d329fe0ba6482bbbc2762c2e532adca36a32f7b38b9e223bef73808a75334c80f353f019c3e503d6c7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4baebe0a50c9467b39d397918bd708806967acacae866232865ceab67598d511909dd3cf990e9371a929ea94d5184524a30f4d4517888b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cc51eb319266a3caee0dd30cff39da58b4e29298f52e56dea55b5d07d2aa88300c6762359f664def1dce8c6d06a2d01ab4fc2f5eddaba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c22b51880fef28f922b86c0645f527a7313143de8ac019245d80805b0fb8c2b34860d30fdad86b6ebbe87f01674798cf194e3b3e83cbf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c401093df3b304568c7ea7f21ee0ffdac593fcaad7762128c49aaf7e375980c4041d0ebd59a39c69000d1c5478cd48dc22ce69700e6382;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe6d00421429934bce0eb3140dc8c34e8272ebc6102bc47566cc752cce4ce96dad5c2590953cb1ef9e676b026b711592ff2109bc3a3c91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb463fe5790c1cb2707f29a558388355eca46192ea74576bc71cc5abb39f1e30f190e9a1d2537bd5a2268c9b5ad0e4ef965a223e9747b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce13f42bbdf4e74f256f22c69f30dcf18aea91a92f4951817db5ce32cb39b5347700e5263d2beb21ad14de607ca0abbcf1012d1bc7fee8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d55a9ad48ce66e0dc3f08c342f71f060baa684fc164fe4a9c10330a42c9eab7e982caeba0587226abebf6c2a02e23d0a5c601dca1de6cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166cfed331614108826a09581df1203b3d8d14083abd4b80b88d707a03210ea5ffeb25c1b4afb582a828135b4d16df58d05a9cf7cea41f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h115a68feea7ecf177efc7b119fb488d091fcf94f9407c0e46d323e47d2d7cdf910504e3c425e1729176b1aaeda8c3b67151b9c9b29514f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9656041fb6150c56ea95bddcbc32b4e0cff9c1fabab5a53e6e037ce172eae8175faf53be42a26620ae4d8a16fe0c6e2e35a6b9f292753;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73d84aee83705cad068ca06242d71209876fa14334078af56dc80845bf2e9ca4d63dfb18515bbed0625385009372e5514d17ffe0d66258;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7916492ad96fad23b5f6ab2f4006a67a60ad5fdc01b56a23bafe008c3b5f76cd802c0b9dd2b2b72334591cbd7fb23f3ef62002eff86fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11964dc525da25fe7eec33fa37f5a7168b0125d57e362c4a0aaf9e5a8b6483e991d4bd62ff3e9e9f2e0ca1a4729989c379cc4dd6d619eb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfed47b9155a21d7ad194f2f1bde31de6030301b916fa51620baf122f23229876bc8a286fd44df6ee15d43514ee4317ca6704f3dfec8bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbf3f492a2599e103e54eb45c30afdbe5947e64c5f1174677ead0dd307c4de6899e8fc20df9cbf06d342ca8ea81a1007c10a90117a6341;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1669684d05c3e5e9e302455983d29b8e6f8474be2f8c98ca3a3c20378dce25c5de0ec4a1f99745917dca50593e13403782048b446ebb7ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18fa0a4768dac4dffebf7eb23fb8a7483fbd9da2fe444803f645418167cb0ffa274af97b1cffbd366dd2c510c612a39ac204565132f19b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8d70cfd10ec79c1e53cb8d5f46a7f59b48369a0b9801569007840ce3dc6da9435a55d7cca501e1edee5aace280709fa28319d8ee75fff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109686695a3322789f7d16a39113b70e2300caf0edfa5a7b5f0aa9cedcd6933adf11ccb2092fc904877fe4a5ac06df82aa5209c0a278a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h283358ca261de04440222621b5cc6373892518ac1dcfa44d2a97f3984b6acea67d41ca63d888e90f619b16f1a209b71ca6d2549f21bfde;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1218db02840cd35b00b979af32b548806985b1adcac79cac3301050b1c546c554982ac5d92678ae7b394c1dc571718808b7f3f3474e782d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha66a4d890bc1a0fa223a7b2b391eb6405989850cee3e3553aef68ac98f1598ca59cf0c06739810ea4ffcb905aa8217c8f060bc2eb1eaa4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc039c02c9ad4e138add5ef26a7bd9ff48e55060c4d5f424ab793556defe669e5e9b3ac4b06deb1bd8e398e96ecdf5c686c154bc38494d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5dc99a204ba05e383dfa220f515058ad8169c1a1ee4555cb16c82e3bbe0ff49d857d5f84e3283b78e50a3babbbc9a89decd9a6fd4be2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c29cd11cd7c574365128d69534cff386f06c1a123d61bd41d3e8a9476d02b699a633325e4c0f09797176b19b26179452146dd787199b65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h977ec6ce3caa0377bcf07b388bea4016cf8fb5a5dc01aa00d0f0e6062d98048ef4a36b279cca1507c96b2ae8330f887bcfffee9c02b0ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfa31fe781c6bd97036c1aff515000887e7188bf7ffd4c64df1e61885d22aaa8eaac0699ea2a135d37e1f98578b4d2723a7e74a700e3c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd890bce1c5580ff5ca9089cfb5b575bb4ace59793b67dedee75c80d0bb845447d90e64c4d197b52825bb2be576cbd8cdfc4967beb3ea34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1ab77637ff0826a6f59c7a73d71e0138a1c4be850fab9fec6c65dde12aca3e4c64c63c4bbc4201ec9558adea52edd252a2f893971eda5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15af7d02eeb2c6331b2e0b27e7bef7fd3d3ba996d13df39bf87d56e5f4c01556555539fa8d5ce6855a862bc969f36c2d8f657f4985fc4ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70780114a23ba7575c2725945b63f5b5cac75ba0780c6b389288c32465c81634f296c611050fa1711971ebe02b64f28c69ff8ce890ba91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192f288774b33e67ba834d0894e1b4f6796c4482af539d6f4c79c68ffb26385bb3c5ce1536f25fc1473bef890ec4f71ffeef3bea3b6caa9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126846d57d885d77c199c587918d2250643be1803fd74d9915cb469b24131cdee595f938b562cd47a8dc3db10f61312f3b3dec634cf4a3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dae29de417fa7e1ca7e1b4a741350c57b34dc71c6b8995f69573322f1932ccb3eadfdc726eba3c462b8586b45114dc8d8ec00d51954ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfdebc126d513f57ec871c845067e691bfe0d64a0873f3ab8677ea2a45ffb73bf7e0b1d2cb72339c99d68758430f70a442e6ec843cd6a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7140c8dedbc220d2c5ca45506c10e56c6086dba3561ee7e2c6e2e15ea73eb6c0c58e5bbbb3377b42c838912d00f55f553ad617f245a836;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5b695e541fc05780835b27a0334076e1406adc87265230140b50489491c036d2d7601a5ee1ab92f5409e97441c1436f9ea276fbcd0c06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181b87c899130b9c9bdd1831b094f0c84e5d04537a9cae966a01cca81a74981814c47b41353b11a19e0455dce724d94dbab5cab706224ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13daef635468b02b16f6b94df5be520bfbe3d8a927ed33d2f2c6fc3c0d073996756c3936e368c497d6241523303970ca5da9dde95831463;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18854663103aad85d8b5a3f2cc63a12759c92ff3d5bce107a5f25d2149a3ea5e14b943551a12bda6e36ec700f9defe34069c5ce25225488;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0acbfe4924f09cbadb069bf5594580aad9ea0d76e0d3b575a85b79a551780f69f566615ebc78dcae35d8cd527479365a37c28be8f313b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1651c0538df1076d6118569847302ef67a858f599890aba2d59389f32a27e4d7d6dd064f849583e4b3ed71c05f0f7a54f9d36db12ddbb7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d0c6d984c1c3099170f76b65a217c561ce95409e8bb8ebbbc3fddaad4c4e72c00350aba488c6021713fd2a77ab6acc8a72fb3a1f1c791;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0a0625f2248c1f0a981e62bc35380ed48b8234583135a189ba55b394b6f1e2337a4da50aa66536380f0e5db325ee9a894e3d7e166cef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2f362954f6e7381c37491b1bba6797b265da63b14482b7859f0fc29cc39395944171f2a436d6a41c100144eca1ae34f236990f82b5d53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd91784f285135ab34ac2c37b3039ccda3b84251f480ecd6c101b8b7dc4cb1888d47e0bf168d15904557b6aa18be3a6bd30c1d3d873bdb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3df49178f969a9390e860563ca24e4c5f759b19ac73abc5cbdd0c8480bdf170e49c91b878ec9921b0cfaa138633b35a1c7481e4ebe35b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171c3d70417a3754e7cb3a1148a0b9f10b1fe67d85175e8745109b9bb29d23df1514afff7f8f20c35ecc4f9308a1ad92ce843d102a6ede0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9ae65a7d4cc7216632de882b8a5ed23ee5c0e68fe324750aa854be91f00472f6dfbe5a92dfc4d71ecf8989d65a9d531d4132be33d06b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f19b6d3c974f70a2efaaf75c96dc06a84b7a333d40320f12ab2ca35cff2bfc0ae2f34fcaf9cb9390393af4bddc8d7b33a94082c13aef00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb70f266db0add1ea663c5326d781a158a7cdd301d534124f370f3ad31201dc8a00f60180eaf7c7f7d5b01fb310c044e78b12596b71779;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca887e062679c8aee8b12298596e18ffc130aa8abd1e7cbcc2821e4b41c3884bd09cdb57be3aeedd8cbaad6ca3cfab916710e4299e9883;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd89b9ff32c80ab484b01926968801b56f8da63182955dd956da5b38ef64dd6ae3efbf2b0a1581b0f70702a93e428dd8c27f311ffdfeeb4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed0682960edd8ce0b0c5c508b69c92d60e023a193904a1fd70205392eb05371aaa0820729d615cc4029aae6bae2bbf3c238023783de61c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da221d55d47de8c7cbe1a88589aa1244bd5dd92d8d4facabb54282171399ec3fde3c96209086b27b45521bd833ddf45c6a4b7420ac51a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee1968607dceb9d84d4edc371bf6c103ae59b750b49f8108b7e9e4291dc5c7eca1339416c152f90b848f2ad5c4af90f16c213452cf3d8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e9e0dedc0e0278d03f13789f2ab80382226d54dd1aeac7fadfbacdd7157290c1985a6bcd03255a2901c0ded5bdfc9f11acac2c20fb81ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15758d06c05ff73ca939d99ab9ea2fbdecb4d35b9aafbd639467f8a432195f6ef7d9fc83a24e26e401a4e05b7561d22a00fab4be3a9f3a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15deea044dd98a65d5756296ca6fb6f7abd98d037107ad1ae896af17ef56bea11325f27e8aab4ba3569718853c37f1ebbf6637e18ab56df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ac22436ac72968ff3e48577aa76f5a7fa66bb20165e45f903092b0bdcd26340a2eae4c50feb815b76c9ccd0edbd6c43d271725bc255fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee80b9fa87d15d34f5492bf8996f57ec11be3d0515adecb120b0c38d709012fc5bb707e80a15cbde1a218dfb8c1262824a86f9373fc6df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeb3db0eb02a571d6b22c4f5390d365f55ad0efe0f2049e2208a265bed899c0d37b1001613ffe76350b44bd4fcceeb90ccb2bd827016a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63e1be32779a966493cd7ab9b7fa63e24a72c67fc489db5b7c5f3ed1d536881b8fa7c1aeea1b1f016fd61d786d1a42dabb137fea426755;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h866fa3ed553f80ee3e50014048d64a9b3208e1ad74e816b4c101b8f67fe97a3e0ea19c79d1866c5a76d17142d338e65b81d12520b66ab4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb388a46a9fc987b50fca296d2172b9bcdc4f391537ed7dd55058dd437a9eac9c1a1578bdbac51ebc9ff66d7de086e15f2bb2c2eaa2ca0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h664867c5ffe5f368649ab9179dcb94d2787388c397360f4a87ec5c2cd1b2f8bb33578cf268e16a1fd69c522305f71058cd2dca28a55df0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fc4138768d71b7e2d4d373127359eb8849a4dfb07fbd00cfb2bb5db1514a25822cab65c4a980f1f0691fc51f2dbeabb973baebb86f1ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1394c42ef2c9d6d2c5464b48edaea8bf6361a21160b2a55dc7660c8dddffafd11b1c57d208cc9316e15305e377d0a6b5fd8a7759902fb85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19853a4c47d79ee175908ad66eae43af3deffaf70008eaa8928bcb6723595d29f3f6f28934aa4553ea86693a076d3fb211e01e5c0890fc3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf217b8f6bb69954f1dc60c7c9cb6615b0fd6cbf09fa09d52069c50b18fe94922849b8d0f8e2c2ee568ee7e2da7e5640baad612ab38d7b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae64913d6bcdf45ff14af485f4e17d3f1b13900e0887b27153ab010cb285e61f61b10509d6e982c9e6c9e48c759ad6c4d2530f247de9e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bad90f7b0f991fa8283cae30aae6a7f3b9cc113abb0ee6fe474788654b10af94842678c4d9d3fbd1c6240bf87fe0983cb20097b98c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e48bfc6a6a205b72b5ec075227276278aa814a2ea2e92007896346efaa28ba8d116f35e9c51394fd98a05b8c3f4f7032e4e22d80ee8625;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6f622a4d041a8d3805fa63c7ceca642a8c1020ff65b03bca187049e37985d1d56ae3b78390e7c15adee6dd369b67d1337ad147d6230d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aff84f9bbdc26509b048292fbdf81f3b076a9afa5f18e775d7c077f35761bb5b83dc07184a981059a7d77139a85acdb3cbdceaecc92fd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a325e448c46d228341f69879a17aa3b29ba327d612b2c6f77dc439f9d55c39de37a413ef7e077a6b01e3c8326c66876d6053d6023a086;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h896f3f19d6c082805333aa6912db3b027c34814efe6b7f2684364d3de466950c92df4cfa582c78eba1d576d2f28833ca1927ccecb27986;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173cd445643da8404910dfabfee44a682259527ec731e6b7749afe14d99ac22f0b5cb0892cfaae0a8a761f059d418f84658fda93e9cfc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118c973943faf7b56191a67fcaa663dfcf1db6b9c8c1989acd71d5e759c1c593c89e7f6ed7999e3815fd9267ead89fb58bf4d98c88ef67f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h311fa1a70d59a84e71e503403b125813c573d54110836e1ec50dbf1a228ffca5fde608e4de5f0e34cff6ee1a7628a9351958dcccee566;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1559a57b81dc280551d8848434eeb70b8d14c475561d6f1a65c0f3a2ed205bb8fad2bb2b48ff638c3bd1ededbd16daa71c52a7f3de93872;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6c7031b7fb7be55f7753f79a3f80e5a715fdb1e4f2c2b39c5ca5aec59f9b1245828c9213f9ef34a321da497517bb0262d9e720556cf8d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c38b315c4e3e96091853f947028897cdd00424b8897a0d2ac4942c3fc1a330f3456f4eb99952d12d30c2c667b61010630d690ee79c39a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157e5e8d35e9f61768e945e97d2348326d7bec0face2fe8c990221f139e4e72bd28cdc6808727fa6520991ee43c70860ecd40264358c206;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h893f2f9fca275ef10bd7bc44ab2ee1066915495787f4f6665433b85b86acc5b9116dc33fc53633cdd2536ad17e9b3ae2643dcf036d043;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h956608ef9b665404f2e0fd9af7ffac78543d9a12cb0fe9e42c58a5e541588526a0657b0c4cfacb882121a810ac46e0ca0e3b45e182c310;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf289389afada45c59a37a503db34d95169f82ca1470a0ed829fd8c1990c61e6ec7277f344b6b9401c088845c00ad499e19adb095fb584c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1692c3520bf4ea8d3c7db2e2c4d9e6134df6b373946dec2571ed5eefc8409df81cee6484ab63000c0c3ebc962b882dd86e29b830e5612f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3a5395f4c37f29460a643b64c5b7f87b5962f538d8512d046e1b51b117ad4f395ed3e00b23bc8339e540bddd39da7aaabd0055849e5ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heecaf786fc213a1acadf6240d51401717054aa628f60fdab44ecd239a060f77f8136f6860fb5aea00ff6d1a56eb1234e35fbe117d22816;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd98bd9946b1b86c1c29fb1c38dc196ac4f4cfb441e36a5ba0b5fd68771564908e26db9afb45e9b9f4ac985738ee0d12b6d92c9e084dbbb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1459cf1f42362a2cd7af3bb8b9ee4a6e5a6449313303b0294684b54d0537ca027a611148bb5ef9985ef769e4e68488ed10c50fbe200b0c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150df48e747b7eca7e0f82b2112ee72398259ece046fd68c331430ed0917f9204aa1075c1d88395c3301bd63d131360d4654bce260a0a5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116a2d22a6415d3852656b43983e466589631f8f1c14af7024e221b17f698d02dc459d5cb08667df30b98ec967f2a70dfd285170986aa48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13285922671f369fc1e9949fbb123ce00cae38ab0719c2ef80f38e0bbf48c2a61c3745c5624bcd39b141c225d10193149d3e741edd30201;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66317faef6f933b04699fdb1bfc8b2e870df7c026bae8fe0022feb3a18c8f7782afad64cbc6db9c7339880f49c312226c5560ffa843d39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fc63fb3ed48aba766f35215c09b6f80ddfd90aba7b031c71ff912ad862b696d3361253e51757891257134d6d2444266b29d24abb0be27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e9bb15f1340fd95a4bb7e4104fa34703a5298723a0f0527ca7c78f196efa5ffe34ae447b55079c719091d156b7c048663846d191486b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h629b2f2276afad95857a65736ede182c006f381ce8d400089c299cd330103ffe8e266e138250efbb977256e7eba026952d63702f64e461;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f158de4fad515073c7a183a517dd74b508fd9071dd783edd361e3864cd5d29707808940599604076c34c856588dc94fa910329091c11a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e025e500ca0d880131ac48f9a9d349471665cb212b963934fcb1cb6c5d5b5e25f0e02fc51211634c5cd9f9df2a109f306a48b19f5a4e09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf71dcffa527b55725095870ae9ad42179e3cdc2658e54cb5c7ac8421875f80df3cdb65882e8b96262242b4559da94b799e116593661ebb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc951c89deed38a921bd1085caef6a6f72b29fb0ceec8418afe4dc051d8c2e7f2615704ad7e063a204601e95a6a0c46f32ffb635afd590e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172a60e97b19e8af178bd367cc9825718de050b10a187a3a45aa6923a6504ad7b7bebeda231c18a32bf3ace71d3119c2a0d5d970199b743;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181f8eb2eea6234c958d9670155acb2cb22b145c1175d5b3257dc44e0a10f5d3b93ac397cbf7f53dd11ba023f08821517bcd7b725ebe107;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h662fb4df8839394c2566eddd2edb7778aeb8a284b6691da57609a1099865f852fbbdf24e641704031372efafdc4c6a61efcd40889684e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7223575b2d837f53c72c1dbc4f0ff62ca9cd0ed784cce80259c2e09756030070c8d7fabc49cc43c0a6c9bec4e05b69927e397620d6476;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae33d721d6fc2b227de8b23198bd00118396a1d594bb14f030ee26aa7be3e50f29b8dc9ed0cec87019c6af178267b7bc2404edb4347c45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105cb5d0640e8049af12427abec07cb5426dde425cff45ff95f4f5195db02115f8f72e5af2563ace73cc09ee642f46fb870a5b94f078610;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd38e48f927f092a9ef1b047970a33063a17eac44c088f9f1c6611dc59dd902f801cca9db5377499ed621298e837f3ff3efed405cfeeba3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1658f17a63e6f12630c200eb665c2c14f919374f9fa1383c36adf4db52ea34291729369b78102d072f296b70f76f66e62296085e8965627;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd307b4a97f1f9b26cd2767fa48948dbf5b504b56826a867932e3c1f958d6274bebb00c107387411c019bf00f475e2394d24e775eacb58f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3f5a822cd042922b59b72fa8e685e91f86b9307b2afffd31e09c02c3300dd261fb10824fb8502ef460fc82fb2bb610b4ae40cd82e5bd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d6ecb669d1c8a810f46da208038187baa635a3029d47dcbf996908274e0fc0ad677b03a8cb6fdc3524181144f8076fda3b89b96960199;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19d2c1b6d7976ae097044d19b26698e56dd15cb309f3ed86edcb9aff9ab5de272992183902290156624b08e4e2bab69bb55bd39804014ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccf6c883c0d4a157479fdcbaae1900cfdeb1054104a00a159eafbde93f75ea8b98e418244d81969ecc5c2575141dd1e5a0e94f94880875;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10667012d923505fa2910b8e7fb43abeeb267da7bfa8c13cfa4a80fd575b4dfaed9cf86be7d9b62f8fe1a3d73df71f3fdfe37a18d5c2736;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1234e18040bdae2de3ae28f8327a9fc4639af4c1ad987ada72ce213dd8de1ea428afc075536ae3f6a057d1a1eced7b3fe9568b7c1d2a07e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6f45133dbff564efe1d11dc74c334449dd0bfbfaa8482c824837a27144399529a97dff404616f46ded01c125480eb36251f4b3f5bca8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c933af273f4b39df4f0fa8d10219569b34cdd2f0e1505941d0b06d6d28569ab00ed766e60b353ff2e9d330ba2f69cece506905d86adf5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34c0881ba8725ccef99156af697fc58e76d41cd41fa242e3060e3fcd3776c44670ac8c7734e767ffe8c17be491e86eaec32428c90150c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b73fb8d80c87c189b8b849a67c5961cde3f1753fd9071e455e1331b4e1793c015db0198d165f3ec51a58a099bd9c3b014ea38863bb969;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha700e105e7935caf1cc2e10487cae141234a7d9cc60cfd92598ec6bcb673d0eb64a4e5bd70efe93210a6f736b88698e46eaaa73c3e67c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc29b2ecad93700d360328e7158ef4f7f4093eec370ce891ac146e93e168f2ff17f8457b4a2d9b8d2a85745da87c146fc531c32db7e8f54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h789a19f265ef8e7086d0a036cb672fc39e23fdbf136e2f7fabf401b22e5a1a1ca3735259f0e7445b6763feedad21c61210d162f0d61bfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102bf8c0f4402c90549f3e0c33d52f46b2426739e92754c78a28c2dfe556f7071535feae9770c9ba9de628165fb94269a2913f4cffac907;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8b44a1c1abdc5ff488129638f1e40eea4af82ae59fa74533696c30505fab495b962907addedccc4c600508f5d19580ae8d44d7fe8a421;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee721482f4a9c9f88e740e00903470cd4c5feaf3bde455afe6731d12a6934e331e74cce4152366ec8938679b79deb4b95c2199a799ea9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0de97ef5161ac2e1f52ca403600642ab6f9a01c1ddd836e4d3843c4b319693635164eac6c8f667f6e382cd2a4968a8f4a7b073d89e8aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha228912dc6c245777ea996e98bc40aa26f471d73a186b897bee82fc6b2638b758cbe4f639f23203234b21d5549825df5dd1adfd9e0a9a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bfa43c6193a72aa2b65f8dce8d586fcdecd40e72d92546b59bf8791c3491f4a7c5014efcafce70dfc810fe71564ba85e2d6c08debd96e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dca6dacbb400e4c965a2e2694b86be3098a6456a565bdfd9ba8e4c7dc2ea9d947eb8d0eaa7360f60edcb7cff216b4c28a0d59b4d908f6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c979c427071d31c1f5a302bbf03406f8f4b983d7907b7ce9d47d62098531a7da5399481773de26577690230c9cbdff506a7008203ffa2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145c1e3eb2c1151de52a79f63f6e21ae52abd54d9179a1accf3cf09cca41e219bf08f5c425432409f9a9f9b1816653f16ccdd9c2bd9a98c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11418dcf8ea10f20e0f2c23497d48ebb9197bbbd66ab3a2bc5498802e49172b3a5bdffb6726b81da02c3656c07a1ee3ff37474bf8d0499e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ee091b91f4a3077670e7d40d9769e9afee85e637e263b6de54275bb92ab38cab5b4e90db8077a397a875c8114e6832bdbedc799c256ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7503eb8e92ae52326784a712c0ad80ef33a014386bbd455b663e63069fef9bf64b365c379df0722c5fb65314648c33fc0453983ebe78a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12cf41b69a2f971ee82324cfadc8c6d5a9c234e6b821bb26ec2a1b24deb3d5ca6578bfb1ee8d67870a7e92a62cdf6175a74a0c5353223d3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ec90b9453276111c4813d1fb22d9199d2365b1185157f7e2dae05e40ba9dcaf72a1f7886e7e5c415f71e10033ca876c7b310d41e13447;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha864979f10632a05e10d28a2805f50ac478ec73cd4af9ca70ea66172d8e60ed6e305ffb0a9e22855b6d15da1227543e0b14c7635da81cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10649abbbf6a25debc4f2152f3592a9bb2689cac26dd7f7f55e82131886d1beb1286152d3a897e305765952208f6b339a3dd1f92e5014a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9c743aa9cbc852a7a7135ec2cbd4c02f831d139be0e4c5e496a91d01ad354a0afadde15414e0ea03cf2e38da5f5241603023dfc1c75b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b986b0dd8709ccbf615ee6e21fb19056f8d3c1097602466724c6c857a178a3adf87fee7a3313205aed86fcda2dbbdd17f055c27d9415b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f05042f23616a4ea5f014e961846315c125822ce0dea9cf0d171f10bf3eb82604ad41aaa2883b292a58dad996da279b7b495417d13259;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba84150e28e4583e430d9db96e6804dfe1bb632f2e1ecfd0cf1690279efc413184e3565ef951c3932441a9a79ad49f1edeb6a2417e100b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f14e1d6057d16018ee46f805c9e414e24197859c2bad1f3819c0ac1f1f241442f7c7543c2dd10f5e747e3db6a57e1c903a281389850f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c2a5fd5a6d631a10be39b0a7a94303fde7a7f89bcc1c8b217574fca594736aa13e64aba518f177097d80a755e6a83282dcc4391b31c2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4dfc32400a5351b6f64ca26add61f524b5f8ad69edb4d4e12b9a0bba2201ee59d429950bf81e267c916b4824da57c6cd64a2d63e8973b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h378d1a1a8082af109c0f5880bfeeadddc7ad3de2c588d2e0f0664bdd7075fd698aa6e7bd5346593414479c5944176be7f3f766b154bed5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6cd0b256f7cafb3587fc6046bdb7c71835cce600a95359afee14f6070d9855043e55e44bad4ca7cfa7ab84783d309c7dd8e5f1decc580;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10660fe3c750c0b1256000d0655a6f2142f1d85d32045bb8942f7d060d29567253b5d0091b901eaa90e428b8f2420df6befc3ee5e4da6b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha249f546f6e151a6946d65a858770a115456da639d7b7d69175391710428cab6cf3cc786b7816c01d7221e52f73b878c4fecdd530576a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h280a43373c619985f27ac5842dc1ebfeddcf8c5ec95cf627a87456ab452d75e1c1ef303f7eb22f993f6d9e29f8a02b0d7788f9283ffad7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h206f195eaf74d508911440907bf24e1a4f157e98514a0cb9a832e92f87a7b82bdf5ff22ef5a80f0288467782590effd0e730b6084fb2bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c17b4a376a13098199ce60fec4738137268476a5594b34d4678a7fddb31c3fdbe39f614f4abb0349351d0344604983bea3165b58e908d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6bd43e0c7e2dfe8072448511b840c5938128614e5e304d1bff2f7cee08e57e340a859ee1cc9d7dfde5e9b8b7acfff86f1c47e4f391bee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7a7a1766ff54253d776d76ce293b0b827b3776b0a252b2e78960b89a872e43388b95fac31d9f3d4e9570a51e3e23786ab74345d62b8a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1339dbffd03a4f76f2e148497f3b8d63771e5aa50a335ec8538ddc3d19d28c8797576001ce1d6a58e0cbdc139977064c48b822b9a40ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b1eb2782721d0258a2e66bdd7def21039d3fc0c7527514e1be5870f683a634fe0f609b3111027d2a223599c95a440c2dec64d46cd6cdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24631bd452a303fb182b3c5f3171dc3c9945f644385a58c03425a79aa6127f68086c6d627dd14c2dbff214b9e46befed6c0c6d97b4cf9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd3af27f5b610324e5fc08ae56da5fa42b6f5b058d11660554f04589e7a2960c0964eb5602beada67fd5753d46e4bc0122c7ce0adc7f01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb219c0ee84ad9b0a0124f169378f15f1fefb5e26a12a2b7f4b776494960d28149ca44e53108cf221f37d66b98f2f1be78435d585ec4ad4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14eaba6cfb5c1ddfbcc77ab378187014fd1c7eb6e0652c0633c734bce6604c6bafe82eb5cde85bcb63dd1a743d6cfbe482adcee5584f979;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dacd31203a72fe013a4babb9f5a676ec3f10db41da88786dfb564a040719877741117682318e736da509acf7ba091fbf5634cd6a5d82e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2c2556eb2e8ede5cde55bc423eaf541770e69c5b17408184ae01cc4086d79b5b41df510432370ce06beb69eae361bd1d59751a995b6e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dd46d9b7f9145de1ca614016f838ba0427c1818d7bbf05a1b51ccd6199c18fc4e36af9cb3276720ee1e553ad05837e70eee59fe435e78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6028ef3f6ee65f2889e5d71391be61091967a2b1e111a95afdc53f000b510341524111486644a592bf4f2fa9cfcf1aef7f8c65723df99a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1961cba0f844ab82ac56adf289398b8d37a1cf45b1d52614d14fd3abe608d9648514327083191ec6c05172e536c70b01f446618758507d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70414d584b654393dcf21082b31b6084219d64d3467580828e560448c86a8bf0b4712b19fa061b5ecdcaa89876d391d1a1b4ca892f3bda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1383c407b9c176c249ef9d09b0d3bc050643eb04c6617cfa7ab9646096daad1dbbf6b8d4da21edd78f7ebc1729bde5c012913cf453a0dc7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2f02d0d4aa334f3a2f6b3760e42b14fb9788f162d953c821d2a06aaa31c678913c08eae6145c8ca93e1ca1b29727fba4c77e2dc57f51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76312a500042021acdb662bd9cdd46715f81e2af01e375d2ee66b4c6ef0a6e239b18459f4da23d604b0e2d7c972114eafa5b751591b18d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he89be35db3deba064d64ef088cbfcc4e8433a79c042ec4b97312fc44711d793210983a3aa8c9c1dc45b6626953ac88de9b2f10fc9ff0f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h767a42da83d70d51f452055646d2ee2b42c3ecc63b419ebd94aa750e07f15766b038864943c9c2250cafe7d21d95671c4fde784d3f45ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123d5f4277399af89a09cedfede76e720d054b91a8e5686a9e0c1db0eecf99def1be4296a6f333abec8bc8acc7721a50a110362ac9f1c18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19955d30e4ea7392a25ed49709a07835bbd40238eeddba7dc6ff5411bfce820cd4633a31a4a83fa1dc63184295ff6730579ea9e771b5ce3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e2392f570d3c5c893ca58b35964e886cc73ddfd716508cbc259ab9625c6cfec5f6dfb605b771e93e9dbc2c0dbcc3340cc6ad1bdea2a3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b1b34f04f4bbd2960f6504ff75370e7613b5ca2b93366570ce4711b0e3311095d66c91a34e0c55d289efd808674b2132a8fc8d2d96942;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa9fea3d680fa20b33a7511c92389d9467d55550ab86e88344fc6636d5bd3286a7022ef1ecb8c0f3886fe3d084c7d837955d70a3e1896f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39b1c102857c3cc7c20139f591bdf88117a6c7b8316f600ea44d970fcf4586f5db081e2856feab777d9f36fbc38fd4d335a5bd8161fafd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19068b7189fd5b8fd2be4c649153b23f59909f813f512e1e46c12f8a84d69a67b551288f6556ef1333257b90751d434362fba4910c64c40;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7ada934f3e50cf83198a6d7f6a862561094e93bbb484378b186c19c5325527ef56868f3ba726e322df5a31e493b9dc0c8ef94c6eb3bd7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8447edb7e93e2725de62cfb96e3e82b9d4ea0d81efc357c45add1d2930eb64a094669eeabac936ad977f5da33f7c8c25b05ab3a59ebcb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dd2a7f03807492724b5cac7ed4d793bedcc9b561a06e1b4b3ea0bb42e7df5ddb9e8c2f71ca195e6e6d694f2a596300290b253d1075ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1515377c65ab54454ee9fca638428639101ff24a243d806b6edd01b8e472ce8853bbd3b16e709b9ded1cbe3b0440a521fb2ccefae9edab3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13dd1089dbf940900930e2a7dffe095024b7a396f316639fe871c5f29406445ccc85e99d4c26a00fb9deee748fc193d20718383aa665c99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191cf581fcbc17d618578e8100c186f3346ca73adf8cfdf79e1d57f1b0bb7eff732ff0592c95e7c2ea2950a39a88ad3003f754868bcd95e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12112c7f850be2761aaadda857faf9f53e77aa7db02be6bf17c63e314e36cba68545426d64b80139a83d00116d2c2e4ee79ebc8eceb2c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c406f4ce94b315db29819266de79424b4e41f05d7b558f7012875c567297e2acdf1b542a6c01ff223ed48cdc9e0cd5d1deab1b3503c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1738fd4a0a0e4962474322eaf2f5721d805c40820f77f99fb89087edd79ac1c23b7225b357a528fc5c3c4f1a3c26d553c401997bbd58712;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb698f0d09b4c91569623e4bab3b001cf9f49b0a5c915e4f0b13fdd09a11069352309628688e8d697f6774eb93a79853c626de4f5a5bc45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6457c99dc2fc162e4e683cac82117ceeffe83e16c433bf74e06bc9bb3afec7302f3ceacc90b04ab5335fdd89ffe35d30397277fcc78f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3832b125437248838889f3dc959f505fc20648f63a172b89e819726da1c7c2808b8c9a607a91f4b00f5a6ee895d207b7e2e5c5caca5e0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf8547ef4e91a2b7a5bb96005d9e28a006853ca5d90a0494fc8d44427dfa541897783d7cf8fa20151abafe3323a95a70201c3bc534c9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab3673f9f8479d6c8b9a07127171797ac90cdfa5c43ae40647e8c304d225802872c42b59b0c9c400c6acabb72482078c228f218fa20097;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d0d17cfd64fa72f26b512993ffa4f60d6affb365d1a1ed152aa3ce0031f6e78882bbdb52a0ff87f50a97436690549ebd67105bd953941;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1403e19312da61fa1e48f3b83eabf8243f727406bd4b3d547aa98dc91531f5329b1aeb3344902616ca6576c50d839fcdca76f469ce0a90b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbf004f2c44a53cedfc44df90ddfd9c6ba1d104026e22a40929d0783ebfa4425452fd6283ea40bc380ef30e1c0a108c242b23eab127c03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11226686261711680679285de561f225260c1cb8453085ed76ee75f363c9c5514c25c76f7a79c10a5c00405ad5e01611b322ae93b68f77b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he50e23045ee7af4a2d7cfdfaff61cc1bdd070ae663c19a6a8ee1aaa64a40dd00796a0f7dded61ffa9c1b11a8613e6435ef9ac5829fddc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d8ed511782cded33b056022761c380287b5520bd53ee51fb2afed6ee231b65f67b620e9c3e0343a17f9cfcba39d3648b6dee5d7c6184;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133baaed3296563e4ce29830e71814ac4a88a7714fc9547e169a63feb6521d23656b7b07ef78c64df11f8d0c75af0e21ef6c9bada2f3a73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56b28204657e4030f27b4287011c229962fab1c83d106f4d52d13977afacf92c0110d2db85f0906d5280c2aee8d921e1ed4f6134f0576e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dbd4735ad64c66d3bc8f236c21552d861034ae755b53377ec832863b35f43acfa2aa80e5bc868913b05555121bb8f8aa15ec1f65987ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12de1d02357f51945f0aa92ccf28abbdd4de6739ce1bf14b9d36f73b2ef1b369d90595e0b2f1003a9b8d1c2abe63f98ac2febc4084e6641;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b494399e96fd22623c330eb545be3c76f4fdd9bce02231475e42705303718fcff8c87e38a32b79973ceb7eae37b57703aa616d48e6478;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f876071eb7ebf805fde4fb66a6099add157334de89c516b2af685af639761b685a69fa0942ff436c10a564fd034065f1d8b60d4cdab47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193b7712b30b4d43024a3deb7810bbba57459415d4eb05b2a2bdf73e085077f60b0be1ad64450ee16f59005d711473151d083b878c1a6bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9588bbf6d2234086be21c57c6eef7f08ed488be6181f06b2d284fe14830efae1cdf5ff28919b6c7736fc4904d0f43bcb5e74b4605cb33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4277ef6a54c765a61806640e23984dd45b18ad6d79792656c89189ce75383b06bfb64a0628b06940735fe4b328e1a7702d55ea69292536;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1e9618268ff4012306092e92aa811bf450f2020f7d4e0878fb15f0eed5357c34cc430ca84af8ebd800d3fed91d78c8eb14085c96d08c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18898a382c50a3f3e44ddbc410a23c4695a6322bd60bb51704daad662056c593f95880f44f6b7a87d1c9f2900c16d42e1e7a6c5f4e0e53b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb949605ac7ec6df2defe2eec7b6a1042ad4cae7018179b52da3a7271e3336f92d0c3c0ed81c417fe52d9763cd1ee1f6c699a73131c9666;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15399883785b122042e4870293ffd9f0bef42d4400bdc1738aea91d3065cbaba1362e5372c6b8ac1186e782161d24273a945773a6a45ec6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h769c62498c11e531ffe7af4787e04d32a2a978d48050cf415e0ebd54f280b316ee8f961d9a98cbb11829cc025cca25fb01c900833246c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd5978c03b66720ad9cc25afca194f06cacb8523951f4907764e3af0498e52fef786f93716decfa085f486c05b84837af39dc7f8a8459d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1add4473623c7818b0f207d83ad5fbab48aebf0728c50fd4309ee03a7ff12ebd85b6447c06b3ccb83ad3228e0ac152be7612803348ea7e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bb8a5cb3069e43970866e60d31259d596968803ec3f35f4990dc59ca8f77e51d9f89b40dde030e633b4a4433a371d2984aa9755cd9b4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a2866d0e84f9727915f238ee6dd90bae671d14404a74141745b245756469efb0b239458a3d42e74f9ec242d27551f4c4b8e334ac66c6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30844fbedfb84fc088921ed75d64596d65e0752c21fb779e9eb22de89c3b5538617e4b23a831aae0b1650fa301b21ae85a1fa427c5edd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cbe35a57010ac37b0f7be1accee2ed6ac83c0270d9ef2b42d285cda4177a688f1aeb647c988e71d5f65d48977fcce441e9dadb49a80c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13644d14ed49669e9f9e37a6762dc2629dd590c7769afe9ef22d091c2d44119b9ca980d6077b5e81613119009a2ac898ae3d8eb350f7c9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e241336bce3b1f5b944785604fc7469bf778a38cd37d93dff90347ac99b655f92d80e2edefd6df2190fef6392cbbcae0ba6cafc5ed00a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47e83e46063dc726b9abfd5f0597ee256ccd9ed2d3e41547f29fcfb10035ce735f99cdc402ccf25482b17a045b8133cf9580a85f9965e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d549b4239b45daf7a301588a4a441106a5c55f4744e4dd83cfe9dc338bba5a1a4172fa2513e75ed2efc508c1cd13743ffff9cdac20aa19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1989c0845571ccd38703780a9a672ec84c8205e8d670fea168f68395f22fcb4276e97e706311c131e1a47788b1d1757cc152e4e41fcac9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ab1ac42f035d9de080ce1840c0ee22cbdd4fdfec53766993af4f21acc31ca828a18c1bc64e8aacdd58a0f8e9761990bfb481274740fdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dd83434c2e91723cfb476f857151e926ee473b321a8f21fa5cd4d76952a4a87ace11392b0e66747b8792c2b4671d7b13daa08977c5fb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a3cfd716b3bde9950499829675a8c0479bdf0777ae1f73a13b0c73d8dbc1efbaafb6ce18c62234ce3f12d4b5d8f1829dafee9996f3846;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1320c2f046db014a12a35cbb36ea5207a55646b72a51a6867a5f8c12c23439ec926a2a5a403871700cc91ce52e4c6e3ced6714491b861cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9ef6d50b8d8d0d1a545661bdfee7f454e6c57ee9d67c7d8777abbda55513387b4c593ccb5ffef10bdbbb79fa626a68e2fe774a48400aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174cfaaac0fa98711a35b17682332c75d504f5481d80acf8e2d36026ced67f548d649941c6c84ab961c9f144943b764890c09b3e0a168e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba7fddb4a3fddd2840ff9e5d2a4ad02b4fc5f33b9b7bbb3ea4d42c5e860983896ab6153b297d81e67acd2d9aa6d1e61df76bd6e26973a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23c15f0ceb2403ce72a5f752009246e32cb5d911a6ea9dcb12371f74d754e4b50be417d658aed418b724abde39895fd646d8ee996371af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdc416f069a2e83371f4443b65a2f7afecc1058d636b0d81e4cf6958f2ec99f3242551bcd737cc645e472fb03f0086c9a2577756ca3132;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h684000ec034771157374d388beea3664827c2fbc0be685f9870748de8616081497ca581db2f5d838c377db74e88f62e63814f9ae3c7ee7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3e0f32115cc5ea844a5aec914c9efb7a2d6de62a3a27f95b5dbad6d8803a06cb1018b37f6917f2d00786ac9bda36db5cf5f361698063c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c7f9ccb10be6b9896f5d6fb390b062a1b3479dab4a092eef20f81e8a13c3bf2c2a3568c9f18ed15741bef7b293c921989a1ab046792aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1812dc9fd0b074b721a38e8a11f56e607ed357f28b75c45f4a719a3f10400d2e64a1435bf31c05342aa8d15313aca432d699edfd3abfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3bdbd6c059d8076ff30eb52fb8866536efaa57d8bf5cb6d067ad762cce18bfc88a7455c986384247926b833a78a869daddd1fe42a5408;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ac2d9dce8bd8dff0b7ae338741f6d621d5b221cab65875cad2f0573f9e61eddcc4b96fb88b43721f5e1b7dadbefb6e296175c87d9f4cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e81c6535b1b8c2355734b0de1b39cec7cc701a66ad4e8b538d5e2194215e465070bbc915a8c57773daf9a42a9006b4df07a57f0be82b6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16063ede2a3168b2389432af5f169ad1a410e2aa99fc4e2f5c57e2da82cad52865875e2cb732ef89768232a2a700757746cc69e7c4b8902;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd45bb9bfd187f423ede9b4acece086d5376de316936bc2365ec78fa77cc48582282074e880b087b4cf6273e8bab38c156d5c395b3aefb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf061bfc796a44acee0b97c7479f17aff145a02a863fc3b9e37d25f33306496ed7e91abd301d057bb0cf57cb4a8cc57db27dd6f569d9aa3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1036e2ae413cb6fd0e0bd1645461940f0dadf3ca0d81c98d08bc6cdc1ca0136efed6eda97b1a0ccd8e81718e040aa43d3603d7225f0a3bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ddec256a4699e0a35dfef5fe23e2418e973c418c5c7bb062a0216cb8c889d62e248acd1e234dfa85da361ae56652e9262f06dfaa3bdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147e95c8f3c4e23d2eabe7b30f698267902ba8f6d6dd5fd414404a1c5536ad6ae0e65dda531c11cfa38ebdc32b788f49dc1f9fcbe1cd048;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121fc7e8a3e5829e5d2738992ae0bae9a0b00041b6897a952e5d9b2717ea5d9b51d11a2a601da09518b231e5acc911a2b2cbe23c9812144;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4aa1ef08ab74b692fe1e087de1d5475ccc7358d04a08779d160733ec06d40d7fffe349cd0c5d7aeff6d2690a16d64a56292cd21c1c1f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f9ee709da1b1b7983e9cc916b714d03f7a6673d6b72cc57b6d77504e352698887b3af49ea85101d86f225cfd75f900c19ed7ac0ac016b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ed5a53d9a78ab54adbfd2cd9c66ec4bc0e2eeea626a828762433989a067fc63663d3caacef1fedcde07630b8d7c313e8310cccc158822;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128f2b395a8d5ed6896b214d365f82f25955c18627b563977a960093c9cd8470ff752dbbc62764bac3003e59a6a4da4443a5893310242a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h365c2441a7570f34a3390a7ce9204b4d43ba402064879c7cbd71ecf9db63a6283cbe757320b90a888fd417160ab09bc545a69d46410a8c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0e4c4b21de5c384dd5270d96399ca65f9ea45767bc356a05b81c3e507bd6bf87642853e0c4da65749a6e70439216c14bc0d334e8beee1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd88c82d1699e01a5b6a9aa53a22f42f81e86ddaf75761780d419d3badf56fd8d413df165e6812a195b2ef8da7102f67785ff9bb9889900;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123b99e8c81e14e565c0945d07dd7807ae06390ecf11da5f30ddd2b4b500398e50ff477b55e8bb8a3b7b29fb050cf1fbd79710ed6cc0125;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8477138eee1d8a93ae6b5eedd7cbb01e9cd4407e453ab48837b8e9b6d24af0af5261dd12dbd1e899eeddb1f22d7f7e0324e4b620330f99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34cd9bb2c0ffd927d0b3fa9666cc1bed5647baa8f18ec1faba0a8c6cf3b107de279b501884006695b9db112c20d38403a309e97d42fac9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177435117c88597bdc608f6fcd46bb52aada9863971c4b235c405148f9622e050a443a77e0f13e3ae9b93340595e7d6f63c6d910224a8d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d678abf6fb361fbc9a95048df9534e92ee6cceb039cf5a0baa708689dce2ba8ffbd6866fa89398ac9cfb7a33438290252003a6fe79f85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ca4ed50f70c18fcb1feb6a1a162221fe34da0bd8e94991e7c6b7edbd62ce0300dc8f6febc3023d780626e01418a31a8441bd82d099449;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11beaa9bcf854fc4926f4c7b17e8ab6de9d5bf0c59405cf9258b12c1101f5910ed8a1cbc9371e77ad992d8a29ad675137329367ae85275b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eaefcf2188db5171432a79f14b1e44878fc2761e2b6e3c53d931e373b06b471fe94982f89a82d452db4c3ee13a701f952666de47815718;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ab2505dad33e6577dd7364e96b45fcb1657ef35a9b81f47e7ede9f1ad09ecadcd433e92eafd2e3b0410f1b4dc07b99e77bc21718a8acf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f37c85b32ebff9bbfc62113b2021ba0d2c58ac9c487652ee137c840edc0afec11f7dcc840a2de267900c35b01317255b8aa434f1135977;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h774010753c9738fbfe15b8996f208d584b7dfce19cd2d2069ba4625031f9e92ea9753ad69ae746c03ea2528dd6187e45da25240c078c66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ddd779ac2619d56f7c5ad5d6ce3a06c91c9476899de27788ab588cdd9ccd1c2a2e1ed589516792b972c1100d2bcf0113b5f9aca5cf87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11251cabea4e5592604471e5aaf4f48efa6c2611e8798251daebe95711110d496a342f5b845f2f4211986bee456857de27b84bd97dd48a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f639b62391695008de538966fc63cf3b7302672faf00ef1100c70c6ebacfbe25f6cd9931cd8dba8e868f4336a04b6bb5cdd6eca75f6f5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h307828346e7fcb4cd02898f19c86d88f5d7982ee7931fa86f42b037f4af798b7835f905d48e0e65707ad5fd1a2a710abb67586ab89e660;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6b198affbdc2f5bc1a58fa863b172fa43597950d87eed2839db50b22abb9f183798d03657314b27a363e2d33d7f08ce5c13f4e06c841d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdfdcd87ffdbd9d0e360da458f947b4c4b5d144268f7ca60b27b3f1451f7eb04e21b235f119b4d13d502017584d4ff1bb8e98e0ea17d27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf53cf5dc7cb6300761e380641cd41f1687f7b2206f7442511710e8733ff316bb0764d855cff1557bb0e862f3638284394970aaf58a04b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e41f915d004f2cab1cc6fbab7237ece60a3834f13f5bd135d6cc052978a7701d2901b524085d0cc102a9b6ca427054f26a4a8276c01ad4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1256a9299ca4ebc217f8b53eb19d20246424facdea131deb435039f6c1728c7777d784e3b66b85fb89bf78d5c07db887b09c866fd9cb2f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c283531a742fe17be113988d254c8e2f37cc28e017a5d606a37bdf2f863f46af796eb482dc897f2a1b842d5bb32bae3f33a8fd1f5b3dd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1974dfbe112c59865c98c5117ff7e8db257507db047d84b2a0f2323ff5a75dd9f68ecb6157aee440a31076aaf0821c97a1cb03b3396e54f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2dc2e827b320481bbcb9a68e301e79bd46fc5e45e5041d0cc9442cf099c208dff6ecd81bde76f86e88defa49a4ee3bcffafab504e1bb4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc548e4d51bd717c0d04e90ce227ec72807015b091d6067a40d55385ab436d5499eaebbcc9cbea087d23bae3f4a39656634f6fba919524a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf90765f8f1b5977b3db86bafc18022ac55a8f98a480bcbcb61b02031855849af020de812e237445ea73722d184d7919773646a114fd6cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156a88cf5fa19f8ce88a6382356069b4e0aea8d6229d1d2fd53f72ba1886a2457ffb223e4a437e1baaa977d96573f9fb5d647ed1650e410;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c70a90408717d5aed89d48940588a86dacbacf5ed61e7fd9d00cdc3f7f1320a0cb1f31193cba7ce98eee6597c69dd77ad2d7e6bc17ce1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7a4ed96319cdb64e06b804791fbff891fea2597831a98f3cc888c8ecc8170c7ba3f4c14ff1494de1447bcf35099b4261829440187e53a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11745061de57e2d025bf90ecc99737bc3cc6ec29bc7c312fac84237ecf1f2378bfe1f6065a01485600152ebe30178bda27fceb9189998e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc03b488cf94396c3b149ee2f207c32e0c8c580562d10773437495d8a6d8304c07901ee83d988355a258387fb7207b38a3e66a5fbf40ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cff9860be040cb4bbab94f3e039ef24893400a3e99cc7134d749c89e58fc77102e6830ed1ddfcf928e71654fe8660b63fd9488e5af8a17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77ac837bb70816e71d3515a58890a5b5a83f80a3dbbe8ae875397f76a397e90cdd5fd444fab7980bf71f5a9c4f66bfc47633d1b5a8480d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a11a23e4648f87457893d89a84c64fe54f04914c6a30b76d0b8555e82748a14641b4f1d6d6155a54a77e35212663604d324a9bd77f64c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77ac40b8770ceb9d7c37603ef322ab448bfaf89f0d901430d1fd68ffb53e62964a98260505a2b06742b1d10396eb0d8cd657fa3ad4c23f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1266e44ba0f6756c7283aa35102f12b22198e085109657d064c757bdc11bfef5178d4ab15371fb9ce1d5d5a36616b94c941ba2100c7829;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f1734410f98ffa52987b382d7283c25dcc604fa799570c060cd178dfdfa6df62c0f754c675ac440a1c2eef2e7217f33d2e992fec93bbc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca14b96793ea4cbd47121c067f889fa3fd8ab63b44b284f20be93e52dc0d3b362ed6e573ff8b6736645d685f06cfe0b4d5ba928352926b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14729d0a590ea06b87ddde1702252e3f10bd6dc3210216988cc8de1daaec2d1435752fde5a7ae55aecbf5c7074046b4c3c1a535eadd9743;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc30c761e2e9b6da49462ed264e8bb8068e4e179e7a171e22b1e87b022e667079b7a4cd15127b7c728a2b8ecbc7c97ecd331e1642012381;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e84d79236085768b0246d36250e1aa139ee1fd3d6dd6cc019525b1d7814489b5adddba11f65fa0f04d2710aaf825f0ff48a70e3c1a0a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e465d530dff0745e088a1ce9f8df26b9b47a79143ad099a5171ff9a7cf34001cce286bd0e83b629f447a0849c7be88e3c2afd3b3600a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he05ba6a5f66319cfbb457b5d99238c9dfe7ec8452b5e42fc4151f3860da90b0f2e80798b5b03ccd11c164bdc462979138b8fcf46f5acda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93ad251bca4bf05d1f4044cc0c1fd86da4da2c6e82da77cd0be524e736cac421f549a342a3c401641978c1554299597fb0e798f7cbd156;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc57d1062dad3801575df630d57f09c13c2a34faeb6334317f046ccfe7f35cdfb04ff30ee0c1e7761cf4f59c2bfe954cb68fb95e5590c68;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f3a533cafa45376fe092cbcb86a430d355561eef56ef87d970cd950ed309d33603956880088d63b2593dab23418290928bce067d0a6c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6678c1cb3727a2a046d9b4cea77cd61bc1f4879e052d4261c3eda8125bd0b276d81521d847c288290b6459285ebf66d649e32920955189;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9fce04dde904bb370e1889a8654b8eef3708bc0eccc10ca72c54cf73014c4b5b13f6a4e38897717bf60918405138b45bad01db4c18243c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e2df3c54bbdfb381be9144f2e84ffb1ca1824ac3fd7979fc9cd3c1d43e250f73c7a4059ca0a4f190930659283e0d725e1fec4087149b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5673e5ed58e2a5dc7cd4acd8f6bccb06a7c4a287fa62dd4edbe59548c26cee3ef13ff5184881455ea4f758b505b1c86a9bb40ed58a524;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b4f205c6da098f214282a695b3e9bb726f1e98517d5fd6a54a96b7603730de352a7c2d4deb7d6862f7761efe552230e3f399fb529b584;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b363ae3a0f34993fa071de5c13d3bc72416c6d3abf296619297be8d8d1241d6d880a1a978a9e1f3274e8af4dc4bd0dc6c709f3a59b6fff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa8079d97124719ed2d9256c2f0d943b10bdb6209f17446ef88f52dda9fe135d440e383c9e78aa11a9aa4276327010a3294278897ce11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164b5475a62fa9be1adb135ef5f4d83e7aa079264cbdf66322f387ae2dc0d2bfd9c9e8ec4786656268aa2d0200b09a99e6c125d3e543ebe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h484b5ef55a084c6295a6f13cf09680dc509f17b6ebfd58e866541a9207a90cab941e835bec40ce745276a2f399299813f7ca8fb4c61ac8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5abaa9d30f2675ba912453fba17aec2e890ca3a7003559b09afd6a98b6c706e76686c47055b9cc5100fb10e6a5eb083de0196055abe8b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf67d7faba73934092dc97c4181be8fb63bb7ee92e1e6b746141264ff1ea66a359553d5f8dbadd3e18412b66cdd717fedac0d82b8991bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha198ae9030fb732b6bfab3d97ec200e3d4bedd0e742028deb251926432c6a2cfae1c62480517727ac9bba0ddbb3fccaae83a0cb7e2167f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7090ea553efdf3f6f9cad6d478bb7eb7994c3f009a1d3d454ea757662687c39fb50074f3f3cf02c6015a6ac445971c5c69b47e12d583a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e8041ea6cacf54939b83f89adfec0be9030790385ef776535313caa7c92e8fc67ca9156db3aa9018ba53530611031b475104a11e3cf2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h497128058282d5644d52aeddbaaf7bdd953c89346333b9bbfa6ebca4b084ac074df3175b92eb99a2daabd4fe40a560feee13c02a744604;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb8fd75998835735ae365d8e4b39913380e0b11380f6722186a6c9ec6514f473940cc18cd3e94b5f7a9a296d61e1b7b821096b13d5f585;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac903ca3f35324cd863bd73511bda4aea6406ff14717c789b7f2b0b6dbdf58ed4374c9d90e312956dcf2011eede0e5fdd7a3f700380c3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had6ac734cc8ae51f5125b565caea5373a1a03f344fc7c232342d62d0b42d1938c9f977b587b4a53c6270833fa951af2df31ed3190579b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140136a31bf71d96bd83f9292ee68833c50e1ba4a27c3b43213d380125a703c69485014b42ccac90e7972a9dee9469c9b8751f2def1ee3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab48890d435017eab5fb0c0ec784aca0b6448e5dd68c8f90fc2b5772987ab2c5db05e6c7889f5eb0c1600b09d19a7810227bf8adc04872;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ceb1d1f9d7df4806b442b306934ca9e3d65ea57ba6ae0969ac35bf595b3bf027314fd2016bc3bacda9ca35902f3400da4e93dd31f361d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e12985a21e996553ac410bcdfceece3601dbccbed70f725a7b84b16b321aecfd41d2047cf9f8f3f727063e8526158de31ed4482d6956f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ddb9021b3ba563c740340ffd02d6bf5c95305a63b7070075b1e2c1b1ac95ceecf20b73ed4b987ff2fe01c04dfed8e99f97e29d6ac4f81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19442bc82c4ed868d8e20bef930504f153900463dc93a63df7a6bd8147a5e38f2272d7ef702d389f3bcdb7c24985fef549a090c75ae3d32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a005217e6751d44e9b37862436cf54065aa67fb737f5cb89f0313d7c4dafe1277a9294c8e1d3dfa0fe37d97c054a9735e4c3fd91dfccc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b35968743c4d837a15d90bac28d82368254fc97f224293ed2ae747356bbfb9efe1d1a0c1a9b8816ed5715c80cc2b0eca941d12ebb499c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7eaacea5215f579508dfbe48d624125d7816d61689acba1bf70c8f7927cba32eda41ab39febc3b250160b6168b2b5323fcfc32f14c8410;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b38dfbc7c750a174003f0863e40fb6a0a97f7c5574259b735524bbeb914663dba2540d9a04033aaf36be89294edfa388ac9c7afa5742b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c84f29872a5843c7dfb24aeaf6fbaebcf37ae40c323263b7b591198857340950adbb4f4b5c88470fa4a57492ba75d29ae77673be8eb466;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had7a43d3c54081c528eaae7767bb4f985bcbb798533d311c2f01b503667b154e4d7f4b905a18919d6a0c65380f2a3a9a6d564778bd01fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha042bd1060df89e03312e98145c2d1887929e1cbf72d83fc00fb8ddaf9281283d69b9877a1d8c3d8cc58f6fb4edf6c3aa264c184dd0e88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f4d66bde435fb68ca1758574f7a3ec8489a7b03db488678485eedae778de0a152654b20d54f8ba42dcd62bb98cc9853c3782b412d7eac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd4a20d22925bda4c472da837ccc89e4552bd26378d08a5fc5d0078c74dbe08ae50ca5d911a05e7df8ccd48865dd634ae1409f282c716f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5b6561b7738ca9f4f7ff3d574411e1c1a1a8e0ee54803099550c59156a9dd3717542e8bb0b6420b7a65b9bfd7a3a41d51c96687f06e1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178c338641aefe5f0ec6a183af2e4a5419e720bc1b3686d7bd38199928b2c87149eef68afbf79500cb32df373eae8e8972fe41e20c40c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h328111a0dc655c3a313cdcc7d2078671cedd70a96f1d9c57150c10c5429a8c12404d5fd4623d435bace1679cd42fb60603a9c0e02b1c98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d6ef8a87211e01bd2af8af60a9dfbb601cc06797883f804e03de88ada2cd8090e34de3340b865da8106bf81cc82a437ae708401ac4ad4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1994861fcec896f0c756947679ebb489dc3420a960bb16e0c57b2dfba26b0bd612990c5d402f4950f8f560ffc5c9ba02f471a8bd09fd8b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbf2992f580e1d8784825f2709a889c9b2d9624ede0233b3c763f6ca31caef794abf19876994a02982cefad73a60a0ed62b0e8bdd9583c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6ec9896cd78ccb1e2d23e9ddec8c30c0a1a58a89f02173484e7dcb4473d04baeedf9049ff311575b5a563d6b96e989447f7dac93104c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h805372e0288dbd762c78ab9ab9bdb7083ad1a4e861c28df78e5c8073843df10f7e313b45d0e5e60a3c072c083a50f9646400d2664e53ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185910285fe22691244f06b0b43d9e2b7148b20b789f2c734ce59ba617a1c791de561ca4458dd6989b9242bf75b3fbd5075a5d1641a7a52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b978dfdd720d776ad8c2f28d32a8bcbe4c3d7d605b10e2a07b042bfeaa2b8e8eb53198197d5a315ab1d08b0493aea57139d15a40a881f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacd93d049e5d81add92b684c03042d5b5c243bacd6e97b3c804d40f206c717c2370c76148b63d51223fa552bbd1dfe349b880ebc7dac41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1f704654f1ffe5fa872144061b80055f06a1d700e9088d79378dea954f80b592b84a251d1f512819e678f185844d95f50193470ce1e71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129c3cc14774f316650656ec7df45be9ad7f0d6666d11cf1fe79431054d7aca3d6c0a60a141578bacfd6cbd6d98af28f9ddce056319e45f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128144f4346c9e8c6a7240668094969143b80de7996086e2b1897fda9f94a346098ab65ed253ab4ab7d80c4590d6dad4532a11d92ef61a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c494012062a51943acd5cd937d8aac74898d86ef3021626e5ee8d3acd7dbab006ee3ca65da188dabda8f25e81deda798f2fe4033de1640;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17806c4098630ccbc34cb018f3a3dc3a6c8051bc5205b41928d79d344f0882ced5ce32e70b579d8ff0f1a7fb8f1adf10e0be411296c53f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7c93ec8a53d2cbd2ff9c0a728ff29d74cbfa73d1d27ecdd6b3c883ba8e12dd7c3a7f2831294dea1a7f1c5f85eb8264582fff800ee05bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e37ee53adb001ccd13f2504295c57bcbfb8063d20911ecaf92fb39e8527c7529b2a3fa9b6f63ee5d76b6b3487bb0b125a29b523191783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b902e65e358ec14215f3fceb7eddbf5b594addccb043e34c7f69d26a52b8181c4057a8819e2df7ec7ffbca5bfd5ee0ae5e627b01fc4ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1214c1a7fa8ef5baa423a3097856c490b62216a5e4d616eb2e0b082677a30f4be081199c002b3cd75942224c1a94370e90387825025f7e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h296bb9b69e78259f03b39ed64bfdd66b418e331a112bc0cc683f0430aa625740950b48697f775a7a6ed6f003dc4d5ebd3bed629464c792;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7514241d2f5f7e548c6585516298ea6d7ddaaf85accaeb3a44e92cbc15936155e4cc0cc8ddb6e583c56e1fe70ce7ca8f11fc5130eea17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d33f58d5915bab5b39b1fbcb4ed30b272b31e40bba32d0ff0f4b8ba6f906deecef8055bcfa16244b47edeea2226c96fa3a983ae96e260;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70c6ca86ec703d4b65f4988571b90d4e6eb20b8ada544ae2943390269f55e96f3503634b6f54e5866a20a470b0a82019def3ef7ed90796;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84e20049861d9ab0b4e30249d58e5cdd9fb6b2856d62d95d088f75c711d308425b215ccfbaee9038b994c1e87891049337c776c67c6e8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d029381ecb0f5e2a2723b4f3327294cc6d47b26b9788f1d0affd11283ebd7feddd232bc112813b22caa087d93608ff2a16120d1f07cda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13240329e5430cbe9f2c4d45f747ea396464ea5f5e33bede9ea0a251eec3fffa0e8a83d9e88a7990e19c995f59fbb1c4ddc44ea4c783acc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a376e1c7a02e8b759ed2803bd22fe9a0062f5251c4fc70457b4ca53b4c0fb8a15b88c6e5784ac7a1994d799d8145f2b4a9ba971cf45f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9edc7add53bbd490c45a577759d3a0a2173b2d09b336cd01835ac388e2502f085c3d2b5396c44981d1fc8d11080be8302d9f6579b2b29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42094237c777df1c1b9efceab13ebce1b2c75d0ed96bbde4952b9e890aefd038deaf06505c43a4c87b8497e6425143408b946df3402b4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab6ffc98ace53b4e17ae3fc49dada044d08ae90fef8f16ca8996d1f60c138e41ce90f78187c781f038893184bc5a0bb8993ebbd609ee9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce490d6c4a31b803d82821c960ef9af26aa2cc7090275e01256303995920bc080ce05bf66dc6a432724e648e6f73aec904f507a0618d62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b66963bfbba83f55b0da08cdaa3e23e58ce8a13a10d40dcea00db8306eb8358ca5e86d70b815d3ae484a7ff4fcf36c4eb020c531c1c8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169c75dace2d74f09571e517c994e1679b24785f1c424f62e4973f7721c44e136ec73a96b2bfa17ad311a4b3b1ca0dbb6a206f01e7e0657;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d89e1027acf5aff3f031684ef3da58a89cbe08f1d4d5688425912dfdb820ae35f4af14fb879e39169b791651095034223c83a3c3a177d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcd5f0ca0e4307e16eb3488300fdaf289a343a6fb044ea6864bfee41ac16555b7052e357783cc7b9e5d23bbff5c779c58426881ec86375;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9bf1abb5c0fccea4b31808777ecb02988e8b45de02da161da8c024033e60a3b686e6194bc0e6e51b45dad7ec41b6ac0a3b3416666ace;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29172ffa7609a5abc479479fe270d1e7a69e05a8c823d2a4d200a27bc570cb9904c3306a01426a2b1e6c740c9e8ab6bb91e92afebcb1b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8bfbf15e5b72bf3157ff20d0b3bddf8dfa8725b2ce0baa80321a6c5b861ea71339de474e21a633577131070df8f7c25e93c1ae6fa4a1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54f4b143bb45e9e495421502e08faf5144da9e2e881e68ac01aee2d87748af1c130cb74ccbb52c6d874efc7d2031989eaaa98abddaefec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6bb88ae7b4c6bc5586005f8debec03de1e50259742ff8d6b3e108ee4197f8c914e5776348dffb356e5c23d009b3435cf6fc393d702f42;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb09ca57903e5f15c13c685b6c6c951a054b972b1164a49e6959348d1fae1e261ce13137f46cab93fb0c9a018ba0ef1dcd55bdb571f055;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc3322536def5f591044abb961c7ae13041b7fd0d3b5ac55958d1bb110cb2a0382ade88d49121892dcaa34a050ea4f30f1bf135576ca63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21be36c50ea3a68dbb6e4e234d20424f984bdecbf9cfb93e84abd5d8be7fb5bf9667ce6e5248b03c5d87f2317e08182780f986134469b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58b5957313ba16e04cd2fd3e156ce0c322b086bbf357738382c98a0bd20c069a385ad15b22bd555262a4ef9376637e83665be81ca21381;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76ec02b2575dd0aa7d7bf3f4b415b1cc671ac697b62ed98bc64c01e6fbb84bf4d61f1bc0931994c4cfd1b73f29a27817679c73b48bc1ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8121cf4b023a03ddf345958f14b24de95f55982381faa8fb54008754987eb9840327e66a973c79eff9b5f0f1815d77e520322e337cfe7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb30cdbee7b92c6bfd899606c9351cc468de2de4ed1eeb5103ec8ea61992ddc3febc25957f1427a82724d99848f9d05cf72cd6640f73b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e796fd6ac685cc77968df2de769563c241ebb5e15662e6ff66161d9150c60001e02fcff7f5fa187996de8c7fddfc0b25682e42445c342;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c7a33a3920a039e073cf8a21473522bc56ef6e2471c12697a80755a9dd906ef3821dd8e187f51cffd3a3826ccbdbbca66e042699c098b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f2bb12ca3ed2e295c82b77a93cb7f282863bb1db6847f1ad92964da3e3868f63b69e104d369fc8f3544c2b7d095ca7d76abad55eed80b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h570f29233581d6b158c0c1cbcef26e8873c627f26de9b1693f23887efff564a69f98fa970393a7c6584b13e04ee99277e81e688f11a21c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0e0ae89951b9eb9566a86ace64e84121267aa51d2e798d38fd2e76cc0a70bf1d951f6efb83f486074f64f32147db04f1f727047dc3976;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106c21c041f1635f34c22477c2e16f9a63250a6a19732eca7af6c82ba2f1d7e7f973127842a00dabd95e2cbafd3dcd2c3cdf155ee9b5b69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134dcba5ea2b965ddba6b43425ab350748229601136cae95dcabd0a8369f100af8eee051285d9f4edeebccce869aee7749668d207af5619;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba000cae384fcfd28bb388c9724da647b23028d0ab045dc4725bb00bc13a204d8d634b244b04d2e2f820dc5a3eafaa0a1139b28b9b1b0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5fb4cd947240763bef6f5cd98719ccccd3581739eaa2ca51c701317d35521336146142937361cfa73a7780e3f177d95ece086ed71845e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a27fd9a7c81b9bbe7059b10d62bbc4eb2fef6ba9ffa10f16a66ce724dc094641999a5ec72a8a8ad6738eb374fabc50cde7ff140cd1164;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c78f563767c3a560b26520936aad77c23d0f43c1f55bf3dce1baaf6ffd4f76af83786ae4901e988340e573eadf44a019f78aad22472a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f23e3bb0aafb73583f838f748098fbd56beb31103d44942cc9e2f44102083dee7968d76629d66199ec5bb6c0da5e71b484a713144f8961;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1edb3cf9786f0303e0248c3d7dafdad5ee15a55f9d7a1269b7d8ef44ed07a6dade63ec5cdf81f08e71890b1aa4100860378f6d8cad2fb01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9885e19abc588ea2cdb376497c058b5295269076fcf1e6fbb076a94f96baec3c2c667d8f20db207ba58d3ba261c3d4594ba16a337ab0c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b612f701887b630487c23eafe4a0e43f726c34487265adee2effe6e6e284a4e4bec769bf346d8a48a7c48eb9af331535168d58beae0cf8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130ca924be1b3ee9fc6bc3a48e50dc42478839707dea3764caef128fc94288875034e467f5d19055dd1c836404db0878c4e6876d202905f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135e9192c5ec591217e7587122b5db0a86cbbb9f26879fe2aa9cf268d6a502d03ea8a0dc25d61b10f37a33dff3957dc730a45d084f8d78c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e4fbb57fb05182c232125c110ae175238097b887ff839607577fa353ef59c8675a8fd10f55611feb9c6ffcf4e353ef75c9e7398e62ea6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae16831dd48c61eefbe8e8ea4a511d511933dd7daa148cd5feae8c05cd1564c121b29e46f176e306a6b0b6f55a384d828d6fbee69f2762;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cf68d314f3b9e6e65b0182bb1c28d858f13e04d4f1870c8b834abebb48a5601e8fa2ba8f3fb19856808705aa40ac0ed239a7301a9c6db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc9c295d4639c637ecc420fa4623842d0982a8851011b0613ea9e418d866995e7e3ddd3a38aac4682837fa28b4f409614a707d4c76be99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1138f50467e72061a3272554aa4f03b9507219be988be0246273093d48dae94df2aec59477e6eb3428d0361d218ade2e157e8a95b4a4284;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2940405191adfe64f8d6cad120d374a554b758c2c6a05c2ad1e60e144973f9e482669ff9e598be4736783e8b260d871e6534796e1641e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63a51cf96bf648d4df9f64cb5e2410f1754c68f2c84968675e506fcca845a4ecee3338aea5f992124e4e6a4066e601514f3e41bfeb6c37;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6910a30852cf120183e08dcb9efafe793c0c944d5dafce600363a9229ae4e39b6f9da5d493b9c5aefa07ac99d04b4689e46b91e6009c63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h818649d1737ab9982d904bfb7aae0f66e61cac376196d5768060900a847f70c1e53c7dd082dd46726b3d6e660675961361f16fece429e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc51076365151e82b97b7595347001fa9a8e3449714de2e56db93574ad1b85787a0352eb6ea69dc441dc52861cb397016d55dbff1cec085;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2615969dcb8751f7fce3e92ca36fa0a909c5a0dd0eb5e50e5002617c697326150a5d141d6376fe1044314275505c5212feabc3e56df2f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cb015960d90b901630d60198af29ca71da2d8cfc801df2027254f4882602b54e36d7e302ca603f25933a2aa3113b3e40bf1e6a6a171f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa318c52a49ca8c719604578e6f8632aa5c3fa49dcec467b38c5a91f244c067465b50d43929ff5bcb11560987a4a57bdab71cacae5dc87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h435509ac75e15e50904f0c68d91e5635512cf219f713d8ebd748c507c745938357fd176f2bee5bd99b5d3b90569a05df56200c79910f3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4f65c028dbda1b4f1f9185391ed7835ea5cd166da4a84a26d6c0f22f63807f0831d40284a541e69098f59d4829d0be55405c57ead94f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f41d16aad473d3f660bb2a2adcf8b0f4adc890668f2cc980e6728c1c536a8d30f4b6d0fa02abc3cf941340cb09cae6cf6e9738848a153;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7c4885e9ae5262b3a9aa89e363d6f072cb97dc4cae3edf247940a870656c4710af35eb4b7a55eff893f57337acdf89d923dcaa2de4e1b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebe873b4d00ff5d192287ff2f44e90e787e20d24c8bee05185f50057dc825458f2a7e12addeb5d9bad89bec98c3f18a0d546f891adc0ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14afb372a20d4846561f0f40143ee3bbc52c7d996ef12a3725e25393361df75ba2762e5022f2ceb4ac8ebae4e394901dcec2d9919d0a37e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19de62522d87fcb775aa94c33e38777feabcbffbca2258ab5cc2af7b747cb2532817afc35a630a2b5e402358f5c1684e0ef86804adfbcdd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0a511f8d6322172585cdaa74ab5c1040e7d32560696a07a38fdd7b278e61d9aeb551c6293d3844417234b60702fb8d4ca9e80f4dfa426;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4fa108a4262e078356e068fd02f7b539ca7745a604355b1401dff0b2aafa039ee903b52d3186314ebbf6a107c0c5c4b3f8f84bb2d0c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5dd37fddcda76dfb3b554189479bc253ce64557dac1237ae88522dfcf8903334c6b79107f40d40898617b13e0bf5a3c25f0ae79acf6d8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3125c4b162ba185c73b5af5508e9e8022451055cbeaa60efa8c99eac3276a723ec32956e098626e17d9684b5af6cb8f0f2b229eff5e058;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ab6ab3370635a37793b414ffcd18b21212044e39d763e501a5ad1bc742999e11ffb3257fe0a7946dadbca46ebf68d869dd8e0267f888a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc3cd511702a8f3dc1ecb28e9f5bb017dda96b2366e6fe517b18e5baed45ed5c2630c69f1a1a3b9de59aa66e62d529564c12d2d121c7d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ec0457cce51c837ec701d73bab2587d4f96bf0d5ef009ab926eff35b10ce640d7888d5a5269ab9789f46f4ef769aaadcf6f9baa02de72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dec1af041da587e510af18797fa2ff13c29da1430659a30aa48d604868f787ab05d908207e08e3b0717d1da86d8becf6a47cbe99035651;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1737ad35ef41c6637fec9f0e26a41e9d0d416a97d4efc09cc4f76c089b1fd9a7152a367b9a2f2db4f679ff423128cd5dc9e8d2cfc016b61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1f5c67594f5932b37da205732fb0c7e7531738cb15feb888fd27292d0f5da2bfd1f55d0a2c8fc5e8d54c931a318fb7de5e1eed4530233;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h534394e2887d1fcf619970aba7976595c570bb7570bf5f73744ffb706975e1c73b35f7797a1b6c28efaa3a30af921e254f54c26fc6e640;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a21ebca8e551c929577475d27d7fe0508b566c3d29491094964a9940d1fd4ceadf386153e712c0fc2b43c9a7316c2bb0a61bf59edce9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e789a30f1aa37919e6e0957bdc562f133dc8f8b1bfd0b217cab394ef143eeaa6cf58d46af61ce602e3a80e98ad8582dd0e271c1b152ada;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1050896167979195ce85bb232ba61eaac804cd4e9d95da146789dd7173e4c293869a8e3c305d2d13a812cadea21c747c789393d41d9dbba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4be73b2905e3284e9de36f15b3879c5feeb2ebf3a20e812414ebcaa63b971b07d6e4f7e0c94abf32a290c087ebd4eac6daa78b959747c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9be2078d0b72a3d3b8538a23c3fc3decd3a27cef062709b3569d404d99210448a2b3775469e4d0cff80c9638c47bacc25df8b6761e8d11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1054cdaf6cd92a4cd221f1c1445413e9e2cc54a4488354040cfb23173cff530f118abdb2d21306e5af2bfeb2422ca69a93b3e9e65030856;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1632326e131d3b15f2914fc2dc8c7b61021da2df2241aae3218462b23295eaf61a4b4ed480eb16bfa7f5afc0b026f32812ad2f371ae4578;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1910bea620bcfc8059f0891cb2e289a8755db474671f29d62cc91de4ef86379acf9b3a4a6998682c3b2323ad784a2e8c9bc76e38eb282f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16679f622ae8586d4561f639a95d769fbf92d78866a8385cc72208438f83625968af2db3d0c93568262f7a27f0e7dd2e79e44e11398e9b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8c2d727f83eb72626868beeade2865aedf207b2dcd4b08ef7c19d975b9c1ba51131a2eb2a620ae7c10f5310321d47c5e25c02fad6cd49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he272b460d5d1ef3e77f3266d81d18f23cc2f7c01d875127380314552fbfc46f9b0c2f9f7f36411ba3132a5656983d5447ba2b9846ab8d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd711a3fb264ba5f9180aea33972aeaafaf906db443e6d8ea0bd678583a11f6c8c4c25b6d618e476eba1690cebc5ff9f10fbb0f4f7e9f2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b52064e6498b027afa8a94ac034d7cb91f9e2db6dd5659747545dcf849ec0d006a02cf2facce309f48a884dbc070b4083bc2fa46af2f22;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdee464e5c14a56d3efea6d4632fdfc89aa03b6b9e635e1c3e40511c03deb4c4dc5f6ceb8a493ae826fad1ce552e84337f738ecd55ce71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77b3c8bae58c96072a2d7bff14a77e6b531e280fdbae2a78d2e58d8467b84607188acb0ab04373e8a6c2fa57005cb1b8bcab8b02a10776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3eab1ca69b0f357f133acda6a793b729db7fefdccd7a3e145e0ab2974076967fd1cd75b98dbbaa8ca7058755dc251ad9f36cbcfadd73b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133017dc0f7fd5fa678fe5d11bc81377a435ff20f29a367bc32f2370aac700caf0964a105b2f982481e9fcdf43d3e64bc635b53a8c4d3c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd64d87eca204ae7da221e69f030c7670f64f06cb0a553ef14d02d5629ef7480b382775f94f359b1b7f59fb3a72153ffa4b3a4c956a32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb6e80235d0c04bf266adbc3c03d1b339bb1d0c836294458768da45e8b8eabc5f2abb0db1c3c0748d5b13bf4470d3ce1a5179d4651a613;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9732c244728236232c08108bc5643f2151c4c97660b67087bf9e22038e45f810a4ea592a86a8706a39b7b7ab0c2a6181baed8cbdbcf80a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ac8d83ccf43b9aa7f0a9c57d17427fb22db7ee3be9b3f59067fe03aaf9f133ff7122b573dc1aac388a95cdd79438e1f6a3fc73b750e21;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he386f4c9fa642f8de6815f611b20d1cd57d961ed5d8d87bee7ee3aac7288795fac0361dffadf80d873b5832521607a97974ca83814b10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aec67cb76ad2654d9f7893fdde59f66780aea604932008163ac2433c0441f7b9dacca4b300c3a41b3b4cba0b00ca56ddb7f752383119fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171834b4efc0d36b16d748f921cba31a9b3c95d822cef602ec80bc209b2e470cb48263c66ced66118fec4c4f0827d8b6f8322b5caad40b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38d8f590460b60f94122c315b989e12fd7f15d4abd5c79d1a1a16379f2d76dd244ca6cfdb3a215096e8663909c5a3a6c54123c791781e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7347b671f43b99bf450fb371a15024955e09df32ac05824e14ee3f4a03a5b0e36069d2b966bdaf7602c5a7c4a6ebc42cbecd892567e16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1227ee81201f411d98b470101ef205f6f8bb3e1122f8f9549ac23deaf377b418cacaf7d9c63f7d79566da0d5e1779fae183c88e697d3fea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd77b246110414f8c2158508f02c29e46f0264246c0dd445787db9dc8613e4b6a525930dbc8947e8fc5764f25c225590f316c1b29a2fb4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he99ccea24e7cdc67bc45faaa8c0995bbcfb5cbb288e4b8f63d6eaaf29d8dd7c4dd3a836214784a71bd7308ae7989a994f657d3a0c6c0f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc11259cd3db98d406b7aed1381228f8b6192a365ba2db397b5cea4b887b3472518bc279466293d8f49b609ffa5df7014cae5ab472b2906;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15901fa28e28c8995975ec9343a9e91e39ff2323ca2142adb309046487d88427f6e233c5d31fadb76ccecfd05fc770a8d7679a861cb051;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dc25922e345ca416e2a0677c2bbd4fb45144a792b4ffe32fe2ac0de1a2407d2661ed666edf2a68ed0d4714c5c6890d3a6ef0d72657e94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd4fb2d015f9bc15d679d2bf7e0c9c09595460dc30108014f0de1d9cafc4da20a523f8c40e52d3c6b797cf1d7045da969e8dd5c911e04b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b76ba2efebb6f23809640d51f0533631ad56df5f2014d7dc0f326e7749d951d8613b9304195d35cf046a6e13abac6c87a5dc20e82d5ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e41686fb83e8d4fa8f6e9bc32b7822895c28e76ed44f497ca46c843ad6df9caf04c1546e2596d508ac29c6b05413c23a5a72543db3f730;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ba7ee18858b3895669bee2bed0c3e83686addf5b2f32aa7f6d62a24ff10f0aa04444da3496540df46a827477757ebebd7712560b471a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c05b73c27de5e3d8f7fade5617100ea750a880593ae83797432addda047c40eee27a5285926e988842aa01737508688a4385e4fa37621;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h546869f3b22bd8e4ce646c04c8ddc8d637d9701322e3060091abb64daeaec621831e9304208ed5caa8855c1fb57b02ab6ed633e68aa2c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2b89db29046c61d18b01359e6b15a61a65907291d7eb9c3fdaa6c33f8b8b88a3168532aea863f048934b10c36dc76c0da591c49667a82;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h72f12743a751e43b3379ba9134818f17fe5bf9520a07249b4cb75ac85f2539cc3e20ee35086e9caa73d0e9424fbbdf0bfdece5b8fd801b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha52c1d197ce64a773fdea73bf5134a4e08d0215fd668343ee778d557f2486f0dc972f45adeb799a9063cde4858370354d8e953c29c6bcc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4c2545697942742a539daf567b54c16b05ae51b2716f09c8e8e8480f6747c82de39a5d8e15b19fbd9c776b1ee996c5b94a6b89e6b5aa1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1092d45ae89c82bbfda15fc2853c71d5be43cd9363bf55121ce2cce6a54472ecc7c65cb01887b1393016049be30eab8d6ef825285b39b1a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fba56b61e9dddd5d74d6cd7356c3431813fd5db949c5c6dc6b575513e37e960d412612e4601a1571fdc6b4519ddeb24f19bd4b27bbd15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e0ebced873fe63d39804beb68cd3a7137e9c00a9050ed7259b2a2a1221e7e46e3a982704fd130787b3b0a151726cac2eaae82a58b57dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70e0d0eef52747866a08069f05434354f599608f35210d13f0deb5692e54155ca076a37f450e88270e5907f8c87baf460b1c9e8b23444d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17714e3c54b4a1a18fa85251ba812fc54ecd362affcac6fdd9996575ee9c0c9301c9978df8bcf1af125d7f7718f5e7d8277277b8d21c71e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b2cc084d4d75cc3febd25f8e0b9ce3ceb2bcc8706b2e24640933defee59b8a871171b7e897b8fcc2092ecd11107e7b7a2b2db4c79a1a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf49c831167191145bba38eae64ba26551bbb4360dc5e3ac1c28e77a3e1af46a0c30922cd6bb731fc53e41c03032d4380d70c238688699;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e500b8571da24e11fc875da10169f5194411be56d2994375d5c2ba5e3632dc69ce69e3f41e8d70fdcc9be6701bb605461325481852f3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bdccf5a82028f77d154c92a384e554085f1ca8c287c9c070fa44ce26c96810443027d15a89d194ecfcf7167dfec04abd1a7b690ae70ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86bb55bf57ffed4717b7c07d12e1a637cd140559dc7adb0ecb5e987cf9ebfa54b54e91c1e42892fad6eecfbb345a1a4c413677cc1526bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd369e541e07ab6233f60bbeebfe61664d9fe5058cc8c54a8f486c0f6817b36eaba238c7ff648ad56ffb716d139c3f329815d00fc0fb8f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e21aa835d7452019909e6a0dd08e7614c001fb7cfda4f3ffaad8421ea415ccd50a03c578e70acfb692a7d8e09a5a125dbc0ab7811cf8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12fe5bdb8047af74f2a0ebe8dbfccc39eb8ae552ea57b7c567d854a83a255b187115bfb2519c6e54221a9519e530c9b57609f8ea07794b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c5ef38e0162e23d8fc6b16f216e41f4482ad12ef778359aa1beb72f53e6a7ddcbf3e8e89a21694d9ae92bd94f6f7648ff1996c7c93b13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c278d2b5f88ee6c2794af1693cb925238be1711e5ce2d6e6c075ec0d2d33a2928f8b01fbbffc548ea1b86ba3a83b8e6a31abe7173ba566;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb771bdb2996d4f394b0f0ca7cb78e0ef3c83dd3280ad21a0a5a06aaaf7523c97f7c4f5b2be8ae3b73f35b4079c2b667bff648c5c8032;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1644d9a3862b206aa31c5f1982362d2fbe780e7531e5cb1585447288f35722de01b0b552afc6fd0367a71ecf9b43f6698a0fc73c19e5fd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15307dd53ba1feccf6df03ed18a646b7ce5ae3c402d12d85f65369a0725dd7d98a8e93758f542cf26ae6a0e29f288c98a037a8345f19ec6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46927694acc2a6527d5c09b8ec6c863a95db6df5993aaa761625b8f8d1b10d48a301c1c60a18dcb991e6f1af9bd1e42836e60b377c8d7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afb1775f170bbd5f0a91d19712937f88c37dc86f2cfbd1e1c18543bfcf4a702d57ef7aa983dd2b1c5f70f4a69fcc72473fa60a14f5662b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb689e8afb20b46bfb7efa9579fd8adcbc7f5cc478ebbe2ae82bc818b5af02cd06e10a1a441a17aa7f0e539f6e554e9ad83a9b1f24bff74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28418a86355d9d0b222966f2ebbf994504f6f8d80211a932a134ee978992c9e4680b572f7ea09eaca0b92503a2f0b4ada88bb0b046fdda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1e7474876fd03b35b2cb601688be892a069b6df72c6b0f646b17e9107bbdb4e2397c8c4e2c470ed71bfde04dd5207dd6fd6b75813d6bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8aeba709f380c7a5764de0c4bd9bcf6149c87d0250a55ce9d802fd3da4c29596ee3d1e1095b833a95854bf16ec3c7d30264af95d8812e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1153c5fc550e68e18fccc6f084825a539cf25b37be41900652febe20d85a4f92498a674e81213894bfc9a98a331d79034ef3adfabb8235c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2fe3e389b39023e587327488628a4a5eb4e5655b3643db55c14c99fab888a1a41ba61f452d0cb8e75d7a38f47860de5e9958511ff9239;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5b033dbc22539e0da71f8f091b5ca1996c4c66feebd3a8189e72ed2c14e159dedd71628ab7f51fdb2c2d657de87214ce982eef0303d9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c57e58075c66c3c3a88f9998d85662c5e77ff2b60c8a9ad54cc14cedb46d65c2ea8e2e60e6dc98938aebd00394af7b31edf3f891b4ac0f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e6da7ca72996df106f60a2dd560de1559df137499ac3de53d7f579cb1c20369cbbe9a163f6cab722928abf4f9492490923f2269ed8744;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fbaf3bfab8e50d712cc2970dc6baabbd141877ee59e8dd66deaf4636fa54f746fc1ede39e8032e1459a318596d7953366eb20944f367c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f88030f92c7ee864fcc1977ebd66a290dbc1b22e0f6c47555a6351cb3816a812c8139ec2d1fbea6ea9db996ddf79b24d0cbeb8656f2e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2617230bb92b55947226753bee2f86c0f8f8afc27832615e05711e2e25b5ec95db8f92f86a922bc44a6f9a704bcfbbcb9d58cdffc569e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88d791f0bad730567406d1ec2f6856956aad6974e15919383ce11e504e53a1ed2702efa92b0d6fdf1b76b1347655092e896fdc717e0901;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h310bff05492b60d8875d0c5e0acbfe279391f557815d03c86c1b0d237f4f16dd190633f03110ff6cffdb725109929726901b75f1acc514;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9322f0a9d7add82478f0749aa9aa9404d959d6efa68f0842ab1bc1a4dd5c3974b1c10650c6c7c4b7176ad3f33183093f7b5c3d83a280b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e250bf1f46e7d6c44f9fece2124ac7f023c4edcd52bf4b3bf452cd6f7339a26bf6ec115642f55bea32738f7eb90de37c577cc9e8f8cd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffa9534458d8a3949772fd2a43f40ccee8356c4953f84bc24a89ee9f64f5e8e495eeb1b1b4c63dc882e53cda2a1be64406d75a3be9f329;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10aae93b0920ceaead301971bcec9ccef911f19d670296d1d7ce192723be371347c974da80d843ec54ab005fbe84925f7c42cd859ad6c8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183e5a8d39f63b48fd2e9b74c86eef7817228c424518c0f9731324b581687bd6f604321235f86470cb2c02b2150db2c946b8d5b11cce8dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b2bbc6feff9f04b1110508e609636579831f0ac8f220f21aeb35f87b85da437eb774a220f9fb1aad2479915a871cb125b2787d3043e06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48ad5b0fc4bd35bb57cf710158b26a81b8488f35b3f6eb68a6045ea7dda72ada879513b38ba4c4aeb0509e751c542453618e083002300;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124db0cf045734f2599eb6596a841bbd438f142db4b36de343e8e8e4f89abf48343876c7f7fb1ffeb28a2fcae3f7d18b4f0ce9976d3c160;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc830e77647bdc4ef738f5413ca56ecc42a1b9614388d0cb147e618bb13069082c09538a8e3bf645bdc60c591bc769e6d7719e4a60f569b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3237ef10651fa0ea4dadd2b7090c90252fb5b793856ba9c7a91b4ba1f395a96dd2569bb1684dc8b4cea827e8a3e961e71b894cf2f87718;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3dc6c486bda6f85db2b8d83ba42a0e21e111cd5d8aee17df099364b07f0e5681d3c57ff60724a2a68e634c114b0bb30d49b453ba1981e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf05aa6bd631f0ae5ae5d9ae220dc9903cc9046ec7dea47f59a06214bee06ef0c5c2ad635fa0a6c807a2a7416b0d153b1050fe8a8fa7c8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1348775377bacc36152b6a0a303a79c184f2c270d06fda8ac1e995059ab07766fe1b09a0ca7da8832bd76e5f3cdfd57eb9e7e144e623111;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47d5bac3461534de380e7d7ff6c9786c922199b05903b87c4bb81c2a6f3953dc301b41a07f48293e1412ec858b399a1189cb8bffc52d06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b02fe510f198dff202420096591cc0c45b6dadfeab451f3caccb8e43ade8830451a3bfd0ac3eee60bdb8c873161869951808b511bac813;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hffb926223320eb7b1bd1d7814d40d81bfa50dbc8bba948858e4e6e459dfb81a92d52d0f30389ee006693c8c8c685c9132c55d4d7f56e64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c8864ce04db25dcce9c1ec697d93ada25b933b27352ab8362ba6e3ae089eba913a3b71849642e143cbfe5518b2fdb8c375a7b9c25f470;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ffe0ce93ee28c868ccbe2cb16843e10455ab34db24b8dc6f5989c8210b4f2e9480ab747157c817cb9bad67ab35f3a66741b2f5979073c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb4a9aa4b5150c67bdc985ef85e13e813336cc0f3b61544a2ec1cb85a0b75123d4328c1c9b5f42c4a4e29c4752af11916156e0748bd31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196ed127bbd38e2603579fe2793c172ea631edb5c431d94dae70f689abac4305fdf9ac1170edcec664bcbe7bbd7538647ab67206d0cd20d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6cb06a54bb36c78b74d5ffcd176fb80009a5d05b892ba993da64d4a4643f1239528493576c25d182937ff9f8326e5e43cfa2c2bda21b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fd504c77ec9475db6931d2f3012a0d9848188e5539612d93829786a82171af41f0e9c8f28dd11753a0a7b0dd9c745a1c932915187b358;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c016758dce0f17017289b4c14acdb7ab6ec043126441d04e2d44504a87277f78524dc4938f3de7979d897972685f7c6900ac6c754bb6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cb1f9771c146d52388bb2d5544c97a64d79ac27723b5535354d9add50f36f570b8a927ab69b5fa70b5ec3014b8897f559165ee21d55b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bf3d67872660f051cd0791be64939a9bc99cbbe06e4ce4668301514cc9d1e67231f677151ebb306a365e4cb0d153ace6e091b8912545e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab957eec3c3f8ca2a5646d175911065eace8403963c32fe90ffb600c96dc5bf3d47706e8279dee81aaa47feb6d91e365a4d2b8e814f18c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19af6a1bbd21cc4e0f161a9cf78d19df0b47a2dfe2f37c98aa4b48554c458729e0342b9ea653a2f45bc3aaf72d4130acb70487fd15c0839;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa556ab62f769ff775f1413eae7d39091cdc986bb08f4d7cda3d0f85360fccdbc5bf0ff0074cd783402ccb35e8840654c234afc00516af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104d1e53fcb7f93cbc10ef23b3558c19cc6e2849d707c89e5b1dcb2648752d32d2d8d4b9946898259f7624d2e1fc27790504ae335ad3a81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7417022794c51272e5b86c8ab1faeffdac12c8969f3a17f3ce8b14e487f5eb7eea3c07b0ae456c9fb3975eec10be41036f46725c20cc0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a986f287bfb52d1f73a44174704a678eb70bfc3d62630afb4988c74ea9610a14105169fd2d2c5f994ce7c526b30da7f72e29c8e4f43ff1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2550e7a7b5b8ee0ee921f1f0a99759eef9a22020d11dbfbc6246605200994c8ad25e1e5caea97c7103094c085046ff2b26fa17a4f88e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c8889a953d9637189107e48101a94d933172df4a9e9a93e5df30e3b3e9cf7204884a6bf29b8e92a1cd03d9f86eafa4f31805472982b07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae82bdc3a4609b752e97ad45ad8321b229eb498a64f61ed85d305d9d782287bd860c43f834f0a59607ca53a509453e7019e507c613324f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1372dffc132dc3d423bb847f40720146db9d55cf26c447ac282506c0da4e25849fd06da04e6d07dbbcc0239395583c1d02b40cfb717345;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5e022be490dcfa9d874142a6b9f28a6a16136f60e6068e2dab0157096d2e2f0e21c7cdabcad870b3dd69f0e0144d0a4d60e34a0ec5c23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3f45d54b21709481e3e26c10a37c2c17bf4f94d6f9e4ff5b5c594dcdb8d206c33e2b86a15a570d4bbbb7bc1eefb1624ec2c299a459b65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182412d2bf093974a8cb3c6be8781b7b05fbdc3ea19d40d33e16efef6ef95d6d6d0b314411a16503d3febdb4ce91bc30f064dea8ecbd33c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19dcb1579f247a3bb393e0d7712c112e308cd3aaca35c0b8a842495cac56a75af0a7a564071122e4da8bbd4da6dc1de4c18aa790e7de6de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a26d76accc0e9ec1e10db7bb86ac7fc8a03a2129d4e5cde482d0c2a9c3cd9e131d3ed6e41c005c30cc74f147bbbb3c1f7496bfca0bad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5119bde95690673dd6510432f8229b22c092822d3233de25c1f15b6280e9e00c3fbd11d6e3b78c1214fe273ce6001e58c632aa19f2da5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1a0a633d49a7b95da72a167945a528e6c0a475450e574a3d84afc967887b88aecbd37c0acd47e55a6309369093cdfc644bd16b5f21d64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf85971afe690031dcf18cc21f81d72b289f91a1559cb7631b59396975715f772e1078bebf6228b7b97399df4eb0a52996caba49bd824b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab194fbbc7a4b773777af9e427cf7997fd4acb689d36175f9b86c091ebf8b2a33a6fbad5f9ef6db156a9ce1e555948cbc86465addc07a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb0d59efcbf001b8a1a5c8f12a3cd980932a696a218ae51ad6acba6e69d6f6f833d67c6c000ce3b0e26d796b9e9764f234f2e59df9bef4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86146f3a3db4f3d72517b0721afcfc12e96bc5dfc2195b2e5aa80d8f440fc81ca5f483b6f6515c0ce7de8cd1bcff04812d9d55fc4a6d78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9125983e2d51fdd705c7c66697b008d89b65b0f70c701a25e07ad113de191c8417c4369dd3c35712d532edd72e8508f5dd1eb14720ef3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha479e1ae7657554b4ccd55541cc7ffff285455c34420d084dd3eb204e98b43e25882bf2a35671b11eee8a4d63c46d77c2244471ac82b2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140d968b39a207eb924b300925408fc791e182c1ea0e2209c637e4a1bf824076aa3e62a9f2ee3032a1ca543454171c5c123994775cb89e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8d2b179ba0f9d83ebfc26046689072d3fd443f453297ea9024a45e533a2d3d7accb9ae0d6e66860b8ed4e333fc4a25f920ade2e58930f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e799fc254e1b7f050963de8671759c6c128fc06725a749621c2bafc4af089adde07f564fad05b39d269f13a46b78f56da43dc2eb618cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7a151745ee8ed48fee93b77ca42ec62a41417e7ac13991c9ab3ba4029bda7fa72c4ac82f9733acc6e57cb6572b6cf10c333797108f50d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd48a160253323cc0b81c772167262ed18dcd5a05a1ec02eb97e7c1c667d0e02169759ef0bc54bd8d50d10c8a8f04bccdac4bc828f4379;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1061ca7844bc4591cec67e241bccf63b5e2aa30d21f78c0ac556796b44c5af930a14aa8ab0a8a807a23bd70097bc7daf0d334756c909a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b745dc85a6cb6abb6084acad07b26810d909b1ae127330426b8c0b5858194b0992be3d58d79f113d603a650dfd4e7fdf8869ba2167807;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b79801e2db70dcd127044c1c41e5fe217dda6d25d17d896469ce0155d3a9029292c1797ed6ae95d36c31e24bc437143ef9d4a3859741d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7917334a943fc89c161e90ae890d512f8569ec6094cb3f17494b3a5f318e0390e6240c0241a829bb1182c0509cebfd9f8999ac983e3b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h25fd7e2cbe70e95303ebbc44cc63d4960ce94e5e470e4a9cd9905e3500154a2da33418bbbb43ab03aa4a9edff4ae325583655b127c48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12220369806a88e7ab4d6cc772af7fc7d3186aeb6047e5002bf4f259b917e3803174fbe3f9d173355609e1ea642df58e3deabfaa18a207e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dba53462a2e734e5246b1d87d7424d366b5749fec0fb9a9b653f1db51b07c92614c8e2fd7919ec11a1d7699074abff5915efb86178f1f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14da8fac1a029d07f5d0d7e067f4c6ee3391d2d34aee353ee762aabe66f18d5f9cf65ed671fe4e5611f16d694058f0e34760c9a40edd2b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1946af97c74bd0cfffa2441739c1a9147b3897c056f5fca56d232f8f42f889b3c71c9726744ee1435e30b49e9e1450a2ed3548fbf96b3d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80fef7e90199707374d9bcecabc1aa346e9732142ab71438e80dbf8a9d003197086a04689de28f0616b2a951e77871be3403659455b669;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a5bb3d3731fc195d2f173317e50a4e505e8bad687aa3a35e5b198e9399313df8122c02124daeb0fa288733de9bb9b27027a9cd05cb437;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1954c561c9565c5299235da6ade81e3144df5704dbf9b6c5195fe261bf00d7d26786dc3bcca7f47351e4e18d53cd7c07426d82e0561591;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa6762cb6cf3b2659c6745da0d92c4141d155004b99028bf2f1d642ad88923ffc20c91dd45f164208443dbee4a389bffc0cf07dca0191;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d7b373fab187742aae985755cc1fbc6add258c6edbbb5875f4aa5d04c42c9f7775e2ff6e745bb93689a864cd2cbf9c139aeda9304896;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116563d90cee1b3fcb3ae0053c7d00c9332ca68f2e819e6234f1c09e09cb2cd4858ceddb6d6c445789a618565d66ec23082b4145ba1d856;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151e9bf0db5f2705438c545d5e8a23d10efbac3b40c82f7d6eb9a286e816d314fe5b1742ed4e44a30e72b41fccd765ba54277bbee0031bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b2ebec19e2fbbe433dbc0d584111ab8e43870c616d79fcd8baec6ddb64ad56ebfa425a186ab40bc3b348e4c8aa7494c02624b193eb57d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hedf2f86a7721f671a5ff3d1a13276e467c490d39b0f962e5dc284c45bd5529b987dba832353761971e09949b6940188ebb9eacd3cfed94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e931c7a0a40ba9a1dbdb1e7893be687fb987b8fddb7b8c3266ef55784be5abd81047bb9ee15a12395838c016de0b7896d97642b9ec999;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e9a8ceb8a41ab6d42e3bc14e8127c0cc704e3161fa41b807df3970105fda8163ca53529e548f6066b01ee3229735b3abea0e69193e62e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb17744235923a3c8d6032158c9273741211294605e5e22289d8bafad9cbfb8fce72db6eed497acd5814725354fb8e6e8c8af703583ab3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb22cc8957fdd3a3507e8d17dada4d17298f9bbbf2808ba850481141575fdff0ac5494f373a5a10f736a9073a23fc09ca3088d40168654e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0f40fa5b7aa3b28f84bd2774db5fbb07ddc6be514e87e40ac874cfd97508e5a0fab3ffce57d4819f984173aad3008b7e53883bf13ac27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ff2bdfe39bc613c494176360f089b85142e673cd1d23bdce0d8936554fe6b563b7f71d0f55820520e3594073bd4348e9ac73ff71ad751;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133f52eb3de539765b351911229b16fe6fdcdfd262883051d88b1e3fabde5c8017a475ad34238de9be4481f78b61a8b9c4961d1971001d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f37adf47d73ef6468f023c94e4f2afa5d0415b7dd03f8bdfae03e9c94029b9b547a35fe390f6a4e95c48a26296178a088bda4f0d1912c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94f9ebfbddcf8f3fbc51df887ccee1418c47f9f38d03c029a530d55627ca25fe32595b7a59eaf5b4ed7acbb37faed9448a9609472f6cf0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1747f0cf2e345ee8f155fa3fff9ad64112c8ea7bc6e36a131335d3ef6c88286793af0fce7e979711591e4f6b0b0c4913459f4c33dc0050d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6f71b92b2503f3689314db94d049f71a09f2b33707717874e67b036f6a367eafd3fc5d3fe5cec273070552c9c3950e2ffcb37f94dc9f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a7e1c6b186d55fcf207ac3122fd64f52a6bb55a30b7911118df4715377f6d1a738b65ab7e411fac6157df8d39e66d757ffe9a31b8afaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h392dafd517fa4e7333dc7ab8c1723e1eff0832889be56408b1b0436f89584f3f20c94201faf3a14e52890b7be7f64bb62e0e642571d46a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b09f1804dfd3d72adfc4b275ead629d08fee895f236981d83ea46089fb0ca80b984f932880d465b190b3c1a242f62c0b6cfafa5886cd5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dccb6d9c38985c5447bdb2de62b9aa7bc61cb881efe6e3c4af6b2c8c4965b42c5b957f8a28e437361af6526810659950562b84bcf6598;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha21a06803d6b3cfd4585f15abb50a8b6ba1fecfa5103b73d43bf8ec0f0efbf2e7d47db77f1671d9b0b451acac3cc32baa370c10ab55842;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1626a882841638509012970e21b644d80217797930098496e307f6adb6189f9733906d33493992372ff6eeb4d0517f1f04ae91897138851;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103b8a166a20e52750a0b50c1c525696fe50337bb3a6aa79cfd929080de6263747f8cebe9068cbb5deb38f8082e5bee23a90ac4fb8426f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b4bb71eaf7a3410a113a465e771ad3ca232e776ea771d67f89e8d3629ae9b63e9639d2d41a680859d097f8446173de2c6ec9bd58557b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h858f58096148b926fbb5329951eaab7f460d0912f16cbe816a78db5a474d3b3df092aae8fc4a059d0034c384e9b16ffb38181c197af37e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffc23273a3a1531534846d4a55a8f1d688175f21efb32f960f50fa0fb548453ceea46ba32edf8a977a2e2ee94266bd5448796abf39c5b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdba57acc69d2aaf60294271b65b70a4c7989959828e888699b5ba88ebd271037147a6cc21abafbdb1927668cd38077a16826dd6c156505;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e7b34a6d49b58debff4c732ffa55ec985e092bf30485b9d376df79538bed936a7882666da3825ece4672d26e4d1bf94c6fa43b172ef12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3aa4da73c58079dac4ec9c81aa3165be3a335990ac794eceaf6d2c73ec880db8d45601700e18bc03e95377c318cf9f3401996edbdfda2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dab70c69d5f26c5ad83b2c99ad7566acc354d0eaa6332c1a26d2b4dbac33dd5a708a806a321b6e36f695b9b967569846a479d59df44c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bf87a4e5c56a339d00a58195b6c8a69e8d65caa5c95c50aab78f57185eeeaa0920552196a83d442d4537dda75ff86fe8ec4cb71995d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194ed8d75c1fbe0aeaf8345475d1f9cfa7cffcb9e0426938563fd0119ec4cc70338c975d1f9bbb35977ce40f1ab8247a4484b648fd4fa5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c875bca45f0d642d1af751cc11bd019381cf1198c95944193b40a6cac2dd886d77c1cb5053b51f033ab0106cd2fecaadd192cdd23236d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142578905a727678de7f93bf3e5aec21404c4b29bfaf06bbbd114ecd37707d7b6274935adcd63ba680c6072889ffe64e9aa8edbb19cde06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4803da0487d73ac40a4e2a0e3302889602da6051363b99fea40aacf6a212c15d5d472820e251573c2a8adf64d3d1c973d4f73f16944ec4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3699cc5d5a4611d7b666252f7e02e0b19a71208fe9c259bb2cabfa38de99fff07123811a518dca2f2134f5a17b20d3255dc2fa000eb6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f55c60bddcbe88078e0ae128a2e623e339cdc37ee3f1d545fc085355ed0f7f547d5f778c2e5f76d4b5a6e0ee7dd49072fd1410b37959c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf07b72f6a90a4848209334ee66a279c408e0f6a6c8c38bdbed597226b1b357c257270d62b0021bd231bd0ea40ad7673a27808ffc038019;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1381923db7ae35b31e6c6e225a7cbba0866946997b46190b027be7dbc3022508601152762eaa1f5a959135ad75bbb45532328801318060d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c91a8a5f1684301179fc82816c15236d46ce769e4f22629aeb102df3d59bcbf8fac3b9686b3a68005377731511494a75057b704fcb6ff8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17110d7bb818bdad4eaf27518daeb2318a7b1ccaf13a1bc7fa4edb6448c6acf464139fc9b7a71232d0b9e353c493ffa3f129aebb659c26a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd699ef2cc9af285e5566232df8eda04b9baa986856cb7373065550b35d8cf47f2e7b2ec908867558c79cd19dc2b3fa034bb72d84efbaa7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ebe5a44444d79f8567854229c1f995cdc2a917cd83eeeda9a1e942474ec5a5244120940a82ae668121758fd850898f99c67181873dc8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121f0ea68dda9e79265b9a811866942786420e546fb34f7b588a336af74828a05f556d00b6511ad81399f841fe9ea09e0cf764119dea9ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93b0045bf6ec35754f9348291a80b5b73ec8df876ff8cc3d6ea515731f4049519f0adea7c93008e30c62ddfde651a254f95068c3b8b6c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab4719447faf0b0e5efc87cfceb791ccce597d229a795d15c8e900f3eee03100062078f4206467f61d841a52472351fb6ea78342685fb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d479036971da17880d934fb1f4d47ee9131adc319df894829a6aa9ad4e51504cfb1540bf66987a1bf1db0d06f69f2f576287d741f504c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147d690b2532777381c603c73d371758e3a01fa113b2bfccf177f3d5c7cc3eae2369a0b594cc918cd2e8525ae57eee80be85da9271eedce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e1d3315a65ee10a83395bea0aa3b65ced9db25c95ddbd1073c5195fd86c0f0d64a38cd2dd37708dd3759cc2bc1577f6cb0e86cc1a4fe9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19248bece29eca30379121dc0f95f0f21863221548697fc6997a76327b4d320192b2058ec3f7327c159ce7ef952c92bd3c281c3dbe1b031;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b0ad353f6a906a7e58df0c7e594a7fe75fb4961607ccc84bad7340387866d03d971dd9e9aa18e0bb7f41701d14286cb12296d1de54516;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94cf5ec87011ed75232955db7198e487eb8d6b9e5564c1bb568969faee94ef9472fd70e83b5f0ade9fd35723ead5e09930e3975d1003a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aed06655d8eb8f4bfb5e6639716cd226eac8bb37c4f482a00541aacbde7957b0c7df477645049645119be73a9293feabfa78583421d2b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168702abf5d02d0f1f47b396944e0fe217d778d4525d6c976bfca4a1aa934d6e47b83eff779d91f2dbc4e61f0199fc198c7f3bd3b992157;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6095c81c40eb8d5c9777622d16c06af67a8998455aa9751b691bbb71846279d04c91c79257b83b452c8772ad8810c72f1fe4374659c8e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eeeba07c9344ea5cb3e375a9e883a5fcf83db8d5b5b8b20f8be50b813761c6dec8dd96151afdfbe8e538615e089371552f19101540a7da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17efe344e71e40f367b0b0716308c0abd3f3fa1f675e6891c6d5e34672e5974adfecdfd5594450411fa92ad61db75322262777379f573ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53247f1c1c562d60336e58274e8be8e14582bbc18d23ca696a68678a2697330b18326fefa850b61cc894571704c20e5d43d5ee59e2613;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1581a5777d496f05934f79ebb81f1f295c829a48955cd9079603c735fadd4260a3bc7e0a032a6719f5e0b08fb14a0b09615c2b5a24abbec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f0a224bcbd0293e29ca06684ddced5c347560aae36c4bb1c5c4ce9f227926913b19d9a33030d4d58daa35cb6745b34254f7f9a59802e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf02909fb60006eb2d5d5c9e51c4ab305896e6eaeded8cb6c2bd449aaf18d4218ca64c07f4541204cdf0ac858355016ea82d43646654942;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4f96986d6080143db3fbb53edda2bcc06184f0437b85f8e65a6a3b583bce176345b975f7141ca46b9294dddf657c1c4e167e83e3c14a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1958e4e9221132a461ae6f47c74c0d5ebc8bdf1287fbde2f6fd705c3c5f5e5e544c7b93362da73b7a4c35cb640ffb069bde9943fd197ede;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed3317d29d31dabcedd5b81cc83d3adf815d7703b9c01ce6cf0d1da3bdb8d3b59ee536341a3fa9d042a794437028cb729ed0754b71fdf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dd074d37f5b2ea06691706cb12fa99fecdad23c0bd2dd03d5ea19ff1f5cebf3381fbe42a46683791fbb5cd0c1b42abaa2a98f4245ec33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1471a280e02052c7cfaab29bb41ae688657a8b8872b0876a55ced65ef1b51714086de3042998c92adc40e54e4ef4ecbf6f5bf8a9169d4af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65c441024bdbd7569d82b0b1cddf76f75b0d52114a0785a9c3398f7dd6ecc2f17bd423e3e3195780b512ef050d8b4e7757397114833d5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11709eacbea536c0d6fe7ad7edc79a7915260a487234dcf7e15a9f5b6feb20ef3a40afc9647b534993802f3270e239b4e7d4b1253dca259;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fd57390cd31cc0b2dbf9db4e2559333362da01c67bb99148d42d3119956231b41ca3358f95dcc3f4c5c5ce4872749d3c1694f552443a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2b6d05d8f9f3b7cca7d2c6b509fa71b5bdec8bdf765ca12a70d6b04d1b9e153882614a44b983a002276cb5da1a617bc9d469e975c2e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170e8a767f72fe80a95c46f996098a07989032e4e3ac756b3c117818e1d8893cdee2d5ceb42d343956c5e53132cfb0f3af9c16f1700a4e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d8a244cda4a84ec2d81e4e361ed5e809b0cd22e431c12a4c383e8704eb53e125c17e757e8169f5b4ecec635d7f94acfab75ccaab474dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119c6d536d7fb8a8c6b83860167d4e965f74f194eee420571d38f2fb05b1fb2b98a75497d5a8481caa84d47ce02bf22de84276fff557d96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8382e22c573704af30c17a275a803d355aee5949d2bac2dad94e4d0cea4a6cf5b361ac65db45770a639705765d4d0dafd5b1e191b77eaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95f2f1988f55c8199414b6d4555215f25332f58c3f31e461cae205ec3c4ad85132ed4ff24a4c9c71e32855888d32874dc2b444f0cbab9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6659d7c21d650118424b762279e71531aecc0e53459da5fa260ba47c40a1120434bf92bfacf8d0292f3ef69085f0fbbf969f8e813ea87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc16c18c9af8e301c9d5dcbb49992c8b9d6cc3752c7c171cdd85b6a58b32e426910c916b3462af976678bfd15a3635faa12cca953d642b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1621517a096c2e953a5cf7ec2bf61ac2ef855cfa829576587ca6f6824514a7b02dee0416ab4330a19f7fa8650df74e5e6efa5bf0405464;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43bc3cfa5d92b71597179d895711a34ace1bc16a9a4bd5854eceb7dd854a580563cbf6c79d10b86781f909921cf0fce43cf46418aa91c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9a8f97f2450c9fcc8bbf0c8d5d916c7277aaa2d5c3fa58f954d854722e84f2b98094a987ba800c07c59a4cfaa05f823eddd34fda26ce1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3d5c1c46205d632161d95a2e4a0d621246a30b9bfb4215407e8fc80f9d1650af8a7a388e1d525ecf1131a685102e1534026d61ec15773;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb46bc656de4c86fb16269a03f9b2e9ae0ecf8e9ec4b70e6e0aed7e4c2309b6a37527a3da9073ed142f9f58b555d2e70c9e92b43eb47134;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d407beb746604839208440e3939b65ccf1155a05f429dec5a12dd2bb963c41bc0062f3ae12e5d98270b87f45c314c1a0cabbc09d754b49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9d71e02353b32a561f7e840f2c1da3690f7fcbfa22fa51f5f2b0d2229d0356e2987e62e6825510c9eda8c63f870d0af9d32fc9821cd44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c00eaa6db401f205e12891274d7e4d3d5322dd8cdac6e537908eb31e402f1d90ad3b380fc93e3fc09efd5f7d16505756c25f4587ba1a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a3009887c55f17b824c6ed05cc552517425602fca2e6ef7946afac7d10f3c744e5f8db38ff28c7b2f709eca5a1f6a90f8a29b8c08adf8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfeae7439472dab490291aacb3c54c9aebfa681602ed7eff47490d3fa17275a22f3130d18399c4263687f3f061477f0742c3c50d236b305;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4997f87f1edcc794566f64e4e23e9c4bdfd510ea9fccf9207d56bf6b762c8590fc48ed391fbd5647ad4d104ae6a9a33c25b0eb6218703;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97e9e6feb4106cc4b598f6faeba043056ae1c58bc778f60f16f740b3863b244b4599d8453a9f87210a504783a6789f93acad49bd47e595;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14737a9ceb807fc030b6e043f99dd00bf8dfb8cd7ad0fbf8ae4b1171ba97176e5c0f9d578075ce52c5f12aeeb69558ca2f68239a602eb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98e82fd83c5392c4cc5fa2bf60351d3bae48dc0841534fce21b81545e2b350c0f24fa2749ba2cc0df441631d9aa1affc8b10905b8799;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h818e100cba1de9fc343b631f7e809e707a5657d3d538ca4d7f8c3c0e86e1d6ce07bfad08bdd021d50242abc093b878f97ed63171758e8c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84a6ed5f7a85625d61edd5ac1db6058521ea7778789461681e6d1bd9b4f3c4b96c4403b2fb6bc75aa2c971d2baf9e641803b4abccbea2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178ad75fc7d55661b50df894380f956a442abb542ce43da9a0199aba47352aaff62f8cc725ecea311113e584d4f809440fdcde1f076c10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0fe4ea40224df37cbbae4a1eb19b72e11c58451f7a55fede24745e4448095687ad22183b90719e60f083eb4dc322cde7acb556beb7cc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bb17d215d4be6ee53a27aaf5066b83ab9ddc366db265af07a5f2f0a0d96e56dbae5cf2c084d0275d03cbcac5112a1c89efa9c676aae15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc96c3403d578bd5c6d49763076d085b993f2c00f2c9f816d5cfcd3d5855f53eaba163d86761c2168f553b2066b4b795451cc8197301e3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3f444cf2addf717f2b1597734d9eeb4763f9e545c9d23b6c0305d70e1f3d6a1ccbfb2458ba29c9661d4d5dcd37e7296dc7be3a9a5b361;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c86b3e6cde7c16a18cb840e8e2c282e8e16e06deb4fcc8b21c682b36e48945e94d651d0f8364da50f3d5950b674932d1d88143da7060f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf70a1ca4087d7966bbf05eeaebab63cad9cd2701331a879c80f1a862019bde6e0fd7dc514d4bba0a619757b9e6d94ea986757a0190ce4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8c4b565747fe968cc08758149631dbb9c4a3f8f3d98a9fa6c0414735f11ce6d85ff6f981194689b0c2113cf93eb031063cd409e99344c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113d498dc4e7f29126807783d9da404b49942d2d88bb2904cd88ca01a22889b5d87beb47fb60d2022bb4ed22e822f61f55d161b6731728b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h422829197dccb4d27a642ae71786c62f8062af5652a778b0c49cce4c34e0b8435f6cdf252f6bb2ef549d30e81837ba87d9b99d26ed5f32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100b0e65ad9d3734a77d6061d6b9de0428f2a4de75202520d3464c5b6477e09e02615d4df458efd243925fd8a2c7b417cae4823d8e05918;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1261f5156e03c0a5f3329ba9b534008bfe0edd1f3127562e85d858f5959a5ee7a358ec68d68f2867a68aa4b8e5b9f9cefe79e0d950d94d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1100cc0d241eb0a621e235b938e9d688b38edfb25dd6847c6e0845b691cd1ef3e11421822742ca92af5dc66c56ab6cab06dc485947ae844;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1076485fd9f82941dfadd247aba57f28833d6331975a4e5452611bd81d3d58cc3bd6a6d3b507868b102d82e92f6b6cd8cfcad37003e5ff8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b66e8061538575dffe33f7a4a7ef577fbd61ec0604ad9bc5837a480458bc24b79cf6f2b42d599c6293313aa9e345882e795be99fecf62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b097bfe807eec3ae8a6e6f8895c1ffaf40096e85a865405d950e90cc685878d92a09a325c07cc560ec1fbcb333dcf47c9621ea7f070d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf16b28014a6dd2547e71049ddc15e2f131714eb5bdce3cf9752759fc0c0e90c7cfc0db2a966f4885fb620b272b89909180417d145c70e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a558d56c1082d0c315a072e40b0d140a70ee9b6db67166740b20a95d6f95b744219b8923ceed19428a97e709881930bd261995ac6b5d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he71185f647c4159b56693ddca2a38ecd9b970a66ec0302edb1e9dd8590d4948ce290eadc77d586559cabb37b91a7a93fa3cd06a2f571ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ee55752c5b5aebde10c8edc055f7477e0bb6d5ee5e07ad378c43e7e700be51551d4af22c312d5b19f1d1374d1b4271db08672b6e1330d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc8eefdf0d4212664ca895068927089b26fff9fbbfb5992908d0afc97169f65a2d988706147df43a04a808c689128ea85d692403f3f53f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef58a55207e76f6fa002e58724917428d6327d8516c5158d224ecb1e7065a449021769617d07646cab270f69bf7ba8ff4f82fa039cdac7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9b0a1e23db9454a9a47c91f9e012551fb07659331f5aeff075ebbbeff128f79a63b1b31f34bdd45ed5336ec1f7863f5d5d635e17055a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4873d0308d670d85f099e6b29809cb71a05e332cf088db8d0ad5b040d3c22d1ac21c0284a1ca4548fca19dfe256afd4d6308e15211771;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185c0c2fa35d5ee2cf3f1f591aae779bc987d492bc8a42405beada08763cd72e798163c3acc1be8353f1307864009e91532dc0ebeaec003;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3315d61fe90fc216f034e025d4b98e4baa5287219dfeae38c92d059725c9815b4d11e2704c3eb0b1eae21edf2b6df6c1537d90fd635f91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd38f4e13feeea9e9d13187859fa5fc60ca93a6e8f3e527efb30b61029e24ac53367e58413cb12cca4a691e688a4c15314c63a723a2b37;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13313eb9040962f4be6396a2e0d33d94ebede38ac6ed1b7a7c191c93cd091a600b67a8c764c5492d50d87164491219d6c3d75b8bbfc36ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf37994990f565167079d1147ed5a4ac4ca1f0ee1f4871bee1890a4448df90a8c7b3ee99ece29c36f1a44f6231b446ca4d87c68c29236cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152a7b5dbb75541b0f790136cb02c9adf5f7f9613d51ead9a1e506c8ed5e7dbe694b8395ec6b5615b4e3034be7700e7b98800409e882371;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2a4e170917458b76aab2fbf6956dc7dc2fe2ad428dedbafac6843ce6fc5d732f4cccff2d2409da9dcc8b8bd37c78afdc7649457acba0d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e44cd4005a5712b61018c8fd90f22086baf1a9b43a4534f182bdfe043cb919707951c70a9df6be742d666804b79e2f41f49323f40f478;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d64fdb5b690066453d04bb5aed8f3a612c4b66193dac726f9f4a69ad2725f0cb349185d24da7d785cfca94c36b44b648f673fb3e1fc6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d369c1e43011c8eb2955c0f7e112e408afea82a35e1f1781fcf3fef841f1caddf1d54028a140a51432b9f3cb9c0b9e69b59902bd00d00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0770827bc9cce1c592767edddc5068d2ef1f2ed76de463c72436887f84cbf7645d0fae8cfc06af43a3286f462824b551451a7648bc38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a18a71bde997a1f775172d95fdd1adecf18f7082bc56dc1da4768943c1c8dd1a77b870901fce2f74d43dce13e8866bdd6cad84aecd8ada;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b4cce31ce18e44fadc3d585127aec784e003f4fb9ccced93d2743f7620ca1da8d94be261e0d6ad42834ce1e91022966993669cb5c4f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cec0e6d9aa54c469543f4a51c7e845a874f82a17cd4d5008e5e310792ae5b57f954e24a1f579fb29812f1e3e68b1f9e531a9e182de6f2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26576101fbdc4970b1054b9e3b53c7dbf60e1f2b3789666d77de03d4a29755bc89650f7af0bd8b7fd2bb4132f3b97c34ded3f04b68579;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45f018b1c65aacd21b6c7731c2fc2259c09722be6e3fb5716d45e63b77cf5c50426ea47d36b9168b30c990c994d482f1c43e5949a11bfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b85045bd066164e5a61c5dc02bb09bb9a4dee68f779254e6495bae0be2a0d4672f541481b664a1b2d9ce1417ca4b9d1fdeacdb621db99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de7ff662defafc4fbe5ed4a1e5a86d0c331a97fb80cec665929e20206db0941a42951873688d07ca817e7cc1fa72387f8c57cec1bcbed9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f82c5d7dcbdf57bbe62f46985823df5354cb6690a12768eca8f043df0eb06318adb23cb03887dca94dc89845e2252195d8f914b51872b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1048a9bee4ff8f739ec1ae941903e37838c7093ae895de82f3ba7590fb814b155aa39f3546f703335b80acb067f8a0fb1ba2b87b9ee06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1f4674cefa3ad8296e06cd0d1189e84ff6b28b015f72b3e3655d9b67e4f92be088cae3e8248f37eb501661d2884df9f0edb8e4490b9ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198a98564d15064ca79c28ecc34ffc891933450335718f1b13b9cc83fcaad98b6958ee835b247c8f2b75f891a12c42c29433c1db1bce997;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0f6c5a128a49ae32e970bdf2acfdba1234f3d65e7ff0f5985174012356a84ca0c0b14111637d3b48f0b32b300e426709c15d61e726dee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151ab6a1d9f642e964b2c156c799161d474205a9e4058beb307c39437eef38b9f3e1d6f2fff4d97bf68309814228c84cb06a907ec63b510;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h697e6d33aaf22ba8f72d1784cb79025b92a65c57c15c9c47a6a500a7b7e22ee0804e26c852c8c88ee084d5889c2a40ada4c23c4dbd36e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c053284f4da0cc32c6233f52588ab0e95ac3d8290c99cfae053c355c706ac852a9ea65290c614f1074633370227a3cc19031eb14238208;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9d5a8cf4e3549d94b5d8cfe714ab6eead9140a440d15d0b6d9149848b81ffb9ebcd19edc119ff5f4a67d3e73ef163099e495e571bfc71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bc483a3faadb21c07d13a0525393a73c7865cb3beaf28be166fb666b1c8956981ba1ee2383f360819b49ad3c70281dc42f68be992280a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1370002ee66d87efb6126eb021eef3d12a1564fb850798ae10f5163a846da413fcb2cd8cf971f9323c7e2b09045a2c6e7f864659d54e313;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7a865bf5d4f8b1cca86d31520820f1373b01cb4c0d868b252873d78fc0901d37b0364b4293520caea00a4109ea2548e294756b95fd6cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae35007eb2e5dc0ae4d1fd2a0f1542ab866b955f38d1492114720e263e6a3e4d7b7aea2e911de2e508fbadedac8f21b329f769872a3771;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ecd99c315da7da93c9d255f594426c3005f51d63693249b768955704b244896533fd91cf1a41ad7b7810a3dea80e354a80cf194e3a08af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7b40cd0a9ee849727a774bdffcfda76368621eba2f44d191ff395aedd22fa85f8259fbaaf635b11564b20debde95cd70d77da14bae76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9ce5b9ff7618efec7c4db6427b79e029e03c04bf6c4be03978acef9f0272c2890a4bd848b5c9c8d916a8d6b067ffe2e98c991bd9e5733;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16832d5854a7914846c11041beaeba26df9bf369243c5b3649ac082a195925921e7f213885eb0c246d5e48021b982c17f97da1b638b9ac1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62b2193a575cde03d331fa3ae05215765a0ff31a7a24eba7979def625215be2b9adeaeb696b594104719fbe82b7b9d06f2e17c2d225c53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14475a8cf9bd6bc2e5661e1ee1804cdb06c94d393a28536cc9e92cc227a127ec4511175820c68c77b178045f0cc822ed8fbb21814d5909e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100479f4acfccf856484f7e89519dfb5483f23b6b88394978113a33aff55f88db960783d0e62ae90bf648b7bc9f872cc37db5607abef7fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d7404022eff7f7f7d6a1024a48e69ea5d39384fa83a76af1c364054cf40366a7b171dfba93f2897c70d85bd9ce1293bdcfc4836216e46;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd7c6d1edf6c8f37f8047d69f8e5cf6980f0982dc1d58f32c6631c1f2468d29578492c60e2696e86a3957fe140f60a226567fe730609e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ce44136eda28f3c3156ea53e46b4020b41e25be5ac288b5055d50708ee4b81899c3e0f29932e71af20ece22bcecdd2ac1db3f97fe323;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6ead1286e8476999bf0bd5ac683474a588aa225551055f5ac04c6322246a1e36ef164e9cc21d5eb5b398a55837cc8e52154066d9a51d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a04c935edbf18d37a6620163b84d185f8c296661fc4d95af9c25a2ac1bed84f2ee9783f57c1daed9f373cabc1df9b853fcf6c70bb7385;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb33fa59a616e0bb0cc8cc142049f82eb0260bdbfc50c1cc8349b1f26b57eeadba65dbc96c9f3c804317d0a68682b60c2ea1880189071b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1261a8b7c6c3da402c93cb5fb0b48375811ca7dcb7cba07b4533c5a29332948466bb7640c92f01cb20884a61e92ebfb475ef46ee30d5fb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10069a006cd319f1d676d8b8ba128b14c1d77d976c83a389bfe7184fe101d35143cdb766d7a034f9f0e9d44fd1fd2b71a072523c2d2edb4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80a4c4fc5e23efc65ff7aeb1b35229e2449a1da8e968e893fc5e54efa33274be5f6d634d9835fc68bd1155bf863a60e40488fef34ddc4f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8e094d19d57ee28d7910415eb7297ed30190122392d201e2f1a8f7e79e0de1cd3637268f058b64287436de1d7a2cdda3b43a6c4e40f5d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c85b22050b49a9504b82db9d4858f489aa80cd7a6d27641800c30545ce0ee1fbb9ebf30b8f6bcfabfb787d37dc0598344bfe05d512918e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha289ce806dfa446e059b13d53e5df86f57cfa1d45355bd5c51dcf071234ee3711d9376c31e754d8afcc14e695a2f57e8a050a008ea050a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186678d4164d0a5759e0feb55ba890bcdfd7ed9d08ad23a44742a75147cd40b4eed96b7994d0589eccdb3b2fe9b7cf52da57ee1aa30e1c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7cf4e3ff16ec86f8873ceecbe1014cb12716bb4b18b8b81505a68be60c115273ef8452b3283a47da5a99c21e006b7b44b9714ac115283;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178e7ed4dfb1b4065d8a383d09d3e9c2fca41c1f24c0980bb7a7a0d5f4c4d3ad42fe1fc8bc5501eb4f1384808c28c5dc8e18e34a9e7ca29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df4b430bd9a38f3d5d8c3bb19417ec0636940bbcacab0213e103b298f3dab80e649a762aafead7923900be1dc740d6d06e6daea48b877b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88a832c644420838b50cf126c93444d69f2a90b7bd587ead73fb756f881c4f643f888574f4e2641c5184c89b842c0c4e355c7eb5fc6ccb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a6100c28df82a78928e32f04a95bf6bf9ecda67442ddfffed02d54d98be3782203ff4d3ef48b1f93b7ee54fe83ea2be376e9f43747303;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3841bec5c99d1568658132d555096e3f315790ba35772bf0f332da1c4de7b7d50953eb059c8633fbdfbeb78caff41037c2ba276d60ff3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1566c14f33e64263a4a75617b6be73962daeb3a73e3c4c606fc61bb801b2bb12c8ee3bb3d0234d9a7f27bc6d21c8ecf46dd60d64e10bd49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a491f65d0d8774ac1f89dad530895b2aaf360ba140532b99c7b509914a9f1dbd20a4a796720697449710dd2a9ec27d731e1451bd25a7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ceebe48304a0ca13e8f08c20c199ff8dc02fc55a641120b06af6fea2e74db4cd0e8e618cc97867ae3cceb8b3cc2a08b56d9188bd654de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6ec943b1e3fcc83fd7f9a0bcccd18927b1faf631ce68615db6b2619aa5d99fce614ee9d15e9df0351b0338085f18d3883841a2040b643;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de2106f3c073996da190b1f36186f243ac987fc32d129b0e940fb6f0b8b68853745795d3182613b4e44611979ac9d1808f6353090ea722;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149832196e52195ec383b13ef99a9a283e36c3cd46e17c59750de8de7fa1e39afcd8e4a76d021e55d5cd33401ab1d4d9cce9d0def07f866;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha568eb50ff2217dbbff264dbc4e73fafebf0839c6b84fec197c664fc92b49b4ee56aed67b472187e0ae042af95eaadccb1a26d146c1b2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcbe6356e6afd2f4d76022a277031219e4cead4734ca6a1777952b1ac3e0fb75d93083a25b7ef032f2a1c7162940a2e2e487a047d793f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d24b0944370c2bb71390bbe169aa00f005dbaa25fce9026bd17844f579fd24266dc304a6f47761f0b043a8c094a9d68ddf73428ccd964;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3e4142f39c4778d13ec775326f4cc9b9584401056eba343cf7079ea3059a90b84af6bdffe63024c3c10c3e52157149b0cf1ddb8571091;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129fcb1219a84d0a5a0ffded44fe9ee851d240b53b6044bbfb43f5db7cce5769c653642f199826526e2f30d1f959af42f73bbcb934520f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79ed831202fd43669a9ab64398be26f801d058eada8d7fd74754387c786d178c813c72e437d3c5c819af5b0ff8e9c79d9fbf1432f54043;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb3820b58580dc0773cc9d1182b1278f9fd14f7676cc212032e7789986220341e265935b2c319c185ecc12cc5eaefcdd2ea66ac79c1767;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b7476e169d1e39164c82051c76a100c364098c14fbbb1a5ef38c6d4f5f489720d97cbe83afdbdca89aa0094d0d63385674c7c7623fa7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f5f7966cce8e01cb97efdf3b459ad3573c50d18955e94e94442a43adc77808c338a97413677453b8900cd8bd3528378fb5c4b9520768a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f69cd5ad12aa4f18d4bf34aab151b8ed7851366069f01e8cc26e37520ca5295bf30b314e6e5802771dd36445e492e9facf77c5b3f61dce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4d731cac0a1c667f336060b6adacb17c49f5141a80040098b7fc555a583c430be38cef83c2e0389aa864fdf2db8d1271fc4a0a3e7305a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee68b8339fd14d50830c42eaa12c17b937651aa2fe22fecfa7f658670f7454d2beec20d0f58c4cdaa8b10b047ba6f5f6b847557fe62304;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h552d58c24439f6aca5805787655bed3a48bcc3a062a775823eaa3c5950806fb5517696b99722673aa7df6c3156e9b1c16f636e9062290d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f31fa32b136883cd96bf76678a44d40b739ea9b9dfbda43f2c80ac10a26deb093cf57356a0e759f2eebd97b850fd83c6ee54c1ccdc917;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69167e2071c1480fdee3d615e0c8a5af9033496e95af1e6b380c8d92682f8cacf386ef0f49a8460592b706f14b0e96161c6513ae2476c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f60d9d90e9846b885036abcae3899e9e0b04787e503fc18ecd0a3082c4b9921d710b4c2cfa3b4caceaa5bf8fb8e3438b0dd2bc6ebcb87d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195907e176a905ca9fa3cdd654b2b1b93f1d439bd2fd1065ecae064b755d2aee04cfbb57891a580eee4b371d603e2c9c960d5b9d07cef03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4f019382a3563337baa5cfaa691a74d8c12b87eecc1ab43d04972539bc74b80a25eaa0c06a81943cd595b7e4eed4e7e8be92ba9204fa3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159964820eb280bb48e3acf8c9cfcf48f41824a85857517bf24c27b70e7d834a43ae54f78200b2551cfd35d45f90c4509cd50f43a777775;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107559aaf4651d7d998455f04d1d39573e0a201b4ecc46f07547c115995f3d3842806cfabf2b7b277af3101ef0242e210244058ff576a3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffc10f176c21b591de01ae5be7e7233d244dfcaa3d0c36f29d3b339924736df80cbae23a50b0cf0ac7d786ca729b2bf1daa126f21996e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46a532ccb837f4a0d52f87c83bfd142912effdfd6a63c45ff7d929c29b57b9866419926276d62c388ff1ac8b2221727d7014f7c3d0b5a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd47a2e769539125d6bf1326c707e71489e087aff928e9b25d0c5b5ef01fd668085a4da32c41ee64329063f344891ce7678b52d819076bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fb2ec278b70094109f8d5912e51cc235c7478438aa5a5cb8cdf20e4fad82abd3e8cf66a68ab2ac7c1258252abafcedd63100ed2493582;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd94a5a69b3c19b38deec1a87da63318d4e871e68a1bbd00f55b448d439a6ce45351703aae47979441b132ace93666287b528cd0c17932;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2d935e59735cd089103a8d62cb247d8a963992f0835afa622397eb3159684191eafdbfa0f523bded168a36f40bbf69a9a49e5b35fa8ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bb660ab52bfafe5d51f255dd7304568141e920e0491e8952c323c7b8b4496089e388424007019161432315f80ea91d044a00c739bc28e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6b23dc763e9886b07bdaf347d01e1470f69fb398feba2d937023da1ad98c3f468f9b03cd412a898910ed06ccb0514e91ed78530a3ed3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97bc655c7e45193b0c2159ca64f1c2a4370f1ab3e007b35331c32749cab93a8f21e43ac8b9bfef2591da7f20d4e6b66f06664c2a9bc60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h148ad280b85a195f2b21f6d6c17f488d46fdb70774f515d95418b7c6e24b6b380d0311f82d122d124eff161ae91b07ba514ecf94c4b407b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e356b6b52ba29e1611742c268509905b7e389b0948854b8196c9f2ea19efa88cc40e87d0df445a28a35e0acd6135afbcc300b94998628;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e6040fc4c60aad1bfbb5a093de3deee7d8d7173d780f10eb623458813a01e04aa8a7e1c5ada2cd5a07297e21524e38537f9f4248361a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7934d7554fa658b715be44014c6223f6d7c0e3ac2eda2c0eab555303a4dae6145a4ce518016f1ad3837795e6a65befc514bc3480e2e9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96b736ffa17cd18ee5d56f069141c2703dc5a49089f299f81484ad6d854dac61abbc454bb0905a5c3fe6c11b1cc8f8034b861bb487e0d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1accf539031a753f6e3f6ee7ff25f1f0bc8eee07f4dce89c187655dfbed81b271e66ee554efa08a39389cb9d3c56d36615ddc1963a645c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbaf016e51acbcc017471ba571a303b61580d28c71c5684aa495bfce0b7543a609c80b1864a88010cf8cd5dd581b7b484e63d28f7ca06d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97feb2d616c8a46aadee13270a9802203af61fd8cc061827f83a8cb20b39ff38a939aff228cea2921bf558c19ae5ff760f1fb99535f323;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9de818b51e5f0e4da86a1683f18820dfb68aaba9c8dad7a9ba2c310f78894717e60c8a6c3c871b07c44476a19a36f11a9f33660470ef6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a16a471847e92812f04fd907e51c1d94742e406894acb93fe234f0c2ce1d114f772038ecb6a3e741e6f30ab14ebe0e41da0ae97ef66594;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e6c93a6dbd86b42ec22591114c72836ff25098a318ea56915e8f45630853ba565ead7f61611023ce100081b9b48eb00585a4a72aeadbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b2e5ab601af05b7cf6d929d7df6705e9cdc459d2b7d7e8eb1d2de67f94de3b13bdf1cc9c10ae7a2b9bd80ff82dbe85c69d5402275a5a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e45ab98bf14c1b21ae1274bd6bdf28003f4cebb9394e543643d6d665c7145550dd0e1160d0816c1c4edc93fcdf9efd59a9402fee0e44f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb526a708cb299b199dc564ce328de8e7fa1b5fcbe888ae8f12e73fe3b3cb4694a2661b2381b01cd81ad067b0f8e07c6e9198b26f16760;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169875b8220cf7de763c08be48910c13ecfe82a8f800148e5a9b18d2023d7a413b19499122fd2f599fb4bac7ca1ef881c7a7f045a5f7a17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13db5d14b09d2871454fa55f5e7360d48a9c1ac2b33f767ce7b38c23dd619a5b348bfe033b76b543e0c01ff49158cb4d418a384cb09df77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h661be1f5aee29f11fd008dac8a2a9533c62bfde6ce583f332e34dfc69ee3ba18124dfb9a371b06fed3e827ff2351af027630d1b9021b05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fb81e7ac86811065e7434acac0725c7ca987ca7f3895a8f3223aeb0bb9191e17268d00a53c4333ad9a66501a78b3d13ec47f9f7514968;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb15215fc3c1fa3d8fb3afe9e4182d858a7ad738cdb4c2abf9de360e92b836ec02506348719cca53f49aff88befa6870d1366d36f4b82ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18eb9437fa5bf3374e8d9472e814e0f3f11d4a6350d17524b8b9f37794dfcfb47bd90e3cb0d397f5541b0d60e2f9e16f4bd3038a157aacd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3f81ac07ea770d0ab0bc0d14728da612bcb7264f68dbaa4cf21617c8a05e908fb3bd80c642ed2f7ddd265e9bf030831ba03818418db7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b44926434d9557de6627670dcae61b3e4b448b9c29b9047b2cd44dbf4e4cbdb61ec7f356f11f6d6ca8caf619a2859ba977f195cf37a16a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb14f32b8cf0cf6b8ada8abe09c1f2f4afe5ec0bb4b6def01d0f64adb1fd15992a055dd4d71efe67607bf703ca41efe2d428ee970f1394;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124c6523ba129c4c40964bd0a2678dc145e6da4dfb399bb341ef8b482b020d5ad1a3a66f159813e983942f5cae0f9e63daebf44fba18de1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h158b92cea4d7861d6b0dac5e6598e4ae2dd3975515d472aabd03f06d21e73ae539e8b7969c166d623d71ccc6205f42c05056c611343174e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1371e25b5ab39dd196acf06577f3c77a203057e885122a1fd6b0ac26ecb86b5cf639b8256ef99b8ee20b99e49bb84e401210acf2cc55833;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0aec9cf05c7b8907ce1934d43e4d47c6f5df64a811f3748b183707a5f70e3078dda9076806ed0e37132ce909e0822c4d1a2efc26105a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31a73702f647e4b9b7f793e2a7e810130e9bb8900ab56a1392e89b71c40c7186ef2a054eb24cdcebde16e8a1511ff6c421c9176108323d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf46c51d2901fadafe20f840cede8433f5861919d6b3c2bed05e566510a84a5c1542c5e83e596638437a8f4b42b245b5929dbd81b66d676;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e01a6668f50d881fcd0daf6414b206139ac36f320c0fd54fa50b1815f81305a3836b5365aade60c99d8896580391a2c00e7e00c38f46e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a5a22b2930cbd327bb9185167e55914c3cba3c816fa9596cb2b86f95d0663331f01d0057331ee77b4bb12546d8410c3e4cd60e782ff9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5655c641e721a42bc61bdb278c64a3b0be6a6167a61f7665e241b48fb828ae13deaedfbb912a251028fc5547db7ab2943ec95198c4a24b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96a4d8b8677de9db336423c1edbfc5387ca8824a0b12f5c6a2fe876f26983b6310caa9eca49791b3d7d227c62022172155c17c485a26a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151013ba66b9f5fbf586d2ecf3dc06e0a9e3794bf0206329c2a118dbd6b3181c844491a735ae8d88b9c05c7fa5f931c2b5813ddc38fac76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fe9011bd68832375316dd4218de8c4f4b4f171dbd511e69019c3e0d520985255e7d55f8c7ecea93c80d178c7eff488ebc6d458bcdb454;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f2c8e2218e90d1683cbe60f6d3eff23514713d67228a75e4bd2c96cc358262e0c62a2c4034886ce6db5a75f7cf00bc835d7407f053e81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc14d82cb0f21f8b3a4b641b398641713fdbfb9a9aa4653ef5fa6eeccbc85d82987b016cf803c6b125ea1312d987aedbcb73370a6c64a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1148be2009a999e245e1a09bd1a80d4b33b7bf0c6e4d0993bf5462b2abf4f163d86801e608abc813c06f00f811a10bc8345b673d616c428;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbfaf1616e06a3e7a7388ab3ba3feadfc4eadd7eb42ca6917404aeade06cb166812e09a238630701dbceddccb1d1048cfc758779dca0e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16849fa8aaa414fc478f2c2a7e15d8c910792865e3ac6f601f48e6496e9a101955fb0776ffcc9c6e5fe27b8b145dce70ab68e07c69624b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1804f99021530b5add3d279b37f87d4a6da2613593ecfd1d52b40c89ea7ac9ddee24b406c7d2a96517dd08f81294ef94a9ac57775d804b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b0c4b311d59f98a3d0bd00858d56e9f42008dfeed2ac56f18426d7860018f8895618cca363dd143d2ddc99694f355ad4d6dc662facd89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heed2ad29a77c1dc0fe70859cdd39fbd9b4d85e4977330be9fb7f42e159bcbf13d0806640115422ec5a2776b3781efa2b4ce8878b0de42a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe5ce3c6ceeadb9ebe9234ac75c68fd4728b930f830914e9501ed7864b4060066de6302f10f86dcf2d09e64ffee09a098b6baca6446a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca52968f18a81738627991d3535c4b2e317c662f2047279927dc8fd410c6303a74ed1e7481924c1eb68873aeeff60e49de1acd2ada967b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122d09f41e93ceb89983be653ad752e0fa9ed05b98ae1f5d6c2703e53e1cced007b1b69b671203a5098a45fedba070ffe075df2c4c8fa99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he709df22bd378e141b2729fc3b148211db6d51d5ea3e1e58ab9a0fd1c86fcd1804d1a7d8622b558b1ddf2e966b97b810ceb8e59b7269ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166c9f27d0fdd959b3502c7e21d32f2fffe7b7c649135b759e8961a9434eb2b6701850aba7dea3d3701d1f9f9639a7b9ed7db4b56d95feb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4808425d4e3d86a97b5512b60ccb817d581da8254758a410fb15c4cbd35928e1e6ca8e4cf17151cd86feb72b644f6081274367ac49127;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19d59b2fc9a115e3406068e909c3bbc45c7f9ad724e3a7187b1906ae50d1b9e614c66565a04f6026a77b953bd27190ff4e91a56c7f6f66a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3c48612ca370b0fb53d7d3f412005b889b7c77a10aaf0aee42ccbea0256af3435d44b2dbda41a1b02a18c660c373db65c3f73786503bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6900cf882fdcd18ab01f82d1deaad1f4c39e8fa8ca8f82c2bcaba32d2782ea51a565d8ccf422a23c94234612a942fe9a6ff5cda36a953;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7454beb84014f11d3e25ec70b38620dbf0275bdfcfeaf93e3a3b1dcd02bba8c8eb030c741894be68cfc72b08a49b76aa4d93b9023efd75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfdbeaba5e487437496c8bbe04319fc5047f511b12a4bf3fae1c0edbd095760e2dea125a67c45d79f6aac054484c9ee5dcc2a909fa38ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16496cd50fedf04c45e62ea0333078e3c19a4e991274ae71a2201b55356f40c6c5d9fddca34e80a7856b9aa5eb081656f9e5f0f5b6c15d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120f8a454f20d6f2d7bfa8e12649fae4a87da6dc9adf80e20ff0c3d877036788e2dedba30312334440220b87d636cdff2e27bf9b5162bd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b364e85ee6756445a670fa56dde3b267b87176c7b3a61f491c12115daf75c2f815a8a80e107f548f15beeb169b0a21e77725f5df4a51a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebb122cb7507a84689a18883e976480e6a75e267dd70335172d02fbe5226d9350f69ff748aa51e3196630849dde27b0aa412c08f555d29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1690be33e6ed48020c8c4e13ad7b3e44236c299e615b297c33fe24b09f88d1827c944c520350d714b558b02d00a1db920e14076e59d8a72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88ec33c65f8e92859c42d939a5a14c66eaeebcb3c53c2119caa97f33d0c7df7ab9cedd12750ec93eaa80bf782d36d656953d627f408450;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7b3228612f8baa3b54d69e3d41a572e2d223cc3aa1c1b13a42591486433d427607337abb213d11409dc5dc59aaf468a69255dd7dfa1b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1365fbba34319a3a686cb6ede716374b44361c85614db4cff5686459b99bf4e83bcaadaecd8e0735f361bcac6bad41d6140ffed73fe50e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d10adb793ec9e04e8f021fd3fa2bd98c03d5ab18160a5ddd5f5115fead4f85ef2c23b62b73876642ecef69a2ede22b6fcf3f54ac94f74e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc36f264ee7709e82b898a7af80f207c4e580942d3c4ef460cc9b43a4b27962ee2e6531e665ff0f0a09da6aa38b50cbd7ce3a2bb64db95d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ba6d133dcd4a5a0118db70e9b1fca364b8e196a0ef407db840e31809a5b45e003c500b350c19619e1c32ee837b3d7c669e62bccf2ab94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8ba495fdc3860509951f61d687724d8a2c0c3fef324b0cccbe80c8dedef5223f645349f52d7bb372410974b36443542e1cc142914c09c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8142729bf0cdb5d9281b9aa5314e9687f6513127f0cd5eefa88441fbfdd8f895de19b52fcf6a49e10083c4f56a45b12874b145ea7d31e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb97f1fc856d97d5ca743040d4c44602462d8f83cd84269613a4da842ddcd5b86e513ddc65598b44f7cee8a249588b677da2720bfa6296e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h710a98485bf94f0fbd4e52be90a2b193c5e11064083bab0a30f0325f19e64a5f5459d423ccfded1ce5d06c9bf7dd7689318b36727d7570;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1495562fcb306475a1434f761b52c4a310265931dc0b081ad81ebd2bbed5ba1bc015400772da9c2ae032785aedc39c4a12b7db18fcc8cae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188c3f35d9bac13ec6fc9c2d1673743fe4c8bbfcc817ebd0addc5fb238af8418fa82b58d8262b2d91b32575a0957adf0fc5de60ab5133e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130e56f7336752750c0e0e368b9128baed6946d17e4d77cfaeec8ebbd1e5ee5d15241510d1dcb117a188ee5bd9b158e63dcf076c9b369f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1844fd8ae669325505f91881298feb6a978fe9a39237418fef038d1cee8199f748b8bbe1304ca920513c098603272c9e6bd00d111056152;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1a422c1ae362c65a4f1f0da6f89b973397a5eeda34b91ef81e20e7c4539df90ceb2abf240b05dfefd3f041b57a6a761f0a2fd5b049741;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27dcec5d6764682afbeaef12a2c4b8e143ea7ac5961c0adb67b76b64017af196645cef8427523851aabdb43e1cb43a2f265291f7c25368;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca3e02980b6313cc38ef3e887b5bef311c4b8c2dfe83262ee9225d1678b94705a17a36d2dd2685cafa99fbc02a2408d45762ea0a3352ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5f1905863a266c09b556719046b818aa7eb6521ec94dc78ff0166e964a366ab461a4b48098abf448564827b584c7b521b79cd2e6f4943;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18993f1a2e2afe33dfc91f52c376f36e6cad3e80ecf9416c4d71813a632717146cf29321e660544dcd4497b423aae2481dcf129b4be894e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ef52583c5be22f15ec25015b84cf5d8a0304247566274391e97238eda1e194ed71adf66bd602a9c56f06405e37ae3fcdf8ad7253fec27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c43ae4b961217a9775573ce96f2fab492f958f7d94871e8fa9a84bd751961a39128d991697b5e8f7ec9ff459250a5c153cad58300ad764;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd3c03c0b0b4e4b13556f36fcd094c6e7ab0adcfb1124bde0d0fe65376ae477f66df4f3b8b2cac40b423c398c75888ea5d68903f25fa5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15574f8f3dfe1b68ff897c316d05312ecfe1b371ef4d2ce3e01f025ebd9ba6be862846ff604c0d0704cb1a204932d30938d2ee3a26e912e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0b97be280ce3d7ed043052b04121cbff9de5687a65ff5ccb74ff4c0a5307f9c1d7681da835bfb518b368d835a2e1c500dec546dae4a9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1deb70372fd332e0c2642fb05a90f4edff1b53cf283ac299473e0aaae4593b38f4bc386963b74fab0a945b9da1103bb558bb922c7259d24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c92cc625262e376dd53623293989e1a44ab6d76b60aaf3bd55bcfe053dbde55b77a4b2ed1a3d64f4fb6b9f853c91759e78a92bd2b7d68;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a5586ac14e93aa2768192c6cd9cd1866195b743cb7ba1e21a663e9bfcc83143044dd707edeeba92bcc0aca41699989966f740c40887e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h427e1ee93df3749c1075efe6c1dac54d36b3c6cc6550c2f5302542e39c6d3427e15cd52a43c45ac4e4be55e7f425c08d49f21d0020fcc4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156b5bca7d9faec4da84bf9780c8d97ed2adc6b788a34749ee741d1f22f5cd2b1ec05b5095538bcfcec597d6f3c55376e35f4a7303ce8b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfa674eab75546c3504a5358f1b89d53702bc13db4dd3417ecfd8594cbc66e47ec7d728e8451b59c323ddcad78a870ee04f968fadfafb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bdab403f86cf461247e6b8174cbe0ca3e319b6174b06c0fc1fd4d3810a6b445a5e27548e5ba29b050835aaa55a29144b1ee80e6023444;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69f82bc50648d20de1ca01b2735738166ab91f84f8c8025d526d6bdaba5c2c28c8b4592ba43e1497ae23dfbe9c73932a01fd7eb062c76b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3e462d7f25430d9995f0a442d7ab98fffe3c26d2656a5915a3f4333640e70e2d312a8f02b50dac752e78c6b95d40d5621741e657e378e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd065956b53c3a5f5a9d1ad9d656a05641459e7ebe9c1f4fc2493c878f39a5219d9ecc9b84bdbfceab20dc310b59a22e1ac37db63ebb557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139466219d9df74d6e581d29d90476a263214da64bf8d7bec83561055cc135b956bb09f0bbf96cae7cd855a33bede4f1860c6426b10219a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h343733a3c2be2797931378530812d55180340738928b1944125f66c174320360b8c8cded29dd93566e2b9b482a3044f2bb08a9ff4d4652;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda113b633ac49c3e62ad0b95dac1929f05bbb86c596d9392865e64c1a4201dcc0e2a5fe4cafc64fcfd2e50bf36ab2551d8ae284a57c561;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f5179126ab61502f2cb13189127d14c91a97ef8a72820ab4eeec243767180b8949338ab4075569502641291a7fbe2e5d164e35771e63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74fb42eeda04037252ca57ec3010c093943faca18b2c6a9a008f211948b347c1cf8859fb34bdc42cc55bbc5e2038f7db8488bf621fcb7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b30a6bae619c320df26175ed08d26eb50e012e7a06cc50ce66c22c89f6e20f5e5360283f2a733223308595fc1eaf9bf88a4d85378e607b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b66c2c03fcb815100b22950def10039c144e0a6c1b1cdf3f6c4ba36233b1e7aadb7f9ad666136a7e95a576cb987066d05e13fee8974a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d0a20bd4095cca01e6d0332567e7bc97246feb92a9c69bc1579293583239fa5eebc287216aab8e713a396f08ed8d9bbdaada69a390e2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6280745fad4d4d1091da8cf9e117b07e62159c2ea4f9da35fcb72dfc5bbe998571892cecdbdda902391111b3190260e02731a86ae7fa2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10be05a9338ddb1666d5faa95f6a896ec740c9ea4c7b607391f87c743cda223b3117de222a635bd9fc57caef83e6c104e9c6fab34ed19bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h701d384c60d0880e7062372f33f0759a30b194127eedbeac93a468b633dc12ae98fbad6940b619306e661988d4bdd362f40b80676217b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e547cfd66d9103029555fd993deea6c50b72f073dca6c2e3c3c6ec59c4f9b17ec5a76d89f31f92a8591c17cafaf67db6e79933a1b809c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d718c46f6dd6867e70a76a10e10a9f0cc75f09ffcd42891f5a62259085ff9bdd88391e5b06ceac6be6ebe18a1c6c030b345cb7cb1299b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d3d4a0ddf0c62917f09fea02beabbc2b81d3794695ad36c6a7498bd6a58c5d0b81c36debf1b6796722163f2957b58e5d80e58245cd51a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b5cc26396177970cea45014513535e4e6b23575aaf9ed947d4ffd69426199c29fba7cafa1d406ecd7f8645b0d7cae4d43815dfdd30f13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43a2ae8b6b7c08a4f4e507e6579ab78c97e1bf2383b824c290a4256be05efeebf737982a60a0ed1d817b4c2d7f889e702549bbad59fa0d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130bc50468c3588fdecfa1acd65a354eb9376b82e436b1917614ba85ec439e4bfcef5b14de45ec063a0809554155941f43d70be59c95290;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf591996690a7c1416652e174280c6ff9e526c386b754ea70e39d7d3bab2e5e4add067ffbc62493706dc6594f7697300c87538cbd608a01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc5b922b513246bf52c0cbb05f7a752a9701303c2158b7add70442f777521a3b3dc172d5cf79292bbf4cca82e714ebfce79dc59c437269;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16600b4000b7221bd4c57ca40bd0b4c495faa2c365789d61c5b6b9991b9f3e1753f71a60bb1a9feef283cfa3a02dfe73a1a81cc40415766;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ff31171afbd15b06eb1b0ec45a5e482f6f81f6e337b3b84119b36b4bbab9a112ec8540d335f657712324ba6f90ab1850d81bfc5583bc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c8e169b5b18fb7b657088ea3cf8c9765fede6d1dc1491d918fc1a84190938271ee97b3b7015b06f888439d3331c9636135487dbd51347;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e37e8827a3237daa33c80a1672030f468b546190d21006def49d63ded698676341930b8bba951ba3a22be0a5b0d9479066cc143eaae69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76d5c17110291d2ca77bd907ea61692bd7befb4b68e8ed52746cf03e0b9b449e3b7078453c1aa001a184713a19e0cb5090d0808ee7a81a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cf62c95e71289ff6fd982a040b204d2e7d7aa18db1f23d5f2361b4514c411187c9866bb47fdcbab1d2b015538d3380a20322ffda4f6e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172d6989e6f23cc3dda49132d58abb6fbdc70ed226593f17c0e57e641456e2b754cbac65eec1f3415221bdf616910604fdb017980b7e935;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4186cc193d0a70487b6792ca51ddc88540143f7b9e6f3fb39cbf9d93cd59f433dcc9a8e1faa3b1ad163fd049622edcbba434967adee169;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1e719cf9f151ff29492dbc36137d27fe6eecac545943c9d6c830d007aa16df366ba63151f7e2a9ef188e7bd10db5374108ec54094a950;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2addc4ef2f027aed70d528182bb11e20fe570d55e43329a8b328cfac9f1a8859b45ec8b5779ffeec3fc1ce9f91033734d6dabbbb1bf990;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c99f47204e4558357a9a2bc727090b8184d6e8cfa4a448e27d6142acca7a20f845ae1b719118ad5ce50ea4fece0b5e404c6f7d4dcfc87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbef318cfc88efe37216660f16d5a70f7340460538e8ce515a9f71139796c73ed2850749108a4abbbdfde82ae3cbde6e24cda49d54e1416;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bfa234f2abaf41bf7e9b9acb14df323fa8d14465201275e7ea0e485cd90130b56febab0853305995217721f04b2cd4c09aceebfbc6d80;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105c9ebbdf0daab32d62faf40a321963cff223ac6765f613f2fd55517d77a48b1f7efe910054950d21d60eab7841d16e73bda55ff3bc84a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf517d2b1ef7ed48ef9cc31b481c861e2baa0520472fe24e6fef6789962ae8513bf6528e028788bb9dd8b653ba1d3013f935a9f1257f253;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9167720df64c9a9fe205072b0301099eb5751db3d950f6cbbac1cad1c2d15617f2a666269b1975b3d27c51fc2357d54c5017e7619528c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f055b73e33e6bc2287c469754564820115bc07b0b69b645f3392e768b0065ff5555a6a7d294e7094f995daf3351b0745989f91ad1c8a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182c6fc8e625a58dc5e60822924a4f0d41f0465f2d48d4680254800f1493569d01efa47b0d7c1584933d109b82a8c6812dca1a799a016d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8fcca2a7f1e7cd7d5de8fbbc225963588cf59b93d06e6f0e2cf56a555705c1e385252a903cae9b8b7be96de4be37f011a3199483a7cded;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f96a76db1d1c42237cb486b1fac7110f4ed57f2c1e79dfd8f613fd720f98149eaff359dd22f8c39fa75c3fd3d1691c35974b8ae12e1ab3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12af3958053116220097ef47e1a13bd39e44d9161623ef3fac346a1217f33ef1837e78745f45a6f27db846d13c44ef7a182810c42603f58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf601b79fc2e786d2f5f0e8b195aeebc8df747ff108f84db39baaace0a3de85ce8fb68a189238e59a957a09814c5c6910b3ddf36da9de42;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15706e8308957e8c84bc4c8967f27cb4c9ed842c59f821573d6de083b24a4e8e9be87a7d8ced3bd871e04797ea8ca28a06165a9348ade4e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9720f9f4120166a802d8982e18e79fb4eb45407d892efa8115922ed02d0c380db4869fb41d7ec549274cf2458c2b44a3ea58cc5aa1c323;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f9ab7497a4acfc8886c83ebcc0fb626b1f4b000c9e775e2bd7a626a9b78cc56cb9d621b8670d048763b94064f6f214adc2769e03aaf67;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd615e03dff9655ca6417a4c9692fb87aaa05ec6bdf00e3b5b3cf32eb87fa27f51c06c089e2ffaca6ce3f0c85360cd4e229bba709c055c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8092d7841d2f3a41b24afcbd69de60e0ed8d4dd3f56322b7e4e93b91f1d73be029e81ead0310d99aa3fdeeb697daf17f9db2a5e2d49e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bad66a1e3a41daed4a5d8cdbdb3aaed25a15fa38d2c881241affec7b8b80def779eddc83ff43500b84f84f11ff3e36f8b781941f2a60b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d9b5574ff9ffd7fdb1a870382efeb9ed1a4fd5925963a5dbac3dc6af8c38ecb06e29293e60372d232796a092903ccd8ab243d184c5bf7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea7780a5ad889471bbadf9e794b7c21a1c514b8e42e4d816193cb751effef2918b7053084b3522743cfd49a526f115d5ec2a68b40a8b66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he02b36a023d0d3c4f713179a21243e7114abeb754da0855005d06c3ff81344045702a84bb8e86e47fc34460cdc5db954b14173c78c7cf5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ade3e1bd7973da5b74074fd01306ba98269067059466ee2eff3530b191828f33f5baf3c037dd5446bfcb6501cc58f991aa399b3c01a311;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb271aca3143626874d753c2ae5838830447bee274b82064f2602f35a3f1f46c1494c4d4f457eca1d1e20878052303657b5668a37c7dbc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89b9a2a676e83c14b804c7342eb061d60ef0b971981de2aa67ec9761c17aa8fc629c4fa1a89c38d05c3f9cb5f9cc88b9dd56109324ef18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb53f02d376a861e29668c5753e11efb84ae998665d693b4d3bd514ed60870ae4051b61bc4654a9649ee99e7c7141ed791c946689f1bab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1094b15a629558883c407e461390fdbcd25da91d443665f95553853dad7b86d6bc28635c2845958fe8a914e4e5f15ee6936367f0c86be30;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4af3020dbea449207dee7f792f8da4194c9ab170e10749035a22c87a4f9203db8a189ead3927870a4401ed1e46a17b4287fb2d133f1983;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ee296bc7c13ab76ad7dc54aae1e46293faae81aea191cce09cf5d54694e9edfa9599bf2653fb6f6664f8012fa32b1838f7bcadb2ab25e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1713b074ba7754549049f807bdc05d7cd9f4bd5dd9fd457e71fca79ac0c58446f2a5a3fb6e18968870909f35f3c18c8fa481c177be6e776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125d02d36b3df0baf89fc03209800f1b1071c852970321fc99a0a39d03c48b9ca5d206f033ed01bee2f58c8eb83ad9b6a833c537f619690;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70603dcb0915e611b2a1626ff359eb392d65de70b6a1f623a3cd884eb7336d1345bbddd778317563aea30a52af81144a80281cc34bb895;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100e2d1e6b4bb3f67e70d213bb8e3f76151e341e71a36c9f1f485e4a2d75c1fb70af20dd94cf811bd7eaa06088558522a106d061c2e506;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de44345782c21827ff03b2eb9e7e9ddc75664ef9b20f63103dc38b08c6408285a54854c5329c40b403ef558245c7efd7514c875e98c148;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73b1f7ee02fd0a814cd39b01530e318a9c43c22c5012f4bd1c6320937587a71db0f88bbd72c5ed266a14f7be14211411af54086c72b562;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1571714e1c0ed04c2c1a6b307f81396436f2f9d22b5aa74e151e946fb9898342ef567196b865966ae16f33733482e92cc422a945d737455;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc4c3ba712fe90736ba8a45d48c04e8b0199e34fb7a50bc570e3f1d6f30ae60b6bdd11e099b3d5ea9106be70d576a01789bbb4a606d6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abba9a2c26409e931b374817f38ff7fcfc5068f81eb0a4b86d8731f35d74db7ba6b8bd7e0ec878edb5aee1e5b13039fe454d6a43165abc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89da7248dc7299acb9b338291764abf4e83c6bec1da5067bcdce8f51f0272a3e3cd7ff5822c8afcada44958c8dad46deac349fcda33faf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5b973455ff38833577fad8ebe35198d1d8442b9f7eceede3381f2057c543be5a484de5369dc3f43bcf34aa22baabb597897660477ec4e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca6017500868b1e899a984f7357282986c201cc8f00aac60a0e58954bc9080a7f1e5c1e4466e767dccde7c8a712a1eb107e30ec24edcb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9314dff6ab9a61a2e8b9961685fe9c6c507bba8c676a94a223211e22c9bc56cfc1175a6369e386d5a54a35a5daf16d943226a3413e7c8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde144ed3a0aee262bac8e1f676f0041fc608f78557906930f8e2031d5a95dd37fe974b99d49f6a46b01c36d475eb71be4dc735a4088af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc84c3e1bd839799a2f756e1abd8c4fb0ee8246854bb945d177ac2f1532a0077510553478eb5454275b0ab7f9eb62fbd2a7e9922716f816;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6df318559eef40bb2f6c5ce9df0eaecfab10f6671e4b836cbe1ad11a9333707d463bd373083cd60f2ba4b370d687bb35fa968e595c166b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f48af1d296791c6a3ce0e875967011eaf8340e3e5beadc29955a51efc4879012a8420bc55c0e5f6af1901a4ad85489c4a52d74440fce4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf71064f0f6498cac1d41e5ef4a8982c9f3784d73784428f6201c0a2a2dfb01b1b87db3da1c3d4ab3a98430f91bd17d82437bb7959c043;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36f107b859e0dd7d60fd1c23a4ec9390c86084c1900e9e638f5f59de9fd00798dca0d12626be540c87d634aa63636f6faa75721790e6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151a7445eb5c8f6c480e84eacfd9466a609ec58ab1f35a443e755d072ee2237ec2547f35b1de15ddbfca422f49d5587753d4b1bd80272b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4d630a91de92c9122ffa3e4769918dfcc2e45670841cfe558ad3252553416e1be41322024865fedac779d6f70128c21c9f7d5d1ab45d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbbdfb3926f5c1733e938be0b08f83617187b3a13230333e02da12c68f8b79c6716e69747df9ec5816180dabeb7abcb422433492c7db07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha522628e667cc7690e29e554bddf8c753dced4e36501f4b9480ccaff208384157dbfcdbda85be6e17503f10e268beb792b9cf07de7849b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71c6a853b729eaa2eb6dbcb29c151876cb42dc8b07344c9a0f42e35310e5a78431855e662fe23b1c702434127ba147d6101794c1182b58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he82b3731989702dd8ffc354eec4d562be2b161bfa873d6ebe005c4edeccb6c454e0f532499a7cceab34b60f27f6aaae054a166e0b1ee65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168c2b6245e2ac93e0fccfcfcb9c8426c5b87f0f740763f522fb400542938578c2d8f1927733a9e6add6798afd2b0270a172bccb782e3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1b7e275628017f6304a33460f256a942497a68cdd39db1bb370c5e7ce2665c8c95925f31468e27d3ffbfe3511fcc412cb00e9d47ffa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1efc84c91cfabb23f2d70ab522a117a43ddfa121328c0bbd824105783b09701fccbc11e05935ed4fda710e427aa068b005422c22d8a98ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf208c86611febee151ead093eb0a78fba8739c3422135789ccceafcb22a2d3cf32d86f56d101d2f7c88831011d0a40d9eb2c0d2acbaa9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d86dee9baf4bbde2b192edf9aac70310f5cf4407116381df00581d92ddb01efc17d56bf05800f1ca3e097e7a1d719ef7b3db5f7eb3dcb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199c67dd727e9e4d78604bfad78a90d8db31734f04e3cc29e4f159776a92b814d525a97eb4961af4d929e12b267f182e4bf88c9b53eb914;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188d0d483d8b7c20f4dcfe09e1c69288b92423d0a7420781a919fe75d531aeb85d0dba6987d1ba80ded68732b0aa0acd3db9a88b53162ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170b16e03367ae4f1b1c684a8cf5999f38e3e8aabe2f39a09e1f285ebe677d46db302e49685ba5314fbf41cfa0a734db73564656f694fad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5440a43dc30d2396ea8b2479c9516ff3ab11984a86766cc26508cceb491f0cdd922a3ae1ae90bf70d6baa4d3133f3206f91e0cb56b11b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38f9b9e55d812d22ce73aa03bdc3a8621dbb3c073ac1421208ff26666abe0a464496527338fff74febc9b65f1f58d935acba773023da66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a75b2b98cbe0fcc030401515298ad4a481b3b5ddd604af3009a8cd06c65b3ef37b7899c9ed12f19e7056e3f7fbd074f51dd37e45f4c49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a15051cdf4157577b7c31fb03dba22bb92144d26aa61998607314fc921a8484cafd9abce0f46b262be7b9e0d583a0bf57f0d2c4683dbdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e77f8e26467d0627c357dee941f0b1d10147b71b1fb61bba6024a0555bab495a967b7e5eece7833247c7a0d92cb784f47c97797720d96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he34b095d9454bd4e04a4bdd2ab421a15b8c500cf92a1acb71925092608591f24bc97bad693145a7aafbda700b3c6c8161fdacfb60e5f0f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h701fe1d85e08b380bd7f40f779497f3a86a6212ad7f2d7ebc7e66048791a011f8cdc9bfaeb2e82e3291f370796b59ca4a2bcb755286ae3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd16629aaa25441d8828fed4c2b96eb5418cb208ca4a03e2fc7aec30083334e8ed119d8f2546781da170c4c8509aa0b772a22d7c95f7b13;
        #1
        $finish();
    end
endmodule
