module testbench();
    reg [23:0] src0;
    reg [23:0] src1;
    reg [23:0] src2;
    reg [23:0] src3;
    reg [23:0] src4;
    reg [23:0] src5;
    reg [23:0] src6;
    reg [23:0] src7;
    reg [23:0] src8;
    reg [23:0] src9;
    reg [23:0] src10;
    reg [23:0] src11;
    reg [23:0] src12;
    reg [23:0] src13;
    reg [23:0] src14;
    reg [23:0] src15;
    reg [23:0] src16;
    reg [23:0] src17;
    reg [23:0] src18;
    reg [23:0] src19;
    reg [23:0] src20;
    reg [23:0] src21;
    reg [23:0] src22;
    reg [23:0] src23;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [28:0] srcsum;
    wire [28:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1efc946bfb47e3e35709a0aa1ba60c555671b9f9f18255f10929eda88c86ce36b47cbbb782d9e4a6bc18b4721f434748d5a0f961b23af524e37f645f3293d891ac4e7d5e7f19be12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c964b50e5cee67b576ca09cdea310e1b5e2fe290de1b629673649b88e91ece16c77f415e0f50af664caba6a4943fdb0424692a50d06b6edef83b6618ef8c61fb24bb21eab5dc01a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2c9ea9dc3fbbae728f84cd9684c18737733ea807f91035cbf4056e0e0d9259aa8954e5e00494ed38267d3f5445fece4123162776782c6bd97112478c922e38cea73230a1dc49c89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cad31d9de74d1e3e7550fb56e3667c7641832eb872de2e7a2d18e0beb3138cb38de8420935b064a26f430ecbb614e6b6fc8db3099dd6745e05269907fb7503c46842acfeb9dcb7f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb62a03099bf2a01b21c534ab9c728b26c0b104c60c9765d2be17442c3a8dfb6dd8dc1a18b66438be79589ee58dd8d4c20afe09343c52c96a902a391f6f492a2973bc1cc149fba256;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b23b24514307e04e9d56a0684bdc6a3920d0f8f3737f0332e3819148dd9229079a7c22a424167573f2ebf95008811c431fb242e32a4ae215e11c478b21ff1f625add012b9adf29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h756e5dee23ead21babbbc2f14a5dc90e2e8d642b4f441aa3353d601c5ec6cd839c59e6d7177eafeee6dda7bf4c7408592c791ef22c94007fbdb73d18a5c5ab7a2721ab398296ed94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c6beac7a5817ca536c51cc7d3ce3513042af47782376b5a365fdd0dc8ce708faffe344fe68d706728353163dd53d232ff35b44e6552ccf48931a9d190666dabc16eba4b5bc76631;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h167443e5fa2bb3fe6ce59acd1be38ecf50ae51c895343f5802ce9951939b8e3e3e61725d1809d807521c5bf81bb49e936dbb89052c985acd056fc82509e498bedae43cb4a4df7adc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf50aa11d0fa4d92450696f10865c944fd6f55e5abc63e559dc9452998e1b292d246315867e3ce6fc66e736719c3e787f357812588fb2eb9d9f03764a50a2c7d6272ea6f9544bf885;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he248b6627bf7c254fdae875e6eff589ee0aabc1e9af9c219aba2cf27d90860eb630ad5e9009904d273e72f00058e7e2722ffae796e0d671f5f5c5aba2dd64698f4cbc4dfaf85086c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d88c5249d0713b78f9f4f68a1dede04be367fd3bb1287e49c8abbb6fc32070daf4b962ace2865f441285a8a2a7a1eae5352295b2891d59f4334b295f2029ce29f244a432293b350;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b89d073d979bf5a90820b10b9dbc873aadbea880649812b29e6993426f882599b37796dcf63ce8becc2fef5f7cf88814de79bade5dd6d90a4d25ac07cdf69b2d67c97cad7da11d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b4334bdbf104eb074ee84357fa3691f151b586abd61292ce01ea775aefa327a1937bb4c203cae6a98c31356ba6f2dd1c9fba8840948f5c0a6557bafc251d3f195a4872d27724cb0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c3d07bbe39b25e1a02dc08a3a216990f2fcf1a64c7bd2524e46763748b8e84c7e68e8b6dae16212e8b68824c815c60d09784bc74be4fa36954632f4d6d7b0755cfac8f8122faf1b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e03ac2cefc8c1543b2bb52f72d2ba4d4a061628498bdc7f7d9fcfc047827735839f2191d29401855b5f81317a3f8aa4a53f7083a64957450cb9a7ac1403b31e78e5065757d905b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40d44c40ae89b3b6210e31d4a6bb75681c17f594ed646a54fca6c76b1a6add98309bbd53c6437d1e7f0f8a8cb70db37f7286ca9fa8d7375cd117c708a5e235b726632246f894e9f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6aca955ed9f778fb6f501c57eb2f4c91c963e45920d495482d40b021d77af6b8089947b020086cc70b792862a518f82283b6f70cfc62a8fb6d7215fc84dda0b864316d3654234741;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3bdbb840a085e34c258c9e29de0ca9a3b210ff75a68125911dd810482ab88a92b6bfc548407c40e3feb0c92a4dc093a26a0cf9dcdbd1900fc5764fc98e17fef8bb14beb8fa7b6fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2d99f19d8a789b08b91a87c4278de7112a3a53879ddc9a3d6c4284cfffefb66596978d043fcc56ceea24b8e35177f0caba5e0874bb241de79f8f303c2d07b01f11fea50a7018b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54678471e4b1681fb8cc53f05390f8664890b56454429c9249c9036dc520d22bb01cac67bc456254ce130ca09228fd1cde279bf9e509248f385f6fbaa309c2a69fac68d50fc0b082;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdce3fa0cab1c057ca126d168114f8a2c0086f1a5a66b45fb2397a031925ec200ba2b576003886650481a74fb545b514b766aa6dbd0c157f7b9b947b3dd369e0bd459d7f1e72e596e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaaff0930c4af084f79ccd7da242bab54a1ea50459533d79d344d1af4dc1f57af5d74648315ba3c88415d416e13c394b65be3ac02db20e4cdb1798f7e50dc7781e1228c93860f0e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a09b8c5d65c2b05b8a2292b7b1148e136b76a6942b7f2a992465616baf159b49b524f146167ff93d4be2172a7b931cd9b89ac321ca867ebe377dac13b83a279c8b91c1c6f577501;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he66b94e13d209b753dd6ab20b9aaac2274c1c430f4f80c52fd7f60cfe3e1b4506e11ccdf4bf8ee931c49c69209b0c7ed91434fb5d994ee84d56ffecf5c2585c086c123b7b217aa02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd51a731fa0c0bd9c59c8e4e8495dc8a272ea8c4699ad42163867bd955af4710fe2ab7fe66b8516833bb77b82c896fe2a642d5d868c4abe015c4ce67c02d9b7376cdb954346d70dae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c5e22ae4c3c602a7bea1dc97c762ddaf1443b82339b97110f6fb7af192c054755d78ccf91538d87d34cb40b320098229b19ad03f24ba357dfaa7bb363b4195cf17b5fb3a82a951;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5b426431a1d3abcb91425823209683ca97c60f30888686e7118a0a87873f4a52bfebc75d2097de56c75e20a9b3f7eacda2650cc5639af8b41e9b168b00d13ac443ee008fe34a055;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae5e9670f9413e389fb06771286adc325ff36face63bc0fe8234b65ab1ddf59b4c6e8f203b525da3a07966b8d94e222c493ffce93c91e2c9bbfb71a1273d230be2b7e22a272e56b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79590b3eeaeb2984016eb0aa8d768d8590faf40f38b25ace6efde5b1a1fca07e360cc0f60b3867ffebad4dff378a1f445189618dd5a2f5c9a7c6ee188af13f3f24a0a1c499376d61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h228fc341cf1e73e7482a348c993c17effbcc7fbdad6b76534d79e6b80b99b794c012b12b0e86b201167c0b47b02298922de1ec13b67ee3abd605f6cafbc7218692554333490b858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2353b0efacd67d20971700798c5663c0a8a23001328af7842534336ac743374242fb80ce2a5262bd222a3afa9cad7b24014a2312f0a5698b62ae00bea4122555b6fdb158a4856c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cca9864f38b3ccd22caefe7eb5c3f69728905b7a8ec4a0d23c598ec32cf4df000d03cf2eeacd947703f6ce3550f568aef78cd8b5d063dc9efca9137d5d7569424d9df5fdb030576;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha378a908bf78c0420fe057cb32702f103a635b636f992cfe28e2ca2267f9a47bba51a13c8a40af90c6c4d35d73aa26a87a87af78d1c5030b371e44f960fe45cf63e1a090421f1e53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a468d3e7a6e47529d342423d71faf903eaf507dc6b0ecb15c9f43125a36509f7bc84890c42e4d69b54c02151688a18d537cc6a6655aa2a65f816022da1ff574eb34f7657925b685;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63f5143361d1e0229ef0044364d74e3879ac68c45fb4c58dfb969bf8357ea970e51aa6b4fee3d952d41462bb9f7c4d24589747e776f19f831ae9859cd11cd97506b7f0d5fa8ec5d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d6f715ba5817fe6efcd88ecf531a0ae073d80d045e06546f3ce010e0e40633476051cb9e5e61524ab2b95bf15fbfc72354f58aaa4e4eb0bd2cdef61f36b6641598d3ce75c71b29f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59c064b12991b53549b538a431d1332e7fe36f854bd17a2098ef12761e0f74c5b5139565f26dfc14901c9dd24806d2f565066ecabfb131e14116856dfea5e34c9e1be79c656700cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4064e4de5d99c10e197c77d82827dc51cd3b6d2730fe56c278a85801e29dd9e04b568667888bd43c7faa39834888b07b417fa8fa82f9dbd4d0a67fa7ef72b9d144c22f99ad5e28f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0ae02ab7ebb365304419a12546a0b069baeb3178f787a8667f696d7adbfec091a595002146b4a042b8036c11e38d21a47559e63e8b107a96a591a14a46581c196a610bb77faf26d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98fde7676d14793f3f2a19eb08aec077b7f936c0f3f62ff24aed7eb74607c3d7b531e91e3c86eef5330cf69b18e0344cfbeb9e6abdc86bdb93814bf45a958640837e9662efbb24d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h144317930f06ed8e72f9046ad21c838f1a7460ecc4e075d3838579d8486084c3a39996c38f355d6d1df167336cab25fe26846bd3b2319ffe61d82cd75945562471dc5ef693d99671;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5440a5e0c676931eef7a0d3eb43f9a9eb19c651eddbc38db38dea53d659bf3da42b41aec93af6853db708ed7e79ebe2e08b96aceda0a03a95418951fd492b1a25041cda2039cc1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17dec057bf534a46a5a2dc08923794645d0de6a39ed6cf051d201b8793e6c72043cdc9ca80f7bb253e66030643e90ffcdc1a9b974361f4585930b3a3a450da84cc0b8e40af0381b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd33c78d4e8d4e5125bbc9bb886667140e8543cfdcd9f55cc28f3f1d4b92778d4355cf1382f90c6000e3de361d618590f8fdb4ef7c4efaa78395be28e1d68fdd81bf103840547176;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fe4818b7992928e615ed0b523ba045b4f1c8c8729a2985844a7b54bdf334b94aac985d8a0f91b424a2a092d97ece8c47a446a12310090327ba2bf60fcaa0c550ed094929b00fe2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc46fe32b9e96e9f80ed6415a70506b252084bc681228d0ae269d1dc55ce69714ca8f6a1f7f20f73a38093d95b2f843de6230a9cdaf3100ffd34b5a2afdc33339882ed807b2b06360;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab60373cf65b0700982351a0934e413bd252f443304f310dc4e79a9c0d722f9c8c3a220969601e9dd89896dae3d8bdf23da8d0b23ded3611896af5c8bf101135f4ef43a5602efac3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87ef371f79bad0d4ebf8e69b93b204e3925ae232e46507bd87d3c71cb52cdf97e9d039b131f9fd7c649f80e7cc02a30f116d9caeb7126106890414e35615c08d28975d2cbb9211cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4081889985b20d31cf1cbe1379d11a7464541b6af41659ab7a554789b73aafaa95379e0cce3aaf3a3e58bc59d10d9d8a35ea76eb0c45fcccd62e408c61c09777b4cddb0432bf913;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cffb9755f231bb81187230f57c0dea0389d3a2a5c97b59ce00d70df991dd24cbb00770a7a0b8618200ac3b163c01adb1ccd629fb9fe2a6ec870276eb6ec23ae6515891d0fcb6515;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbcbffc77f59172129aa737d7833b5d6396c35de2a49fae4c6d3d248f0d82e156dbf1c3354c925323a99963b715209c8142edbd0908d13a32d47ec2af2c02d5dc59e8156c9726e6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3311c4be1ac3090b542be6756775cd0c2b815da5677e5808d92d79cc4eec9d4388b0ea5db197cafa9730c843b55c1264d818d8c49fd502e4cb3120625c65527d4ef1f00ed27babad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a09e83c2a865ac1071a9e42fd7b06ed7e6d8cd485fe5c7c9311ec8fcdae431e5fdb613bdd9eaf44d2d27ee91d3d0950290a14734ca1583b387d87f7d7ca82535b7e470e23c0207;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb55b275821b51e69a32654fe36ce3b6a89d25f6e6207d05663e0ca36b14e576e06b5684aeb3b8aa03aff0b030ea6e05f0f7c9615eff817802b1875ca137c9b830c5a41357f17d08d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6299c9e6fdf02c4c1fdad8066b421cc9aeaf7b28cf7e348f35f336bbf4e6e65a55281afe90fafab54072a51d426f2fe52675f60449aacb324886633d4bea1d80f2df8eea90de48dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42658fc3b6009fd88adc18fc9992db333cc7f86092d79eb544be77bc66ab07a9c09c18903ea707a230acaf3ada5088dd012176bfdb375dc0dbf73c1cf5a6a555b787ad950133a3f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e54ebdc0fc736895f3a4a5fc8b614a0483dacd7328923fed1bd57722f30bc3af8cdd0d32035bdada68b31da551cdd70fe07ab0feb7a83339af3424be431661134e34aac9a1d7448;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3cecca05769aae90fca98a682b0fcbd718c97ed956e9409ba8aa5c3afc608a05bea69854cbb74f184ad6b33eb20e15b19303340a1f8b344b3d77a8ee05445bbc23b0672ebc077cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb588c860666f23d439f66794b644de88764546ede2228001f1cafacfe435807df63a9a3e9d2fadfff9db7bc287d1727d713ef980ebf10706e24c213e8b54ba0cbe78a43405e0442b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b789dfa5ef9eab834c83774542ccd68aec5b12f9c5f535fa11b6a828f9fff35bc6651b6096994fd12bf6266b61477d86d127c2d76d2421ae3176053f7b70c82bdd28af45d13da1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5a3cc21ca68ded9d908093ba4cb793ed75a9420c4875b56ab75e6a19ccf381df7a5689193cb1d665eb304cec2bec65f50d0d27aba26b79cfe7dbe742892a04d74b84d377640eeda;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d395e47965c958088ac76007d902a0990deb2ad0a0125f21f037ab77a69f7683f0dff57841d5ef7d4d80a2395bf07c1aa53b142bac41265c85733c57ac123488fa24d17347ab7e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5b78ba7e1de55ed49b8bc2053f9b799591c4c96b8c7385543a27b9b70dd3c74bcd0fb2f56bff5e7263e17d853912b019890ef0829cd62ba8213783be964e12f8df401be4dab240e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbad0a62857773e7c5f8b348b314aa9db3cdfd9f6d0c169f7f307af23e311739118df70dfb698dfc8a6df84864155aaa8d177ba5be8ed86bbbd2cb7fe636080a02940f0bfbb83ca5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2c2b76c72904ca27f1ba56342e2482848cac8cef541e253d275d752579007cb29fcdfb861d80816f670ceb91b2b6acda7b8502b0f3ed47696472ddea87375e1b45768b419c1d199;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb150d14c963e17009e5c03ada4fa234364841c1dc03af4fa2d0cc1cf8d2f09e4528c427ce028ab8cdc1bda47ec1a6d453157afa5508dc70c58a5f6f6f431536c1776c58c316c9bfd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3468b1ec5c724dfcf60fa28e3f10a2de4d17ca1b6398e7a481afaa7a423ea963c97284d1aea6d151624fc16bba32b131499e927180707ef4bc6b3fa1ed838d10c53176c10482249;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6692a2af1a40990d038790200d4f5198f345adb0cf11a267f1787eec115ae111887f30e717f77dfebab602f235b8e6cd918d6986db2459c94f1cde67db822eba53dce020da7e634c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf14aded3a46d5bbae16d3dc0943a9c7c777ab56eb2e3cb4c076382b999c040f3087a1ec16c9379fc90f0d698cd0bdbe7a2e57724ac0f6be023aa0645458b37c5adb32188e7d3e4b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd5294be48d10eff6144bd8a449d6c060f21d9574b22765e83ec4eedfb6b9236ac94a8fbddc117a6528de0ce9d56c563e3d81faaad5f3851aa0a98ccf3fc5cea966c036a90ea51db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h442840b4f87c44931b17a2779e97655d0173bb716f58000428fe9998fa131e5e6b2c077e7c4b699430ad51f9f236fea9823e8fe8f9452f57404716ba05ff4d9aee47249bc41c6bbc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h877fdfbe202f9e060e3631664f10005fcbc80fb79dc7968ee3f89848ac5051d614d42c807a5744ba1c7ba03c53613ef714f6f78c0b14f9417289580934a1321e5b7b41126b945f5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb664b98b5e8a06d43124e57a8dd458c9ec94b5df375f82e9cf66e4f60e58137fe11868e417cf77ce8a99e9c713ac6c3d33a462d08323428f6b47262044ac28c69bdf72f2f6c5f65f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h763839278e465e505f3f30f5e2791a17551bdca06969c617a5b2406308564bcc6a9d7008dbbef917785c519d4c399090750e3a328b04cbe110d18bb58e99542b9d6f99bac3c410e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8789698e3b7d9f69cf15dff3c060fa3f2ca531767c8aa467c05f6822bb91bf832ac8875d4fa618d102d763ea8fa2227e9bf0d460f1700458095307c29f4360a4d6ce2d9a3e8500f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h919a45fd0a3919e15bc504e6ff8c8ec8007b0a7800eb14efb59e5f46201d3b12ae1301cb2790ad7f61b9306a508c43c2c2dc11d5f3452a48dc3760a7886b009763d4c68c8988877e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8358e346cd8d1ac97bf7559e94b9cc9e2424ad62005f3498ef7841116493f089ca198a4492872b6ba830fc36db1125dbcb18cc67d1d4a7d82f5a81430dd7f66148b36465789a187d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c694f2a1d2bdb90fe42af8fcd3c22e339d1e0011535a7beb74c6dc2083682bb50bdcb1b0f584a67590649833ce7f987cedfd0148d714ab8977013538f9b82ca92b28abee1185263;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96534e7a0f614322ded6e471f9bb9b0d7bf27db22f72cbc5a3ef5ba224179eb75777e5b40477b1560a8439addb9cd5b4d0e06638c24a93b5d9dc93b2565ce585f28e55296d4dad39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7895b2f0b5ca0b3850920092f8ba1db39cae0af7dd1b3a338e92650ee740f4e632082f0e89f90e1a4c2cfffb08ce055ea5265e23dbefb9fe51f6ad1224fa21eb5bd28d1f33202c07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdbd3d0819b584935cbdd0725689a3e39ae0847cd187d23917be85dd3adab5472afa008923ed7f73519c2ae1e3b1f5206c3509fc26ce1c04773eb32da72d8eb63c0b878fd696253f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ddbebcff41a550ce7710627e195b930ea13bcae275acbaf5f3ce7e3d6c88e34cb2182adbec495c3b9053183e22f85f4d6d361b137e3e1d10ad2f8e1dd81cb97a3b404058ef80da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a97270bab3fd2797ce945c3d17bd3aa59ee827f7bfd7cfabaa148d2b3702390d92bcd5d8ab591eafeb289ebcf952bb54932847dd6640dff507eba2a5e296cdd188cbee4c1bb770;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfc7442d2d0d67e1ea1ea9243dcd03c9762417e828630490badd9b14300f1ed4639854bd617daf9fe18eddf51a646c62f6db53cac36d2eb1e3ec227bdd12f8aaecc0dfef34ed0877;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc57483972a83e44d34108527012550d4f1a9861d7852700eb16e5c403eb9fec765a611dbe1c8ffbb61dcd5ac45250ceb7b744a3fc0ee36beee2abc108659b1b31548320476c9abc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a630efdbc744ccd282dd895c6b15e83da56ed3432a4bfd0f162e24956de85cd1a18f676e7ebd8f444580ff98b95f42a5e4ef1d849bbc0ef9e1fbebda83f3ab25a8cad91c22bb62b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99be9ab2cf6a61d558e4f6cbaee530beb57a7cbdcb77964186bdd91a6ac6440cb8557eee7d0e93283df71e48a1f80138c2178355088f65453a709ebaa8b2d6b2e312d5bf2dfeb5a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2b8b4cb0ca029f5091fc068ce563f5c4b6e704de11b3f540338e53b54a3bf54a42a691a48b6c7be0ac89a0d12f3e0906e1415daa6d28a1938d1b7b691a650dbdfe02b1fa97af51e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7e19826cfcec41d3d8a486336e61d77621e3a60efb3e7222e661021641a81c66318e8e05d2c3345f6afac4aae2182210e15e6feac9bf6aa4144e85215b54728151a2df5d26380a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0e99adc12b5ad91af4596c6981a5597e939b3e16871d9595337faa371781f6d50381496ad9399ef85e491f4cbe96ce2baa8862144fdf27f0b79f9f5686a8d254ac6a0b862215717;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he793076992ddcbb3041c7b48a33a1c867b48fa3b3475d78e8e6bc87b908ee193af2fd655c0e99f4d7648cf822a5413d512209ed2a1121b9925704987f9707bad8b4d1da702d8a7fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63551bd725295ab4c63d9175134594306d281ca7014912227f8474e924fa4e071523de6d16c6708051ae2b2d541ff25a67df8a6b9896fcd715aae74d751ddaaa16c9172c7f0a1e61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2fddb0691f5bdc8d6194384655e6017745331f3035eee1dea307f7e5a954ec8cb2fd7743b23ceae8b40996efe1b86d1ddb5cb8452f006980830f325475707e63ae3e50cf336d1e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacb2cf5e76eb13ea614925018499ac9b2e292ba6658edf0d51825b580edf65218ec6fa88521032e8d5c9a7c3f509184b57e5f73164b1630f42c750a7e25e91d7c8cb4fc9fddcb239;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15a72fa4de1e40e725960b189e6e72e4d78463f8c65c534465218fb852afb6c57578a91b31d85953d0cf8985e77e35a3e6d495d274a63d82cd54e26e781941e221829dafbd8626ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4185840d66595f34fbdfa920bcb9e71882a73f81158c9099891bf105f88c22adde792abd1582ee4ccd2d0da0aa3d1001669e1483bfe4f6195af2875fcabe817904ef4da0750acf2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4c2befeecf44ed6eb15ba1374c07a106eca459134c7f588fd8944808540c6386c882a14bd6bc0ce5dd1a959789fa18300acb892bfad234658c258c6fdc8c582954aac31d365415d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c48e8fa02836655eb6aa510f2ccfaf22e0409652a5653a028668bbf472fb1f5455261e4f2c16e2c208e36c2ea0efb73b66a9fc6251c93601698a1e2321044b952abbb3625d8338c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ecfccfdaa5499179b2b65609ee4245f48d8aed2064d03fc5edabe829ac9eefdcfbf3a75f691496b9be489b568eb4ad455daabe6dbb64ea799420dd8f6705f04254fc120cf79ccf8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cdba5606728788fc8b40f1b8545bdf4ed2c79f6d7e6417144e244d522f027eb520c0e4b5846c5fc512f0d136bc14753c93311ca53903f67cbd18ca025a56b533a479815d5bffffd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f338c529cd30ee1470e6011760c256fe5319fd884f1a2425d0af5f6fe5bd290faed113669a0f8741122dde414cfaea4a54c57bc750a56adf074432c8e622eb7234f739391455e96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f57e72113ca2a425a34bcf3249b347f4d9e6973268b55f76494d8be7646cc6fd1ea43f99d27d81bdeef5df5145e490307bc337c567fa3a911f2b0c9e08acdf71254cfe6f04f4774;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cb593cccc16b1279f7de323a52cab3ac4e75261ff275238bf6f015fd0e654e2619c955ef72c02e5d8248391127d645c6bd79bf73fb44e8740cff026b2b15e392faa7a05d9996f76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a6d47dd5afc1fcf509ab5ab40e788bc182ab11721d6b123ab34648ba9198bada3f554fabdea4885128ec2e5985e1581c1cc06c120fdd105cb55fe8d39ffa64ef2b2974e07e43561;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a44de6af1c7fc188524f70ddd16b01ba2a6b7132ad630f446175e2a5bb2fd9dfd84888f9e9353453af45e646b9ac33033343bf39968d4953c6a2931b861f154c282abc0270f5dd0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd24bb79166be73c5d36119ee56f1c9dae952ca0a4f018af9d6e460423a532367bfaee08cd37ad7e731c90ab339f816ec1aaf3bfd78ae599b890e1d82264e8e8a89afe992f333897;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1222747a9d6804976cf340e1fb493f40c09e7d6fe813788d11dde255b2189c9d52a31cc647a5190c3499ae51fab1886d1521e4fd8de2122d2a2dc42ee3df69303113de6be6d8ed72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f4a63974aacc90a8eac3b90b51f42bfcc034b78f7574e2e748ed039a5d2da2c1b2dd7365758002ad1ffb360abc48d369f81a951aef61f682885b7c4be7f60ccb1f32a5984d4aa21;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56e68d5bcbf15b818fa156c757e74babb529f88f6edded190bf2fa40d50df8a54907bb8591fd6275e6bff0a753161fc731f88cc31da1ce6992c9e78c69a204e39e1593a3096b88f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a38af4704d047d5e1f7b8fe19d2ae5f3382f250352685501bd97fc3553d40761e08fa72f4f02e08a61c1910068ce1cd0cf7f41f155cd8ec4b5a6a2b3616893e1b267ce694b3072e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e03f8875c5d0930171e6888b6eb1a82a8a292e572cf35d9573c3b5fd2eec215b6a2054130aa476a5d501afc254db0a45fa26f47a9e7b37ad762bb566c05bb049fd88f583737d186;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9fce88337a5bd978867f0abe695c73b1eea13000c2c8fffa24453d72e3a14e0e4704915c45e495c3d8030c8d1ebc53cba4953c777b4360f556078e268d2f0d76b20e2482fdcf5d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45b84b9f855b27eaf670b2ea8f12fcc002aeb592da3b1e48fe96254628f0eb4a15823c89387949ec8335915d21fba65af59bb1ab2a997a1b152cd49bfebeaf565bae4cf2b2e8ed85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha733e9456cf7f571a86022828191afd0db1616c6c30d9a9b7e8ed3b87431b3d96b8b480b20ed124f48983bf3915e451007c6550968fec32819009fb5a947a5d68dd2c0cec1605fe9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e1371c59b39bd0690a2cd703c48a1b3ceed9ecc328f5d0c5d326408815ed6135250c994c55c56cbfe9acc9ee2faa33c30b2266038e90ded3c4c2d482e7f0ec6e4839f60ba0784d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd53752305f87ece450ba090191ef0eeb1a4fe88645b9e40479e69f2e91518ffc9fddf9b3a8ddf49add9e2f6b54de29ef205de814fe0cb1ac385345cde8efe671f0990f9cd16e41bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdafd071078eeba42c81fc2f552c69bb0f4aaffd18dc21ff713bb1d2404cc2521175643a62fb6bc6ef48897a64063d1d6235e98a659e26ecb3c3ba6d7c7435cee49d5c43ea8fd7aab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha27e46adc1012ab1033d9bc5d83bfa05707f970052d8953aa42d1c7d373f5b2c4f0e5756edddab69e4606bc2e0c83534376c5461a39bfbee51368be8fcf62044f3e132fc5b464793;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60a3c1424c2e06a2833a0089b14c4e7752b0323357c680419b85ec5af7ad199bde31790d214018e01a412ecdca051f3b7152ee73f5b6d03fb0f5a1dba5d8f23100aecf2e8e625a84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4ca7217f66ee7e42920869819d6a6a13587668861a3e249585e8715080ce3ed3c4c3039f140798216ac0e7af81360b3b7e8abe2ce460a0dce566f72a8ec911bb32fb7276d115bd1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d2bc12d9ddb1003da4aef08a7b5a5587fcf33408376373ff3d539e2ef25f06017728fd418f02ce96900aa86edd879e8edfd09b610394d12f2ce974f0814a1a501932b1e2e2b358a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he690a84e08345d0736259f11a088972cd5574c9f4c183fd7519d2478ab3dd4063d321e70d48babb0e85ed761aa032ae30c3384796077f5c281f56a304d58815f595936acf882ee48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fb0d58c6889eb74063afe77dcf3a6a107a373ca67d283b7da0e1b82314bd89a1df3c8e9335a438e18e05251914406e0214d831734c126374f5c19c75fe1c26a2ad950517cdd6961;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h557da63a24ee35ee916a8b1ee4ab10632dda6489863c72e40f73f87260433b4995b250d2b668912613baafaef81f652550ccee0bf895c5af9c4a1d7f8f3ca5014f295aac909b97cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a600f25140ba813616d75442ad47a03e56fc42ec144ce1d22b98ab74ec33a68bb693d211ebac06f0f3a5611e0634da32335608c153714b3fb8459cce42fe720ed98d48b88186cb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cd960f4533d4a745d03965de42ac582706100bb7ce9d956523225a1e284ec0dda451d7a4eb46c1d859ef6e9e804f0ec21abbbc2e207fb006568bc09f65fe6985261896572a51d81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59a226b5a74b49e7299e3d983a22a58252d749b02cc5b26d89b0cd202a0debdd0a6f6adfa6c302bc63f11cf145e7083bb4dd27572e9b7114529f2489dd9e57bbea91249e73f75a6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1e559aa20fb4a47c943a0cb8eb0b34ce1a49405e884b3328e182f8a6cbce0cce535b2f1cef212f425a560bfe1942df6cf88863f8aaad221b87d658fcbc9afd5ad01a718b510d7dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99fc5fe0c1b52d7fe03bd1cac725497b3b2e8fcdc45fba2d83e0c01b8c6c0bda629ea9aee3846f9989c7f08c34f8e24f2ee23b2dde7681703812d6c4627cfc0e0537dfa24eede3b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61dad77f628a4b2ae42bfe8976ea659ef7c7c26da8a5b8e756166a4690402ed8290e151f4082d78350f00c5d75ee46ed436f3c728f397dd3bc675d33be38e923882b928d69e25729;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f78317565e9d2565698e9af5a2039a85795034f5e14a018b42572936403eecefbcacce745f2a593402333739fa9f0fdac7c11ea7c3f4de7d233685fb9c7580b5b55dde4e3710f4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha47136bdb34bc5a6d9853071727e41c67083a75fa162a85329534d0ea535be8652eaa57b6968443b71a08b8c5bc6b6af87d0767179703abe904f9017168029343e8c6bfebc4a0548;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e673246754d2db38d8df5ea852c104b89eba6642a524dcc7ae329381a40b0ef8755d7390e357c60e5fa0be9af6c9f925c7d251fba54cda6a5ea6e7d71dcda2a66f30a768c912fc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae12d8332e30bf6e0d80bcb704667604b6233104c3a9ca6fd43806e667ed820c3c483e3680721f92a01515781616c568d6794e47adda08e48dfb741c4e0ef7b36b18d7b5ba6e6f64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd96ac0e60d294a7c5d3cd0b9158ccdd0a91840a759c9372cb547945a9ea6fb45938e08f1d1b527fecb7c1c1878bd784ffd243dea56663b6c6a5434fca7f70f7bdbaf45a017375d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd030035102710b037beb33d8e104de8dea39b1d930c43c9f2202e6c4b4ce453ed7a3c908749934afcdfc275cf9883f292241e3218cf570f61f792f1a2f3bbf7bd08f79c55774f752;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6a24a1ba7a99498c8930b81522559d43e37d46f744813f1901a424342f1a93f24a43d475ea901510c1a21349b7da3cc265493e07e8fabea8e18332128f5b0849acb4c2d68e7bc3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f94415115f307db29386a5cbd78712e2473f4b303a0ebeab86861419ecb83957d68072276a4c8daaf9bacc8a553a86d33204335f96dc1e5dfd5e7aee1dbe0b68b699865d0ef63ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfca7cb7ed14591a5032edf27dee99fb5829421890f72c45e352c7ae701e36bcc103f3d2e41bf46a5e9951fefbc74e202888d141fe928ba33d7f50d70298f83a6fafd09726ba2e374;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4fce1f7fae93d6fd34397ed8210b6099b0fe2017ccc21fa6ee4e9da222d2abba6db8680fb995a774a3091a56f785004fea2c8e3411c11ab7497bd26d526f69fa2c796600e87cb7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h325034f9670ae1f574e83cbd44cd9e6afa42d7ea07e622e1c25ba333f0af8b52b0bb60bb20d66f6af456b36372be2e9c78e3491ddd603b2fc8dcde58d6b5386079ebbc39fe717870;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h685e0c0dcbdfc2f640ddf9302b7c45480131abd4eef8e143df5beabb8fcfe06635782d2be9918f1cdc2d54a5fc106d3d95ff659cb3fe0f51461171bea77f05363329f351c5aa10c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb91d71b06721e345916128222d6e995a6db60677881c6a060509c2974ef3242e59055a5878fac7c56d06ca90576260774203f3da3b7660b1e416c1bf8560ba001a65e8462133e48c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9bc72509dfd580de52797315378b85053c7f4004ebab7f2b38fc300f1a6ef7cb39f90f9c05bd618b7eeeacaeef9c50f534e3912ea1c5130d0e251e9d711c9f03e6e63288ab37941;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba137f13a6c6612ff429fb32ceaa9d309d9234183f9d56c80e770025bd81e29256cc23108c09128f3f807529a002a0b50e91a12ec1f14730c0355df971c54b31a288cf97650ff587;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e630ae14d6d954710b680b0e45cb90e181c5beb0d78b148cf6f7d951073a83b9f7f837e2f018b89818ee06d45ec044de530bfa3b7d689665d85c9833519043ac4fc9674b65c32c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7ff0a2aa49add7ee138bc3bfb031c47bd88d0984dd60e72c215c2b7d6f8c093af23d07f3431d355f2324aad41c8e37b1785e98bf6e319563a3e0c95f63bf71d18f2c32eed70c7ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27b2c57eef6a52a36d067cfed342b8520ed4895a2a5a43d69fce01657e14c5e1313d6afe2faa84f0b578de9cb8aac939c864923d3e166bbf95533df6ad22ad4994650008696acf31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfe804f0c51b751788f3e5c53b74e7205bd40b2cf8b883d1656b8d5683cdb626faace4d6bf3ab7a2ba82190bb27d53cc4509996e0f583f90b2f0b0ae0e594634a93082168ba899f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff7c710d438f0b70729bc95d66aab1246840de5b39d2dd33cb8ee8bb193c35528160dd5712c4aad8c4e201f95880aebd61eb7331a0ff327ffd30db4e0d7d937bfc40980b158d0425;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2022b8e606c7543f2f68daa1a434f3372c836c6fa272a789ab9030fb92b3c640a86b225ba85f1f57a0cc8ea0ef98d30cd432019189f9e86f9899843358d77955b57fc12c98080fca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h231714273e5b94b0b05a38e426f872c0a3d33ab1da57bd4395242b89e639aea08c26420956c51e8950906fb9de66cb0459f6177d019ab52bfd493b377f33a904f2d52485017e0800;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccbe6e317586407ebd3e1d408c1ef25ee4625206a9d5633ee5741a09dba956aceb1049ae36d6d16e41b1d4061b3c5adb1d9b243e5267fb61504a981e9573d06bdc5774ea80a6666b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ec8a182e69291563bb4f803070c3687ac4083e513ee1f37eeed3a85e5d03d1b14c8a9323104a2d9886915e0c1cdf58de65947bc85357778414f3a95c6915fe69b607ca36284ae98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34f49d96e92364d66900e23c383595ceec6d591663541a655a0f1bbba991fb4eb4911f3203ee50a6c7b3b2e04beaa21471bc0735457dd0a8aad7f1acc199cbaa6bc7248ad326c5a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85199e0d35dd615eca77ba6426ee94915d88a360a1c3c22484604c6c61d908f61dd904170d2f8ea1ccb207d89a3776b81f5e963af56d10bac4cb765f9c1780d1e813dad43ee5ddbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf845a3f3fcc7f2ab6e5711628d45270f78f18b9a7d89078047db1dd91ba3a4eea58f7c4f37ea020d9eb064c4e3e9323d5c2c7b7ccf6e355e9e3f66bc308d5c7eea522b6835ddd38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9a2450bad0265726b9b4d7a3111c02db268a5a74fa4791439c1fbe57375758fa7714e32145c795980c4bd1bdba36f9a37becbe0286b9f4a2ad019d1650f116be35513cebe7fc0df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a330583617bc850c19059a41dbc06a6236b7e097f4dfa77f9e84d551f9a4ab2b51e5c46d1fdb6700445183051e1cb55ab914c6852ab59e763b9ec48cdde385cbf2da1bd9a312c10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff12863e36272b8ddbc7e7df18c8439c9be2ee10a8db7fcd7fbfd3b12037497b60fd2e0bae5ec761b61b627cb3ceb55173d78f72a176b7c8dfa6d0229dc691dc046f02b5e0a63af6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h537884b46b14446fb1cc9aaccb0ad0af52259260c7aeba6b99ce05b21141bd447f0e7a836ad5b69cccd0b0ac99b76f1b6d943a83e94473f4ed595e842e5a9d8419a392bc429ef8b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c6ca443d8c2429c6614e743a058cb89fdcca3e3f1d2fcb37824fd9d4fc97d3a25c7f77307912ff0eb33a9d9bfbefc567aad53e7879bd77f4c40c0e1f27b30b75999d29d39c5c131;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb3ac2632d3fa3a93bc37fc0b361775d8e6acc3620c8a801b75cde82adbbef01fe649559125289dceaf7a188578a06287566b110ead0fe7dfd9e0a0582c91b89695f8f9084dab48d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c5891f42534b1f9549f9bd9ff8eba9a367d02bff51f6122b4632ea4000cd0e9ae1808298e998c5ffe83c97955b5eb5fe802844c87cad34fee0a3f59f6b5a90337ad6b75fbe7f21b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a17c210a8762061c6b1659c25ba9047432a67dbe68762e02f2fd2e6292f0381e1563b4bb5117bb09ad493810f39db85c61e67afd4667cde66364bc7bf8b47e216c0b078f0c5e0c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc79e5eda8a6d957ad5de4847f8b59889df3821e9059a1e18c18cffa7d258b77c4d420cd4f7ccb8cfab47e0159c8848cfe6e2b77204708265f409f5c0169a3d4908770b20e70055b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59fe852a177329c2198c1828e378e177ccdf34507046494c76ad364f2d5374826c1606c41e424504ac4cf12e2fbde56e246c2fa17a735b5fcb82a414018025ab9c421de683b01ddf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab62e6e7307ba9d19ec286ded43f4e7c13a50f98d720059828bbe3d24694d78cebee70ed5dceac232eff8e88074bdfd1bf6873ea3e4748db77f49e62919b8f9f201b796b011aeb16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc22b7f957a2e861d53a9187ec41179127a10f3f066a4721634119bce807fb37522cb74bf870fee2184fa9b163e8a1680e801594aab024f15d0385d00cf3a7da2a52d87b932b467c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7898e48d4f67404b0b9b06be2449207df1b2f9c3ee412b45b5fe06926846744f41e3723b906d0266f780267f8b7165f8aedaa336243cfdc83b21217455b3349f2cc0f1972a2ff79b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5e95d7536bdb38e8f93fda6c0699b06a9f8ea4f21b51785c183fc9f89a8b1e5ba006e70fb8d94524ab55c0fb365a21a9e77a9d6018a25063126a2f37c9dd21282fdff2afdc8d9a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ffe5cedcb844cfdecf0b015a2a8f4071818357e2b4e963b59b2bd65594391fc2e671835f9dc0cab87d2bb1dcef7596c0a85f1c7699889c28200237f522dbdbebf9d9b6c2f036a8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf5803f81377569db7850ec9eddbc7a3d4b93a6c42b1ca071dd5c3318d1efda0c4fe55d6a84764bd5c4f33b7f10dd554a9081f2260be12c1f0e64bc36fef3c1e10b5ade4a047b89d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b523466466e3f94d56c499a84002588922b677882c0df6e5d715736ff59af21a6098af2996092fd76182cc903c87b7aa0b385720e98303b72614e8fd2983e5f9e90f14b3f17ae74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc5f9501f730c09d8d941b51050d1e7a7794ee43b24a047fb822d01ea079bd8c7d832e31c349d5cb26a13190dca825841547a4b5e6416ae4ab2042020f6ecc0d770d9da2ba534e12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h395fe6ba31256d78f66d13cff0a10fcaaff7d72d0e8aa2d85ccbff8420b7e873f4a733b8bd611f80256b1d60aa1c4d551d132ec6f1fa51aad87b7ec703a2f20f3690f9db0ba9bceb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee2331de6795109a6645e8037e45372fd042c30cd44d0e64f5ed4a7e863dc16c36870466d781866447e4e03f09261da9cbab9babc8ef6281e29540b2d3837cde976bdf1909dd3aa2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h675d99f39ca1456c8e41a28433b9d1bba4b774ef1ab77131d2cdbe5f14008327509c17ce0b3575dfaec0b40126da489ee3d848b3651c62be45e7a604591255ba506327a4bb20d562;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8472024aac3c095beb7bf4c81a4977a44315430bfafddcc084ed323c7485a5ad26d37a38424db3dde612338c944cafaa6902549c0749cdf109eb79d66aabd2046013cbbd22c0c35e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64e9012b00664c775a80318751bd50dd1e217c4aabf728a775c7c4c3cbc0a20a9f2ab520c6ef0da8f6511c80521796bafbf2c3afc74cecfb9637369ff23473460df97040791f00d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc651e01551dbdfa0160ad019d8a366d60b6d8a0696e2f34aceb8daeb621ff452f454947cbfa8506975f93f8a2f055ac9ce66faecd32f263b73fe7b22b148ca38147fe2f866b26b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f2b21aaed8cd86ee0fd10498f4e5d27d58c834b9521843a965ac29f6f34adb167f100e7d91333abe553032ecc195cddfc06006a17e2a511ac6dd4fade45550e8d29496cde0feb2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha781211fe79d523ac87ee8a67edc1987b75d38a9d0d259a4da8fe232cd8419523efd8c4dee0e48180492bcf638148c57b48c01b7761685fbb88dc0a1c7b8559c1c79140bf4b6f9af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7642f60c4ae5d5b8bd1e329ccba8021bd73c3b0fc5cc2d262c84066a00e2aaf54152424fdacac08c97ded4f2a1abd459a0c25dcea93a7e9e8defcd95f5d3ea22db9b29f87432c372;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8343fb092bbb249f6bcb322368c6f7c5d28639576f9a2127222877b34ba8c168d20771596f6878f31a1af7e016e939632c8e2c7bd669effce06e750c9b9056b9529134f8aa30231;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c7c88c8e16f71d4e48bf6bd68aedbc33282af5950adb960dc9336bdc8f28ddffe9cf13dff1d7e2c22496175251f8a363f8ac09b3ac7a8153d940f8efefd8fcc6d316d7e6b30453;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8f3fceebc31bdad0420fb20c901b9240ed70a52b5b45cc4122dc43e7cc0d4510b05dcd29790d77b35a1c70beb03d3c2acf8430a816af22e6f9ea308dc40f07e0422e82fd0dc86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd609cdfa0ad932d2c4fc213d4e5c1ac36f2bfff5007fec708c6aae393cea60c1ada1eb2473135d067d85c9f460e9d5fd3427369de50dac1e8ae54e666e20e0e14d19b8bb15444477;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b60889a7e63d93d8f25750b510762d43fb6b44f471bb9e118c68c16bcafc4b643c487ee63fdf8b3e530901347f9fe98ac50aa6e1d2af8ba5d0e970a4aa9e65c740bea8dc91d54eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48bac92a065a91f8c199c090db63974d389b71317bf4fcf71af11b54bd1b54212d37039582ab8511d897ae687a2c7ea0c26710471f6be061ec9ba4f6a10a220b5e0654c24e1ca643;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a848e7d1ad718c62c75882587394e5f82b0905c4edf0303d9b7b557d13bcd8769f803e387215e5bae20c05a97defc0475f34edc52f21c79146ac20e53e612a098ca2975ddb5bd03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7398340059c5c839f65de8381d4eae29f10ff4bea8ba707196d6066dccadd96791afbbb01bfe22a44651e1c5a7d7b3791c39c037aaa57e37d9cb294e60943ac1d85519815d38ff4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h655ab01a77e518bf82ad7a05d8db8879721a86db114cfb58744da93ab167f6b0462ee0d335910fe4ac575ccd2f49283e99bc14bf05477d1698007aaecf27bb6d58a2e617df28bd8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h389c8af61af003c540dfa8c6c9da950bb293835c84bceb3fda1b620520dde876cec5bca267a288a189eb73e50a933665e037edb40b5135ea62f9e87f3763c74ccc61c819f2ea7cf5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e86f808c93df24b367ed7f0dc75a36e0f2857f9ae3a03644563308ff05c5cab5b33df1bbc4880d656651ca4f1cb233a0d930c49551bb52facaa8efd915cf04ef477918d23578a50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52292d0f9ce28c34ff80aca068ae3195c0f263aa756ce9dd84748de7801656118e41d18003547511dd1adf08ea56921b67c587b21c289e75cb0d8d739650b73d8b5771e7464ec03d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80eda63e92cd151c4690476d5174f8480ad0ea4fbb7a3b2300a0225d75d746972628a7f469062f25c0883768137027ead048f60883002f9aba38d0a5c45c734db372ca2642b9f17c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e6c4c4d891e1f97d2a4d6214f935564bf04c39ce469a9883c5ae93610a6da00781b1c2c99890a914ce10ebe2c381d9cd5565d2aa25a7b7eb636b64e5c284f722bcafff6c234280e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb60735227329b9885af7d6ff04d895ba3f1e290c4afb113f5df46ce73d0a2070cd3a06a3a551636e551fb9fb9174e56873fb238122360a90d2e0e87d3d16d5381560182c004dc79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7425812073cedc093c2578ef623ff2bfae531a99f4a7c9d357d1f9eec9d5922ad66f69dbb742503faa7aa89049f4a04ff185fa34fcc0856d8ec66b074af620101853d30f923a390;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef225704084348c8c08acd56caa5b214c808ddf6c49f3858a3ba0810c0d2a01ff6e80f251be6b1ca7f11e98f9109a6d546ddde6b081663958d48d683a39ab4e9e7ed0e1d4eb5f354;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ed6940b14a58cfa54065407d985a6527eebe1154accdd6d3f83e29c94ce1660dd592552adba3a12c3a48a82e0b6e4efc44eaa602108e1de74633699a3bf72dc5f751f4ce60faa54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd289f82ed2d54eba1d13b7bb9934e47b89b4cb835f92ee88ece4884c97b97257e57274fd9d444360caf194a0fecaef1f1f79bed43419dfae830414a14a0b03f1d8facb39e62eefc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829c1ad449e987a0e3621f9b05f405be22eb0ef7630d2bacb18501042468d80d802bd2ad631b631a5b83ae6c5d5ca37e3b812dbd3891b0914cb06ddb67a86db9e726177b3f1b3d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ad23b42224904308edc26180e790b5b021df96cd75b40b1698987df27a5461c7bb08be761f23af7ee7541d13d92e940bb99266cb626222f44fee20fb6869be7a04d05ca7d60f27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc1a706e70781a3fda7ab714b7ae6b2071dbe2b3b612388a9c02b25b73ba9a453fe9d81932477982fac6eaea7ae086164a5713ecbb4c36df2a99018d03d64a33700f5464ea4ef895;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2c48a1088ed8c38da4bc93569e953db783e6e76e5033bc7980b36dd3babbbb749d7b38f1e22b4c26ab67c0d7ee870789cfe656d083c4b70fe4b1dfa33a8d4b502b13d07e0a835b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd7e158419eb22b27b53b7dff953bd0d5eb1a88f6816d08d17355facf9a7ac1baab1155b84e890ecc3c17e5ff1f08fb0301eb611598d77ddcf9d5b07e55f34fbbeddd926b4720fd8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4616e2e6c0f1534891e5cad249bdf00f1b271e629903b36e51fccbfcc6a58ab3dba9ef2465618552ba289dbf48772054850242ac9fc099383b345f5ec77ed2d535319bf89ed6fc4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha184116f38e4f66d019c364f563737738684302af261166d50d6f141f6324f1abe0cf34e7971cdad532a2e4118b14ae3eb93f01200ebd2abda6ff2f2e86c87f756311adcb772bf29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7902d890dc8b9360e832016624af1d2c01ffac8ec116ab2d067f0cfc0b90379aaa57ff4c71f67274f78e40e6b5e40082ed81414bbf0d81d55540c7719ff40f59a352701bb3797e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h749053c9845d52d9dd3cf3a8cfc9ccc6227ddf3c38406f1f6a46a116ceba47e1ab4aba866d5b22dd3fcea69c0b643c010a0b1eef3b06adb2d623f294fa020026468932888bc8c828;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h581bb85a51024a41a78d2dacc71ff4642bb613a98a82a2409d2450829aaa0d3cbf8b2bbfa6366f523ebff14fdf48fea33cfbf2c84371779149f6891ce55ff8ed90694849df3a1c8c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dde587810561ffe202749c517adb228f7db2454c6d991cb75bad52454395f9cc45a52f4e4b2d9d9071e2c634ff7e1fe136b76cb4c0880ac167c42de68ba4c2ead5895ef44235634;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76b7dc1528a92dce5893fb0c3422c445a5887f3d49e2ae02dfc3f47212ac2446d04c1acbb6ee159d5c3a1bbd62ab5e14dd91afc7ef119b70f7d4f14f5cbde90dd318882b161d6842;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33304695031313376bd42f4e220b886f502b90dc6d17e42adfb8bf7975d894fb7e1e7efcd5a49efa3b1d8f78141de253313b522069cd0eade6b5b78fca861aacdef9257b3b395190;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9da5fadf95fbd1858fce465c90fee44abe562c2794adf70eff464bd297f4c42062c30e521472a3d55554fdb52f1549a65b5511c3d866a84532fead4e5426d4dc3df9ba8833472e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb79f74364158c3b038eb4c82525af2e88772982e59b05bcddaba66102247b208e9f9b4de1aff166eba280ce76d8c6251d7aa284336d343d39584d31ce3bfbd0616362c5a3b374e84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6f000d3431c71b55b6fd09d619920ed54e9f32798a05fd42b2bdb734434c62e6bc873e7b35703f43e4765caa85c8aa1ac6c55b7663b47a0999a63f0350a4f8038c4dd4d9d9e5ba9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55024197dd04f9a40c9fecc27cfe9aef64c9937c62b49ded21a471431041977cee5aee5bfeee8d2a6f884c09cfdc6b47654ec517df46b120fcf580019a44b785471515f790eb96a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fbd57a76455d3147563c4f82ca3f513604750fb502ebd46d3373ebe5ba033d359567754d0ae354f109f78f6dfe4be21b02b2155359e0c1cbb4e0d0356a803eb2305afe83a3c2ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf68833a039cd1e9bbe6dac0e0f116afef7a5e4c52a6583f273e32adca61768f08aa0cf98bf9c820031774b77370e84d5ef3bfd792db24cb38f9c7987f50a5b54ea260f409e9a5b71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46592c8930e5bdda1667216089e0708eedfa6b20cb7e586c2fbc7cdeea3a895e7b7389f4644ca8fe76a7a26a91a2044196cec9e8494c53073deaa486e1a6545edc7e83e27c8eed03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h359a7c4681d0529599c5777881f10496f848aa3f67c9200b2f8a318954e8a5c16f4a8906afd21da30b1acf07b636b13b67151e52d45678de0aa06cc07eaa95edd5788e7e689528d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c303d253792915a9220eef9c84591bb5bac248bdbf171cd577d052482d25e1c83b7c7fe9c8b7445948495537b7fbd7c5708e9930ec2666e1679dbe7eefd2cfb7d88837d328551ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h279d495392dc072b3dd0d24c15506f1ecb764d3b04e449b3e8651b0a8553e97829a980a219159097bc118cf9318f0970d055a735b066a08dd0b15e7da86ecbcc524eba418583c762;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62d7484e6538182ba52c7e236754e62ea55fac5264628c166b46baa8217c1adb735c7c4ca052d5364c6a691649e96c7264ce9a82f98bbeec3802463765cc7bbc7b83caee5d5194e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h203a81bccc5dd71d1bd823b1c918b26b69991f5c21dce4f2b35e49d11bbdfda39cd30b01f1073d05f2f5f8478fa4a1541eaf0c64462078ac28ca939767e464791bfb23b25cde42d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4b3f5cac49c79dd3ba6f6778cd69989cef6ce09577f1b009ef6d77ab10ccd1df7d7d351b6198caa75aa4461438cf4658fb5f17ea49eb413d61844054a7eeb6225e24053b50c32ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9accc7b451af1e4454b6539c8b93fd8ade2212a1508f8a21d17cfd6e30af299cd08913c6b7ba2dfac21f60c7c013e093d7ac2207eb977033f098978adab7c5fa16c7fb2759ee6b2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddf0c5136e9060eec00a480ab40746805f6bb13091c833408c21107ffef50846b9bd013475feebd66efb3022494ed2eece004a565a6d503a281d01c73e7495f060d47248c4b7ce51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc35c9bb84bb326fd85fbdf0ddfc74324bdba03060c9ff6b7ee0dbdddbf9ff33cc856f2b00d76151588fd1864863a7eccc2b099df90306512509e1832d4a738196245133431b3336;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe9460a624f6ddeb69507ce5d313ffb5c8dee319c920fdc99471d5725c01f9d0af78be660b63754844fdf84d282b2fb954d051106ce0d567b738f8d4410f06c882ba5901ab34efad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b21c3242e17ba89ae14250780df4026ca9a02592c2d7a81cbbd90dd83609783d0d64b284b877cfec214588eda662bf6c2c5765f8d95276465b941ad451a14dc5f8a755eb7558599;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74861a4dfbe798a31bbfded75b0e7645e7932bdd6e00a507c7b1a3f8f071cfe1cb1b0a06ab2a13bb914f033ff0c59b62a20e0cf41ba29a372dcf4b13ec2316050123155403f236ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf399c96a5cde100052819bc1757be5255667c6f3b7ca117768737784dfd1dfabadbadc136ae3a1d1929a3e354bb12cfe9d438e06135652f16f004d732c36d010c9c049ff13cf7c4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1be721ef22c63d7dde9900be19adab3862779b1e9a2057efbad8e435e779b1683b4cbc7acef31ef58c2dab1d09698cdb612c0cbfa9370b620a4543b74d199e2c81d173852befa82d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a90715da1cb8b8e6118751d6df01eb6150361bbe9cb0d8cf3d69d5b1bc39518181eba12a1e75e0b4f87c9f7087b021f0e35c2a572cd3ac0c697b74d76fca26ad3183e6da6a31ba6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40a67bc1bcdfdc60f8822b39e1d05cf02ab2fb52f30d97a8f8f3d71fdf8a546b3016eb12a46d1c6f3fe2736a32c0981f2668f54344abb9d96e549010846c0b0b1445bf57e81a7d05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4e1f503cce06a03ec2fb6064fa776a1b7379ac01ef74f304636664fa79cfff612e52407d6ea1d355f131aef16aa2b995800284996c2cb0e897787ee0f588df0852273395da20c16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82d287335ee3d60044814f28fd92c8efb7ac2a2cb105b2012a762fc9b572d3c00e4dc93744431f04bd75c3180b293b3ebdc4e7eb8a06f8a74a93ff6641eb13b1bf417e5eaf503df3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82f6069d67e0a834e1de6dac79df0f75502471d1adb7cf02bef948ce245bccef80b8a00cc06a47d8e7e5f96185bbef5fe1254e3bcf8fd7150c400d0661303c86e625853afb82c28f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0b3d662d260d6be636410ff872ed4f89f0787a93734aa690b1c1cde2689419f341e7662403d36fe618557419680d2254577da2bb202af76bc5bf58ca8844f92cfabbc2eedf3f6f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he488a0df84739b11053a1c848bcf37fa68dd0172244b51d8e67d3ef6abd7888b8d1367cfb8811bf8c0fcf5f6259b6c105199d6810b15aae562d5c39b90e74d2077b799db95ebf191;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc2b8ae43f17d2ced2ed717ebf0f475dce32e2a5dc4805c754cdd8c494a0a48575110e14cfdd3c29f16a9eefa07d9d3ca3656dbfbfcfff138eed6b1fa708c63107b2e1ff4924e5f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda286ca1e4bc0f5affde9bbe65ee1d73e7869690a269ecccd104eb5d653c77ba83d5cca02fff25dc1a9ae43a93ae6d216c2762644a96efd2ecbdb48a560fe979bff48aaeab3c096f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5fed46916a7c04fe61e9d6ad58609cc0e4927e1553f5cddb5056f67f4ddf4dd71ef9407762968cdfebf3be99c6b49fc8b485510f89064a021f68509a6f91a6c820343fb92d4e0aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1976aec1b00096f654678db42c11f9d7ceb6335a874b079a72996fcfab4a76ca1d278f8dc6cfa06c1c368ae25251b94a90f4edec8aae79d2767d8a697a086942962267abff7321f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e6606918cbca7dd48e80d37c09b68a715c72221e7fe1291f5e13f0bea814f12544e036c9b0d6b8bf11a6920ea9a634544a6531120a9fc4b07d87142c83f7837c68e7faa4a5efb51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68d52954597aff8f2526e2302a7df6d23e6472d5710f4962051509bcbb4db8480a84eea0868e07dbeab18bd29f20499066d936656c28e680e0b70e0d2de6b46e59a872bf5f20357a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b4473ce7ef3e7f552d38d6c031350cf6220f1e8b470fa1811748e8d99ea11265de69abf139c2f6734aae069d30e4d049d60fdb7723dd023a32f79a23639a710b7032e3fc304cc83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc37204e81955487df70dc3d950f603006607ecd458adc5765715d6d9c98498e5f97644a988fda9d315670193f12b2effd584cc9921b4bab64c0d5e84dc468af914976d5c0ab9c99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e13cda18141d796f61d94b80349e43a7b7ebead81753105556a197ec8fd64c676f96a89beffe9166496ea0590cd09af754354a221e732a7bfcd822ae49a175ecd72a04d16ca795b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6203a831b9008a96c2c759abcc92de5562dcc346623293811d8486fac9c5439ac2e405620025d8aeb9ac2e5f1c5881971b02412824f173c4412b01b0e76babb3e22a2366bdc9ac9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h523614da8a69512a5b66533c64732c8592d20ac1a558290f735cb659705d9be6e0a130b21b4fb85295950efa571ba58a8099a2f5270626c8b2c2f787bc800d8fcdadd7df708d0e2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c1a173b88b6e2f866e7d1d4177282436496a0a415a7bfb10d850df6b37e17efd3482126e4173c9fc8adf1eeb758dc9c46ce3c30c6e4fbbfb2eb6fe5184acb0d561326d9e7795a61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8676f3db4a5aea2f9467895d0da12dab647fe988cdb555b2a18af3a66459591606a9b4654bdb4a2e82902c691eb18ddf31b12fd273d2de6d53fa6cb5d2cd0c9c5e20fd107bf5892;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15d59273547ecaff7dc7fd9b9b19aa26a75493fdcafb58b89a461d5fd15d51a7102d131a059a9506050b3bf3f9301cfa9dafa5e18bf506304488e3facd1250950d4b949099716300;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he84364dacb67702cb1ce4a373552ee3c8d3f84f971bcdac6fe88b0b1fa036a4ab247290780df1d6f27d49a07cdcf85d09ba70086dfd0b5719784b74334b7823fe1a81687470e2287;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0ebb4d84b58f74da81c1e90ac6f780360f0e5e8f54dd12b82a03f6feeeadd3eeace580519f4145bb50449836d27588f3e57071f8bf86cac2e14257c8dcf1086bf22084cb5a5e60c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc364a49c91c3c4a307c5627747b5c5323a3ec7bc004bb9d9658f1cdf3b8f24115977f477a76965d68386ce59ed93fe2511211a5237011d0979ceab8ba1512c767a9a0a1b8030dc5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31fab2a4fcf2945466df62c09c4e24611630aa0cd87ae6280beee01bc9af34f140240c4f2128c4520b1480ffbc7dfad42756c4f28d948b2f2b846db6c66ff2c976fda1fcf6fc31e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f104cecb594acb2ff608ef9e326c7474e538753e77dc6741e72a1c1d8602473dcdf0fe7f36259dfe8899a792e6df9f8cc0063415836b40deda7fcdc09a073e1f56f5014e078e985;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80826f2907663eb04aac32e261557098bb40205c8ff05fb7977826edfe5a8a11b58e87b85deede0b02692a831f4c62ea5d4059736c007150a4341c55dade665183ee56a527cf7b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c391acdc7d627ad3b295d9a2f778c1f2f8428d83f932fde25841d68f4f84fcfb5308ab443b4b153f79763af2617ce3aacb901aa82a1640b1d6aa274b70aea231abc04dbd6460843;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6f9c29d9f8fa8d19b79bef12b1ca99c71551fa209829101bfbb63c9a3644117fc5026c020e47ef96394c6202b18e10c4384089449dab5fc7a505d4f6f4343180b1247f0fc7f4d3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf11790758730ee127fa9c4a28b42e0ab5c16222e0ebc638d4f9476c6793d934ece00978ecb595f92ec55ae76f954af3d9dab470d24444fd516441542620b5027e37419d3ca001487;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78b6d27de57b4e8cc6a8b0f4ea87f42148b613eac8481c426eb28f53ee34ef8c40b3a3e3a19a7a3b5329e97e81c47a96a2a79fb587be52013aecc90015a9897a3e6428850931e3cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23a1ae6ae95228b630908223f122b458035c7b5fcd17beaf1c1d9509b6a4d678e4d5d2a71e49c0894b51d3f2e96601e552d204fd3bfc2b7e7581b9019a4c594c9b4323ee0972a045;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1351baca1958db5a2b06369b9c4e7af15c408dc91d6dae016fea829f7128c2376434f20c7319b2dbbc82818cb14a106df52e2caf99c132a9495a6765c2a4b300cedaf967f527429b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0a038f84faff056995ff9a3c8165c3e497bc525cd86a276956b185c7b154132330f9cda9a3ecbe21d7cc898eb6e8f3066bfbb59630e3ee3f9ebecbb97b78f022b05af18e24a4ec5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4246e0c352887324f162f11d145b4d4e05e59f832940b04982f2edbf4b19cd4b7b5a91eea63d06088be9d3898f34d3a56150b72f7064c7e387ed92abb8ef84023556723927f5f2f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45fd53e3e54af63d664635485097bff85cd7046ec55f02c37d6963f8013d16ee81556c87f6e4c50c73edd27dad4d302f4571c7768b6663b5639e57474d5e7530ff87ceb0c95639a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5c892adc2fac27a35b05b6437053dbf88b2a8acbb6b9ec75ca2a98d44cbf5363c23cd1f2debbf029e757bc4a8e8a60d63dd8383faa356dc01e8bb16b382e0f19fa866661daf094c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf83e1f383368958709f36a70d0010c83749add7b9a4328f2ecd27e2ee98901973dedf4989844228db00302454487a4cf0a125720e0518e735a8305ea8979cba6dd4752ce7d247614;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h997d0d4ec939572fdf5ea27911b83c0faa6162fe0ee3c450748f6efa064de7c530f7f2fe2f81f69b70284cd8f09445c9c3ad4def09810395e6ad543b9736596712b1ffe43624816b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d415ddfd9de1a1beb80b9fe1f4b77a7f4e7356edac7c32c9d8fe01a398d3f6fdfea788065c0d78f688862087469ce18357839d5122150ca96403da850f1f75b5fddc284766579e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h532d36429c4024de241655d97fdef2ab292647caaf141ffac2e5be25db573316c4f5b0698e975980da9250a3308091a505eca84b059b764a427be1165c06c0ea73f1c79f67af8f9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h691fb78a2216583758b52006f2d78be31a04f4a30958749fe3ab602cf4e61c40bbad567fc564d3ca9ddf641c73028432f17aa1892af894b473e9000e02573fd2829d196079ca6f61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f91d35d4fbf22bb458ff7abf21d9a02c73967f6b7600c02bf605121025ed77c62ee7bc4626b87cd40b4305b4a5d8a1224b8022b734b102e6b9fd17416256462ca6bd00061dfb14a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77aa0b3d4880418461eb62ef2cb38891994ad2a726424cf1b6759567e98be5ddeafd2f13b2c9a16b0174bcdc11354a59015d3f56cff7200d48e3a9ca3bb28b316a0fde460be7de6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bfee2dd44ea0f2e67af7d8f45e01f87504ebc3a60c7288ce33f3e4d3db6c06f8ff4fd721ad6936ea104e43671ca11fd653bf4177841b96edd33387914d981e5a27b9d6737430e1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61f3f4c7b5ac4351386a83ab97c160802cc1e3a59bef5255cac6359492760874b0883ccf992ac8c20f7c95369e10fa793d4af2c1bd713d11dc0bdc21e80d1cfb3ff8884e6a3f741c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b0c7fcf4f5ab6af20a676fe5e63c768a7aa3863819b3884926e47b4eb6b2df699501873bbb53abb068e411990afb5056ca57f2684649443996ebb398f9c4ea3994c9662e4de83ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec1caccccd0fda7948f4258aee31bedfaa5acb441313b57d7b90ce18d6a38f5894e59d7ae2d9157e3c6f37e109b1f8739a4e2744b5174b887bbb55097d3326796342cc370a6a9e04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha46327b9834b0775c475299c343b569c7ef1507748aaddd20c36f4144e146a733e2495b549cf08b8f742fd076ffade96fe861c38de4d9a504a33451a0f21e192f05c7d090886f3eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86933e570efad82aa90f2f250bd5db1d42035240e872aa5fb3268276e0cd3d0f96ad31d092e2b6ceb646f09cb1455dae6f59a2690b2bc74c4b91eee20e90845cfb4ec32abce7a6bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd6e7a7aafec9c60b91b0bb8fca3bfd96aad0a9c5e5d2adc0369633c166a9a1ce95c4a0d0e87781da9f09f50437accbc649a09f344a545d9ea6b374aab70029b3ba9af23993c8ab6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac7e8a4d507a60837a9ea8a3fdd56bb9410a904f7f607811ea537d8dfec8d40a444d4e757fbfc2e5a80c7dd34167cccef8e6e2bc0ef08ff48e055327ce045d8564dc40b8062264db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h283508af201dab1ef5b2f097a079e635b962db267753fb22974836d7e7f54e2b590a59af62a1e2ac42ec0d58604ada9b406417f9ca36d7bed528c354af5548d4905eade8ab9d29b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0cb85db65058c4b1a9fd3da0880b1324ab533b295093f6c5f127536a33cca71e651b04697e000255178f599ddce3b8c18408d6ba357372ce19c6440e9c59f12f7814706a13ca4f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he38461ffda8848d34e10666f2dd4996546068e7e005ec704f1359707409c943ab05859d38b58b216affb25cd6bcfde649028ec37ccf93ce33dab6371a6e6240c57b497ae00a3ccfd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd62e000e4f53f8468a57095d9180c18e7237c830360981a6418a46cf42cfdab0f04f6e958b6b7c88e6177db5357e176582d000b5cd5bfb11dd5c97f821d909307f4f57dd273bae9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c7a57e22c82e08038baa5bcab6cf3fb95186985b2b21e9a84df1b3977bc4b7a76684ba9da506a05d5cbeccd823f3d6d274aa878e7e0d9772c0214fc4df505b190ea5582ae4c1a62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd13ac104cb5f5ded99f9c12e5000d263c990072d56489e3c0d011efa0e57b74d719ba53f43a8a9a2198f1f32a4fe7c2e4b20dddf26492c0f71f7b0f8ab3b4e3602a59176cbba09ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba5d40bdb1e5a6cf0aff539b2dae890e82e8ff665e20937dfc2ff2dfed6d99a59ca3a3b377367b3b128e5df060fc5bf84fa99122dbeb64798f679d90e192bf4c1276d01be1e1d599;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h818339f63e1c3a5a9e76fdd34c781251572afc9f8b82f4dcbf4971595bd67452dc9ac6724971313cfcab4de4e0ceafdf25e29cec6d550a22debb996936f36240bbc15c507ddbd7de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0271616a53efc4b244de2e8cfcbccade1dd237797a1e850d96b9972d2ef1f817e437d0934b21b4f38c298a92e04ffb5b16a8594525fb8a23acdb728cd99197f36fa3e46d7d8ade3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ce68fd512c578ad11b8d2b0c32575f6e3eb8e6b6c0d9b454d28f70ebef3a0865aff2f1108a9ec1b13a37984d337091c2566226ff1867621001ec67aa0ca01dfc5b41613ab59752f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c28bb710be077d96104650c741e65d7018094428dbc308657ea18c542ebe8e63fad567781c5a6899e074982b20abc5bca49f83072cba04f31729865e98431ea0662c1e2274eaec5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he63e500a81cd03b75dd41e58dc324fc8a4c7b8384e0f386df92d9fd5b7a93b61ceb8398d7f0ef7a2382eae4f6402c51411e589d8af0798d942fdbb833694287a5bfb2d8f8b5d45bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1bc5f0430f1b62bad821738bafcf20cafc1766035c4388dfd920d3eecd64065f4925e9aa17cfe37914c6a678461a05ec16027f621fd3e1aad635ef9547b2d92191d6ad03a33e610;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d09a446ab091cd4ebb0f876347217e424367cbd4764b0aebf39f3e9d0b6f6145bf2ce5e6eae2f417ed7c7469441466e516fd9afe4f930e83a9f905f0e20ba7ca479784f94e26695;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha38efca3aecc038e13fcacf2d9653aeffa505d61266ef0ed783c8eb4f411531b2302f4f54da0de684d9f15a8e2c8b7c91495ac546788e0ed5795dcaca9cd6685b7d9a61f9858444a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11c17f08be502a0069ef0fe05c9ae42fdb2689a41b955edac6baa014b439d103c23bf5af73e20b37a0bbb65a183164848aad7ab212b19e45bd604747f0b158a09b909fef8c6131b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9e0281bc29056d9d92599c661292c863515c6c5c8456c32a23d6854638a024cc76aec3e9ae9737ac110ebb50aa03b75145473d82bc101771019646089e0830f00ea68e9bb9d3c1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7bb9127d71d1727bec84a2b84d3c2445c2bc3aa5815eeaf6e457e254d6057bdc4798312f36aa83e68e328d78167dbeca4b8eb3fae1fd53d1949ba1200d9a5fe1f0006ae5dd3902f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0bbf8cc8abdc6e86391350804e0e2acef12938160a45c2904720a44e16054f93bfbc57270e7ee6bad8645969a77a57fb11b85bbd7e12f93fcf9889568696712e0e0b5a8d23eb11;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf60aa78eea1c86433a31a4338bd1ead86d172b98ea4fb43e113bd7d8f3c66e6ea9f157e8aa120b389e58f121fd6809c50e32c81e6e060f9806a0f0964f6cc3eb9cdf9c88a0e77baf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ba0c167fd7ca0dc29268cc407e3727838596ae23b541295db1decb752b870526147e4d71fd6fcacca3782840b3d552165b01c7c00356796157fe67995af20f8804c54e4012e8fac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecabdf0e2f65b37f9443ba821ce76a1f76f968ead901f3c1561551a3a99548ab5c0027d7bfe0389371c4a650adca31fc485483c747475f0d9d9884756386c67c51e8def90eac495b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7c08800d0c6355a5ed946c3b3a68affa36617276184354ff4f7a00a17692e24fc4bafbfa101027a51534af569bba8598ec4b41c6de23d022f37330137fe1d025938553355e2445d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cbd0692df776781ef02ae0138ccdebb9eeda1b8963bc58cad3ddc5119a01995676ecef5e8bc6d17cefef9ebd3a1360494a27cb0fc4aaf678cbbb2ec9c2e30770911531dc9ed74bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac44409b130e1c76c5da97085468f686fe16ee2a097eca828f806cbedb6c8b4c49773d44b6f91f1d1a1d9724718b22379a3389d47f902494419caaf42cbbfa3272fb78b59972fb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96da0be29d35474a992d41c0e6ae0e4f88815f3828e5c7738942dfc1667c220891475884fbe3ac702fbbbae45a484905296bd9bf275d2e6a4c8323c78b26166d0544aaa4979fe55b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h345b5434b49ae6440f49d0786df1e5960189e03e9b7f82f15d235cd030203536395071161fd8f44e53091f94df993e55153b5afe54ef84123de4596f045ea45ae584deb3d6173b4b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3037808c687002b76a84d7aa5c97bc2d6a9fad40d496d9aa7020b5186361296518a3a69665ef131a18125e6f089b94d63a71cc0bdbcda91db0880d31132f2bbc07e19bcd2d6a262a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95acc7944da6d05b4750c1f1b6ab6784663831e3f426efe5a4144f53a5ad2b00d16597cd451c3c94c4644129c538e9b6cd1b806aa081ebdf5dc055d26e0ef9a0a284bb787b021c53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ddde99064df48933ec850a0515d6afd0939d657990fbf4e4cc577b3faa24ccf1e3c4da5735f7f1d6335df7af5ee42ae0936f2f250d6c109bfdfaee7f19409f828b70dc42c80a827;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ea3725bf93bb4185a8a1b30f16271a860c26dd9980419f8538a031eca8d53d46b036890c221a187b91173fa28d286706995b087ed7b121370b68035b570cd68b4d79c752bf03ebe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h288fb987c2a12e9fdf3172afa57d5a0034358d66156966f05ac84f7aec2e5efec9ed48e708da4738b335a3b44a59c97c656666775e1b4e2d421161816cb050c48586bd79b4a96e34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9817c5c5de9b12cc99660a3f59e8cd275f0428bff2871d86061a03c8e461d1330105b46e043d0c23abbb5713141b209401bac9ac9914cd97fd7257460a5be9437c151caa9f1a21dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb333ad749e07d152d59926383ce3dfe53f579a1396631ce0dc249c4f4834af683fa3f3ed029566785f9e5ee50bffeaff6322d9b68208fb284a1ae4dc891caef156c4c47ee17695b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9902856a6a49a71b511b1158ffa091fccbdee7eca5bc5eb00b83d0c7dbc5e7833ac1e23c9064144568a0f0ab50dda00e004a43b2e80b3663f5a4fe3b9af5214d66b00a8bd73ce2fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9e46516527393fae9a772b52fe8f227f849b9f693cdffeb1d1ddc4c359cb025f4abc0371d9c536d387849a537db1076a5195c1999e40a63c5eac94beebfbd8165406a4586d9d152;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4da51f2129e7965d6428d23bfeff86106125eea1f3e94c61a1c6d25dcd714d5478db0fc6cafd1f8edc29c800fb2044bab10bf5bf9ab4cbb50884cbb8d81cc6834f7f3f7652df2005;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd06b070ddb01d291be36e1519f583884aacdc9baf36f15b4168472b6da26217afc41c9e487b243aff219658173b56220580bd05135be193062f8b51a8ad873fbb05ab275da8f657b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34ca7dfef1b5c5c4f82106026d2b6ea4d7101625ebe1ea580d2f3a3d13f9208bbd180fee6e5624a42b25ff630557abf9b0f307fc31ccbda6c93e53fec209ada825bfc7afc3f99afc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27d363157df231bbac73a7e2f87ebf5929add5ea3d0269ca733cc5443dae0a38e80fac22ab7135df1dc67a96c9d956d8e4006c3888eabf18ee3187621d9ff98f65681bd6efcafb6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc271226e15d0dfde655338d77f413969a18b99722da9deeefcbe6269284d53876dad5b91e3563087cc8f30d41f43a54d2f2494717f146149af0c613a9841b428a6c692de47444944;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h836364b1570aa7f97bcee1736d47f40848f1b8da517fe622b3c15a2e9cb89dcfcbffcec421d4bb4b635cf0273c23f0d5503346e8e5f188b84a7feb72eecad01a29e6cb3f335d4340;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2374db81bcc941b0598f756b3aefe5d5dc64ee67de1764e73dd7f1cfc814652f827b858203ac4d8d1c45eca971cafcbdf33a2899fc0c9f89fa055807e12f400ef8e2586ab5b19ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2207fa8aa0c185293018df5d9675999cf594f81536b31f134510650533b022755ed8badaa9c3913083dbb28617a685c583356f5a2db3d235354712410d054028bfc07b8e11a4899;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f10957a5a39bdf6f51321e73df659658383075fdc131aca09a1e92c1f524468e66f9bb9efcf1c5dcb02bae4318f8b5c3c23777d16351f2bc68a9a00158452b0f2a3ad37725134d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9508dade7a8279444e3800ed37ba845c236ab6d1287cdfff72a2cd8413c5f42722bc5010c199cfc2f51adeb0c015a82df5052be699e702f2c324c2b4275d786a0d5f0ad5709a1084;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3114aaaec65aaaeddbbbe0ae2979ce4c31c6110015c61a2ec174dca130ee93399943ed321530bd9903ef2d80c54862591e7cbed6615768fb16a2005f09eefa54746d90dcd763d0f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7a97fcdc333e920445d3588b9615210612e3cea6a359dcbe546c88e71c83c9f8baa9bb1b530cc4f722e477bfef1382bb22aed7e2a94090bb5295692786a648599106b1bfea98998;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbd8f7700e54b6b72f0a6bae200ff87326e7be94ffc9c4be92ae42a5c32e9f4f167c51518bf37df80fe34683006e051a925ae39d8618028deb6c6f2fba591cc2e17aa5cd58e63900;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebf415f4b3b532b56f1082eea1892e80d074c066722d5c93865929eda2095d403f0ebb1c4dee6c51282cf2954888cdf055b638c57a367ffc7ca17112838a1e29df0394b2d20b4c38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a059e385bdff1b4f5c79dd1b0f1d47ae8705a68d8113779e8fbd7f4aef19e8c1ccb4626db20561f314ba4f264485abe14617a5b5ed30153a46c950394332e6a1f84e4eac40b2f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f0bcb717b157f4d9e11f6b9bc9e3a42f30f25ef6986e43219d5a5b3f7e97cba07ba65a1f20a51dbc80b4df82c601803ff9239a2df8031749ccb298314f0edaef558b9ba058702ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd3b2d9db03bf5287285c4f7f52d2c66869ac15ac26c77e6a48e4e5f3c00d4d284643c36692a82c2531ea76d319e3332b6692ca1dcb4e01c0909b63696f579ce9a917ba97b7505fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha403139bab49154da43d3d1cc8ea5a7be04d1a68b7981eedf5a9c3e561e4974ced880ab4b519615dae1b8b1c16b63e1f28c08441b177f9dd27bfd09a44f797e61ae4a71da1af0c60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha219f3e383853607b0ca4c911d567c687b9bdafa1a66e6d63e06fb3eda181dab4f29f66e011ef4c6ab9109e50e9efa537e5f548c3a61a9dda92694822b262fb3b1aa2564c79a8cac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf27f1e45e7918d1af5a85c982551b27ee4d34177f2b8a6cfae0376cedba252b7fa92398daf6423295294e12f3c56b15b5ab1fa52294839cb9730831cb0e75e684de2f55de774c0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4359289bca9dc713f430f5e19386e319e4846a1a9a33c0c5f2a9db311230acfd8450319b187a40315d554dc6ddbd2dc2f219ad6531eb6ede63315c691ff5b3e7c782819114fc029f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc85982c114bf7a4ebe6628459125832844ba0f099dded9b276a946971afef527a9f2f9dec4b89f929b657a9e848da7a0bd54285015f17a612ef60df65dea1b3d26a80da52289ce81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbd8f680b8961efcd6c4b6321265f3fd45699e8d1ec6f04af5510a03e861449061fd1f1bf3f0715fc5f35c29c321be7b2a008728e719c64821045a495f7db1b68dc05b94d3103a97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd033c2b4a9bccfadee851e9df5fce2d1b42836cad4c5e3852e118baed3fb226f36fa3d293c1f6d104364c7f69df321bb7f9687c641d648646f29e9452bf8c5fdeb973daad66173f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88ce7ca15724baa7744a86f802df4806f705e0f741fbdcfee9e078099aaae96861e01a852f6e09a4d092539d45fa86067703f3bbfdde3846d7348e5bbc867ad9741e2b8e7d0ee8fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a29970770d1b29902d098346e8996015beffa2fe5f6c36e6cbb1ecb5cf67fc0c21c64aea05954920b92326ff7f86eb863d623479c5cbc715d4f577a291a45481d79f2b44aea8762;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5462730a18fecf30a0fad2c772c4f83614954f086a80a3693b18dbce7adf7708fad0f42c54f22fbedc879171135fd56003a35a388da3e43fccbebb924d776aed4acfa126d7ff830d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4630cdd68069cf005f3a52eaff84b5c249e6a3adea065950c21ebe5fd4574c7e11be781e0d3c448612e2a8a5185e5f1063d7794ddca30a8a15bcb08e289a81fbaf4f433a715c7145;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2da2e40dd938029ed16de48210a580dbf6abdec03062cfc3bbfbc62f52260932a0cc758194285ca3fadd2f9530d68b4abd935c25115500053bcfa4e171046cc4c91421b9357ea55;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5403767173005502939a8056fe1b0c16ce03d3c019540bcc1f1c0171abd66fb79092a26253cfbf12db3ac896d4ea3784c909799b8a99c7f47823ca79526ca1c68cf85c919c42cdaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he48b99e003e58c2a444977351e3292e5099777af2a640f3683789860dd2fe316adc96f4a39c3100f404dc6a0052f937d73c081cd9accd545c18ebcce9e87abcd15fe23017f818934;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heab3de86aad5ac048c356e7c6e0eda8a3927fb7792d8f6093aae468b59c06e65dc1feb9c1085434ea3de5238df6854d2174066381165782f115c5efc4fb5f2eaf6f0d206cc46782c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65568fb8bac4ebf70d4e61ee3a3116fc8c529ece6619ccf33146a3117eb2f4645805432e59491bd358b2e1976b43ce99ef7667393cf51893df07168786547e69755c71da72538a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32751f8a76fd315ca9ce8fdd0184e2b237e7d779baa22060d69e758fe4aeebefa86e3ad22932138119b55a68f95c80d2c34e4e9c026adf253b5adffd185ec3ae01a4956b02dcecf9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he111da9c0c774c78d35c58d3bb952009cca834cce299e29bfa2f2dbedd10ef51148386eb4631105411d9a738570c417dc4e11e68cc2170694736fc0a769ca971979ee5d045bbcea1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h933b0e81af21821c150f085fde8a069f3449c27e5274bb9e5dff810f55263fd83779bd340d405a8e5505f4a99ccd2e7c7c61206eae6ac3b6498589490d14cbdfc041ee9bd7e66f35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0d13a676053fd9c60f990a81653188c7860dadbd89ff7a975a4525aa4069346ee00dadc9a85042eedee120c21acbd1fd1a8df7383d82d0a316bd5e4afecf4f0c4fa56be8cae9953;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1eb6d0b5d1cca004d2eb977876a5d44517a08d544a959132cdb5c8b26df6a13d358c4f0260f6854d55a9d0285ff03fe6923de1d211395bde55b5c972211977c64d9f40f27aad215;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca715f51fe2e80f810687141e891569234150c9e2fbb199e506efc6c5ccb2a1bb1571f0620130ddb6c1572e5015aaa33342dd1a67ad7f988998bf11d264684c67ef987d6fcffbba3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7705cd84c4fccea70bded2254287dd80ba3c6fe52dfc2a7231d7dfe2f6567e97242570e6bccb072bc5dccdb1898428b1f6d3323da5dbbb1d1707ccfd197bc3c408179804684d7c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca229c7ac7bbe73265129607d7b56c3cb59ffe9bb436c5b030666ee87fde96fb93e0ae98e418e7173018fe6480c2afab01801b4e2b7f956f92d4ea1f04852061933dff03e2d53eeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4b94031f29c4e6502b0b00d25e3b8d2ccfcdc8fd11b0cd7b1dcb591da988d415a0ec9465357254d8056bef4b0adced0da175cb4246d6b704f078c996c2848216cb68f20a1041a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h930a826050799612197721f759b45311bee1d55c7161be5ca88526d291d5cf99ad5a5db7f919132f4b30b5b39250cc850c894e89e5f316bbc5618b6c737cc643d74acddd5049cd0e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5149e7d848c146310c517f42ff4a72aa5dd4b641a691c741955cd6a161e9dbda9e1f2711191c1bf0ad771a70d3216a5e1e3e47597c0433f8a048185e30886338fb2acd60db674cfc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16ed40c296b65e09fa4ac0422b9917d5f39c01f76c1334ac79d0a1234af5ff5a1914be823a7cdf40cd153e65432933c4de477734ab99ce31d0185a03bbc2337fd3ea86b713fca1fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he393a70c63dea1c9425807c29cb23497fa261c8deac354e996bae00bdbb683058dc78753b3b2328a8ec1a2c75b49c8968eaf13ab92f04dc75e19c112c10c5fda6bd1a77ab4dd84db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadc81dc4f898889273cf8cf6556cbb6ad845dc8916ab4c432a6dc30d5135756fd4bbf328fbe52db001805e657e4ea9d08e01c9e9a027160608aa8bea531236fa7e3b19cec4e13f66;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ee720546d469ecc1e372b133cad5db868d26bb76e33c517922c0ce1228f37fb542e4779d2030f489c4ae2a3458f8f2a55eeac89b54348cbab3b79771d81b4d790638998703ea98e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha42ecc11f865d2b3b6822da7e17b465951a7c2b3f3e4eff4a7b8ff8613b22413b0502b575e5d5da807e8016d12de6ce5f8faa4a200ce09dc56eeb9e59bb78f4da8700ffb9089115;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbdad24f9233e11f244e3136f307c2e7d2ac3aa9a44441c9b8fea474895bd282bb960f5b6c3f5123fd262fae7e4e56a78d25ba8bc0bb0ec6182ebfa41b1e338d6233805d9806be3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44daf015fd6307060e418706573e68910cda352958152505fd3d18ecfddef93863fa4a0ce2ea1025b140b491d7bccf64005343377cdb6eb1386dc4ddf4606775770d1615831db4bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7bb49471b1d58f12b0cc963517e89171051663826f9000f339b2769cecf17dde4ae079c4fa094c67490f9de32b45cf5269ed813c350db8279a86baff75e9ceab6f4e48c8e1d4935;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb796f25c12fa0def034747389d8537053fa6bccb937003df728f5a728f0fce64ec497ba6fa6174127248bb791267d05c5dbc78a20175a73b6b3a3c5845f991331acfdf87b37640a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h259c08c7ff6645703430a29c8c054f3071c119eb68ab561ae8533a2605bd4f4d53a6d90b2f37ea2de1b10a0c432b9516c279749a5aa3c0a4a4a0eabe640b38220f62c844053b4402;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dca871e1e724463c58f111f5bbb383721e3b7c66c23f2bddfe8780cc725a02dda62c9dc1b6bd69d49e792f0fcd018ae35292c15b139c43a7c20f4ac1ab374cc86b121a72c666cde;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ccfd106d32228b7d3474755211ca46f988e5a52b579b2c02a75308591e13d8eeeb3d4b1e34e1d9a46284ea5a28290df0ae97e2d5a8a08002d5a47e9d088fa4c6690c8349ef877b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58223df1efe633992a03fceff067ba9b767ffd8850f35ae78f10e1d1262e850dfb80b9a19bfef6ce895138044f2d49c9bec956639baeb5cadb8f8a57fcf7e76d1521365780b876b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1e2792e45d771c60c003cd475bfc0e3cb147f955000d48a72d512f5db400c4262dd2fffa3825f011c72443d1223d83f4d703e5d0c68af6dc0a29b70746b12593bc77721e8435b35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heea59b53dd5a7e43ab15a415a20bdfd0545f55cbba8a1661ecac1567d39b834034bd16b401e72c17622847d984ed92bee9cefbf807cfc12cff7bc4f235188fc19d2b4cb14eb025e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb0bbd686524ecc4cfac024d3fea6c2a065864e1f70b440a4f46dcde1355b5f28fb62c682e0c26c693cbe1ae3710d96a63c515e4d17910b026d2b42ae805fcbcb84e6e980e4e11f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf0e49685b78b7f6e34fa8032ddbfb7d16a269f3e9fd354d69df04f27d0407bfda984d0e833c2382f6f03dc7d8883f1c0eb7be0f23a6c098a7487c99f25cfe12f5d4e602acd03895;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h460d9a7ec22c5c4d65b8ce577af669be32935909d8b7f03d156b839a40ff10a01a1d45ead93fb64b72802544e1298657693c3fe164a7915916e4ce6e3b52d13fa16a3719878dc3c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30e845a73a793d57ebb5957a48f518ed4bfeffe033655c61191062be203e85d306814b466c5af2b6963eda9388c7ca9a4d5eae9f4d524b8163844236c0bbf097b5a9bc1eb2ddb6f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0d8c47c4b2dd7484a229226859647d87f6a5511325e795f1f840cea36a0b9bcf6889940ede15fb25f9d62594e3b360547f4bc09634284e2731f5d281de49ef22caaffe6a7c3a80d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49c3b89f20abae787a614361063ecca28317e2d5b2c72512590f9284acc9dc9b95cfa87cdcc2564abcac6355803cbc5a3fc356e6ad3a22996caf556a7f2c0d2d5609f28b4f60c9df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c834ae8448b96d1e3740dffe1fd8c28bc89324f9329dbf67f6a9ba87a2539d799db5e492eaa2a7d8f19570cfba848272d399b04693cc1cfe9ac0a2f129033f7bd1016931b5aef54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76715acaf94c103727ebce86f86dac0273849e723d161e7ad3474664d1618404e4dc0e9f39a9f23886c68f578d64aa835ac0a6aad27d3b47a1992b62c3574461a5114af19adcc061;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6c1f29ae819a9a4e2b447cb12e3479549e1b8f01c7e36a6012a6e783ebcff112010b19fccf677bbd409ae3c98ef9901e6da4dd48ce4b8a1e584e11850347b8ca120ccf4899aa1f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6bb6d47898afb2ef68323a5660f53e88098c67996bd0783e4597dafe160b890366900991f9aeb4cde3312eca4b34cd1c860bf76811e13d2dfc07c756648babc5a7f41b5068bcc07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e3398fe79cf39705e9f3f18b76343f4c1ea479f87976f86a618b0d8d16a9a18d317da78dc26add59240d005708959a13d258dcc7cc962a3230ac127847628e1e519ec076693de9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3439eaede1180ca3e0b700216c6b3621495ecd3a013322a2741490808ff04f85bebcddfbacc52c0ff83133a977d52d29b0f596a84d935621e9ebb416ee4745c9d44bb2abbeabe6e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc45c3e82a4bdb6b4f7f09ce8a6defeca329ab9c25662c8542286ecddcc81333d692e3e28f3f884c58af234c8046989c111b23e6ea4651a3886839876061f91265cad2d0729ce46ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h275435214239a21421fa16686da635280511edf9fb583851c0eac8d7ab791bd12f4702bc506c21cdcac455fd548a666e0a5f4d7809bef5cc1d80dd06987b236f21eeb22d73bb13be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8889bbc9fddcd91346926011c871ba1795aed70d65fd43fe492db41ee789477f23a2da9704932e5457baf73c33c13e16e8f2363294bb62ff6fb576b9a2fdf9fd5c65415e3d2945;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h674c924282b4220597a82c2156e81c1a1460756a3703b97f7dce1ea27fe4555148ae0ca9cc3cd2a27ea70b67bcb2ace0f55ca4f4885d397bf36faa65aca09f5637345016fb894f22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73d9277ba0c099cab855e02f775f7687e10a1a6d3b4d8370157eb174b3ce6e637d58f7ac0c2f95460557cdec352df135bbe96b3ecb256474e33d1314343f339dc98ccc3f8a2f9b87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he24987b4a3e15a839ad909279d45c865755577c4745c0a725e3d76ddecf0e15ea9c61fc9c4a15faf1960db26598f5f1d95e2121bb62a956d9d5916615a767d4e7f6d71c9faea460f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a8d4701efde30d0f0cdf5970f0dfc4f068d4123bc6b9ccb62edad38e8324aa9441821b721a9e65ec660882454cf5c39cc51783f54d941fb6e4975f2ce09657843bce3593abc9f99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19f2094774e4f0e5641ff86c01963ed8d279879923624fb07d55304bfa3979e906c45a41bfe59cec3ea3b5219f57f2e0e50e5eb51332c3e114c35c12bc66a69923d7b6d7ce990c1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc9d87baddf34a79a04e3e32d4bcbea45f926ef46bcd73ca63ebc1979d7df1f64bd3aec7d3590b19b25f6f3563b7b8fe782e331fa1c3e6a36fcac461ca72de08421a23f14105ed0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90f7c0c888c000da5a0548d392472542bbaf95b65f46a194986906c5a0a33eeebc650e43099f62790224e831486b07779118d9acd6b28cd629518d29f2487cda90d36f6c56665388;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f2341b5617519a2ada38fb861fa7f8147a044e8f3bcbe914c8eaa0470f8e099074e4817ee91960adf2e221964c8b428cb7648ab52ed7d0d7bb36cbb6abdc426042d75ef40472289;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bcd313b6abe04a457e545c8f1b10ed5c8a3f721817eb36c264dfb973b47334db46253862ccbb8255085fb134296519a96eaad9ad748d608e5ad8b8c22bf49642c34ff362b516cc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae7dd32dc9911f1371f8199d8d1dd4c0460463c2371bcad1b5043523bf5d71a0a8af5c361e01e25ba4a1c7643e2fc03a6d428a823a5b1598582a4d82bd91b6109af8859fd57a421c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h125280134488e47109a4bfd533fea07c665073017eeef812c20dec0a78e17657190e51d0e9bdd94114c4252b271487a3b4bdea06f1f2c422b3ee54f330ac27e44ece1b83be8c324;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0d4887f4f50559e212ee2bdd6bd4afdb92f11c35e54724f71b400c551801b361dc470be381689c06efc3a438698589a7f685e6a81569d31f7a43b31004c0d381514002e65ccdf8b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7d3385a1c5b30374ced540ccf0d28bb75dca685a82a4260bb90ced70c1f2bc758b9553b9ed8e5432b80f6f6f7400bc2ef858635a33a343198fc6f53cc7a7483c7a55a98a25e0895;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90d60670e68b7265eecceabbe5b99faf355f28452bda0decdc1e0caeaf18b2de236df7306002a55ce64090065caff2437c1a03b64abde486b3932429b37255b8dc4efebaae577710;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c78ba44422b1b450eb57d5d551d4b7caa003c1381827efac30c20ecb542de9329cbba85cc8a816b7963e62c271533a14828f05010b53ceca08b3baccac37e37d8c0f27fae2e554c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12fc960222065f57eee20b6669c0a66de43b7e547008d761825c1fa4b44a03b07521ab6e1d2d051e859cb01a2c2d8affe2e04e52e81e34da4ee436c5593aff65d4a0d0de800baf1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e9b9ab2237e2506095ada82d6219935384578ff3cc82da48d74b63bcb37371bff7126fd747253f7dc184dd163ee3ee1d05101edcd1eae42629d11589883e3dcd33255cef63f8608;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cd5cf53d03b8629b899281d977f8ce6cb0e9bcc5afa0ffbe169b39c08ae2b4378505680309e9d84f4664cf22ba64e2d327174180e9fb950b99cc23a25a9bd854f7c3f3dc6485234;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26885fca70f963f0702e458e30a04b2effd385795512d0bd334ba0dea62264c60c8096de0e46357d187b898b8f5f4ea5b6e35b8905dd0d1c1cf46d9214b9488464f2ef040dd69836;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h226c4e319bf563d1c7f360ff1bf9e1e4b635e0ff056364b5d8660693b2f9adf8faf0fdac3327f162112630b117899a450f4f6be4dac89f28b4ac5048351ddc9e7e8e16a90196060d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4690c0a27a2245e0a045ed3c5eb1b6c2c7b1c617c7fe251f97dd64262a14e2a85f04a29f40dd9afac21ef18a89f7ebde32de2a033397d8e7a898dac43b2cabfb58ea207606be0606;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c5b8f35a1dabbe067cbaba8fe6e7c0fa77d7929052b254fc388bdfe0d8750aea16f5e0fc8d89499fd18959c9820190ed3dcfb611a1365a7aafa530139fc4e7d9a9149941e95b4d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc338694b65c5e0c323be4ba74d2cb5762efd206d62c30729beac27ae81ea2553a81aaad6190b57c4cc58ace2c13f4565bf036cb8410261beb5f77ded09088ad58c2a6938aee8c161;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha17e76c284b7b906f6ad5b453b0bbbc290b20a38af44699d2818c0a4aa7e74c19d9f52e2259a7e89f20d71b8d515a21a7b98e55a3c79b6b281135c9542f2febc3a3ca80f5698e70c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20a107d26c1bca1835a40c82c1fff1cae4cfd94ebad8333615141f6e0760f280906d6adc9fcd46cc72637a1b738bafd4fb955623027731dec378618f17767f632382d9a919747bf6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2edba3b9be537abaa3fc272803fb5681ac528fce5f9c813b1cbf112b327c58acd822f2938a203710e895979f32e7f225945de52e02cf97f403c223422633635bcd8f661855d04aae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87c14f11dd25cadb3fbafb84e5bad924caa97a93f70439ea82c5fa0aa3ca6dd6ca332e91215c44f53fee0ca652a371c5eb39e2eed938b98905b77bad71eb2658fcf131e6ab07da7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7def7a53a62c444a5a563d2172d49eda3944b13c15c41cb68e2c3f0675457e9d0736493bbd1cae4a3e20e8af22d4b94fac4a682bde53e08fcfbb81fb41dfe0c164f67c95b787ff3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h761b7b408147108eed7c1c8c4363818f4b07fe7cf55d637a08cab9eee6f129af37636db5af64cba72177886c78005a2237d833e2c3b3d04d90e5e9e06a449fb0d31086725d9f4a0e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5d23bc815fc81d0240533e47eab78fab1a4093d121e0a26012a8c7952c7bfddff27fdcd0e807e49a498494b79bf45d586686e21e2ecaab885e7e0be1b5a825a839882ed34715460;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4672a714b1335397bc84e700ae30b2fbb07dcf639ff95532ab944627886a5cfb313415cc67645a9004310d441e20a9e851821f0d25b39f58139ebf2f15c6151d081b7a408d4997b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3606e004486001fab6ec08402236dd8861ab059312da6915d6834b1f0853b53a2db67b0ee4428da6442c3c8320a49289433ba1a040bec81eed6c01e0e35a843dcd6f417295ee3e53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4980feb019203b70e4ea4aa7acf0767b581528055010739924276afbd1a5abd2375b6f03b8d8624700ce7fa302c85fd0e77e8b8181c04fc6735189168b2e3770a174df8cebd5eedb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e970fceb95600ea23623e9bb1f264cf0f37a1aef98fc9f0136ee23d20cbd1ed1393c8f1307e52cea8621d60b4220f57ff8299f4304a10702e0969a971943b85bfb93d97f23be584;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4237d4f7f2b200379183f6e11bfd526ce76c4d4f4a320e733595a9f036af42c4f706c234eec0171ccf5a27ca5f694b831e9ab24c2ef8ae3de1eb593cc95d3f607990d79d51aa4475;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80077126f9cce219140461516a708c8aa5e0d4bdc022dad7f00ed09058a7046550bb86918a8b33ffadf94508c2caeb350402396f99d6fb88604f01564a9ffaea23a71d46c54990ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae3730d1042e359b5107a17b7d9bea85db653998c692db98d03ceffe589c6ba8a37e461e80dc03d1de00323cff79ad2c716c48bc451026435a41489ef0b2369f60d1251de15b0655;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23af2533f050380322eeb067ebc96ba07a9963142ab79ef3acfc114ef94db4d9f8ca3da81396c99298e9db483c7e34a8ed8f38858ccab8fc28bb96a9aaedf9e894f858f8e2a3cbac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe4beb568b0d004bf7a60031f09e1c30bfde26b1a7a7bc2344646bd5cff4e73274f31514da4a7334fdb661a09a98746a9afb7e166ea945a7207eb299439964d873167b452fd88e53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heee31928a543c7654136ab2a52e3f1af0c0672ee039d16a16305624d441a5bb3f8977581c6cba277f556977550aa99bca35e10c3e1e366f59297c9346d0d12c1a769dda8c3bb874a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc15348f2cd589455e3da1881f78944a295a00a26f458a4ebe2c94cc5ff52ba4674b23f7c044848987bf68d000c88938115b76a6ac81cc3a3cc2e4088378bf8dc5f050d284df75df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c7f473eeaf28ff820a48a146643d2454ba8922dc28e7804466f95b81e88da52de97754cabe02be260b9303710e33830294ca5616dc6cab62f1980bae5c1a3a2c07e68fe47e69a69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b2ddcc9b5d973928c1c7eaaa7364baefe0d719e52e01ba91829abc8eb7d213ae4f18627ebb7c02260694ecd92adf0f3bd9f69fea5b26352b3c8d795cb03a2f42ca24625303c1eed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3aff42ce3685a0e2ec554f0c2f5909ac66a6f82ddc54b3806b07cdc7b8f201292c9fdd8ec76905f41c2d553dc5f18fcf4fcf2200f81e4c5a03bc12aafad889d04cd87197f0aff06f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12e4d301912030f38f0a1ecf0b239ba2d2727f7edd425c20c0f40d9aea026895bee659b4ab84de4c9ebdfe999bec35f40ac44c6de5df3a4b38c1c24831c4104618615990a486cbe2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4f0ca6fc23681592b7d671de290461fb8a3feaab83abd50386386a85efa5f52a4c411b61c3c0af174c288252e58a25a7c984ec935219fbf0fff4e083d67618e124841e4598853bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e59eed521badb8c99ae6f98c2368bf1c6912406748f50c199d0c3785efb59d093b36952dca59826ad7123994c155ad487b49ce2f405708982e8b86f2f06cc99afcf9c50cccb9a81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a6634b64cbe53c76565af404cf25ea6266618fa5ac80e6a5b243d8740d7fe4402f83f7d4ce08419a29211fa6b3bbb0124d384f908104e7a6304fb5d5bd0f3ff74b18eaf6770493;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4feacc6b4a6ef366e4e46089f5e28bbf841ecc68a0b7f2e1e32875f745442e124046cfd875907adbf254522cfb19dce141e72639e38e58f324563e64558f301c69829617a731ff54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc9d69c647d94079a56eaed7c4d8d79d6ce2013198a3a4b39531d8392b8f26665d7f4faa3a3e2f4f9a687c610207db97b256952fc42490551b1d9dfeaed7f74f4892c4cbe178adc7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56ea06053d3522c7e3bfff5e13d80b6263528bd7d20411332afdc3414c5d1a08678b4c3043dca516415b44242f87e61ef10ad72377f649fd3e416e8810b3e9a1d4aabd0fd61e4274;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c1a716ed1728f463f726ff5ff55098dfb22ebdc7c786061c177e6aa69b4db5e8262ef210c526d20b05956f62b32818427a59bbf48a545caa7ed47fd5bcb12d3aff9dfb53101c9d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80796ae6b1596e06f5d1ab78125e1991f344e17255f8c6731610eb39b157971e4e16d6c111eea4d157faa49a228b9a83f438f56557d3948bbe833f7f41c0c0648185d5dc4d359ab8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcb883e4cfa354f578905b43099ea8a7380db00c1a3a62a4c31d10abcbde52864170514c3b8149a6fb715ca9aa31601b121306f510783a7bb62f91b3dc3fa3c6478111ecb95bb9e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fce45a1668bc0e85095a33755e7909c2e12916bfb9018c29d365f49a26371a86e354b7bcb9d68a9ffd8ee1683292e95823bf44ac92e6e78481025a26421f6a2ca2c5c030fceb602;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6de2eca4ee429a6c02179d71da6480e92251d920094b69f24b47244baf5404ff68530e8350735de164ec91cb0c129f49f386cc9dc46ba104b92a5580b5e1bccf8586bddb107f5881;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he24461d6ac1e2fe1bcc73ddc830845eb9908294f677f59484573c46de2f5351b02d2981ed69241a1c831157080e6d0ab5c3d1af6fe4e7374aecd692359a06454332dcdcb41a3afbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h566fc847684b6d5604fe725775e1c52ce6a9772bcd5c37ad367e3aa7e9b6942b5203adb5de359bf9801d94195226a8b9de0aedaaeae9af802f04f2fa1c76a7d5fa482a8a0fa500fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11f0a57b6e46d2b45f5e7732c442a5283ca6acbbe5c92c29b337044b1a74bf912e89dbb897123d6d5b7da37bdcaa95654a3356e9c5b4d3d8ee156da84cb13c9829395c4dcfb33152;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76fd8f9ee9dd065862cc4f00bc06746ab3361c72ad3446ef4b6c03c35aaedf8b0ee981235d6f2124158129195fe2228cee270dae11f98a3b6fa771afe9c41a571e0a7065cd633816;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6578f053e678c9914c369ef640b3a380944405a73d647b45903126d160d59f27d486d990426716091b918b2423032c7934528fcbd62af7491e86f476350209c224984770d1349bf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha73f4b1c057040dbe2733cd1499f630ddf58b11b3656c911cbe15c80746dd4db6df71ee80c03f3c2e06ff3cf06d83b67520b05c97d2049545b3001f5cc6598d50469885b519cc745;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h806b3ca0cb00f494a7945b97741bfdf2df97a228d8db2bf98fe30b11a5203aef2ae134c98e21f8c56d8278f2c74b92e9a7dc493afdbe69dccd24f37fa46986e4718b881a0a90bf35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0260bda5be84b8206e6ee5ecf0e2698c49f5a430aa370677972386077dd8413b3c27abb8d965fdda382076e31e6fa2c642614030a326d0d7babba6d20678c60d41470d93e7f1e29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1162114f8912a85de4a090b4cbe40e831d887573ad59391a69385472885d03b9addc171f8b2b91048e084be18036dbcaf10c63c217428cad785a2e0f86c070f6033b500e7f0b9fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h771066370a9e86f86c838c16dcddfe58a132d37b3fd8332e23ff19b93d5ce12b31f1635f10b7096d3fedece7bb23cf6b57ddeddb11d27340e3644110635925289ca89a16872c4e6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8944ef1cf4c20d2093f0883dbaf97b613d90ef587cb06fa4a01d431bddadee903734ed4c83168e4098ad9adf8d89dcb0616e29aaea7afc2cebc60f1dd7bb5ca1414ab66e069d77af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbc6081d7cfef5d71e023bf666cf8e6de1475a3e9f5145a9a2076d0de21082507b98cb4b04a82661dd11a3c3d8cd06fab9aac8db49b02cb111f2263ee711f7efbde610202303bcff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44add8eb84fc9f2b72e5600edf36b22c01f5bb8495e0c16b81a52f816753725a7fe214b33f7585759243d3c94f8e3bc48cf626c8921c2bb8eaacc1c8b39ecaebb06b74ac4c50cf6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ded19e8843a5b0725e842708a456ea0ec86e612b5fc2f5bf643f5bf63ddddd20d01986c1cd6827ed421bd4a4ba6f7387517102a4c752ac7f6b294c4bec663442263b5383909a0a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e50b8767aee89f3cc4ff491dc7195357519d6002bde8ee58b9872083262fa5aedaa22add7380078225900eb98e4428ac930abb1d9542dd3987ff6aff38640d370b64a7c4ae4195b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb978f36d342ce3d0fba89fe067699427affa5865e5da556c1a53420dc213fe78f3a4d247362212549979d36688dbebb582592f0b73e03a7e64a654204111c3638d5c321bfcca62f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf78ae6e4d01278afd78fa235bdad308e0b02978fda30e5c70a08b4dcd88f6466e62330b043a68587db8088dd2f6417672a4b22103995a4762304addc284be4dc7471b7cfaff58f77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcda3ba8ec6d6aa1ae7292a3f036f3dfd60dbaa6964311858ffc2773d5abeb8c838e85176202cfff307a488531f52cc57d9d1c676209e2d0aa3c79215f9b9d63d74d7a9dd3d1db494;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b386e1232699c29c5449505869d6512fd064ef2eb1c6ca9cf142d5ecc8a31375b61acfdd8ddbcca20207884cd6f6288f6205be743489509217da8f87e28f2c5a4249f4a60c7f7c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf867a473c84d38e02e3b570bbdb8533dc2ede93a0d8414f995c9715205c200d39e74c3307abd9843930203b6e8ad249606fef090b411217ba5252ed72f8bcfe448c70fa09ee91d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43dcdea02fb2b9d8d1e1a39c897045cbb7c27d3ee99731092af99cc8259d55eb43fe22eabe7c09e26f87907e8f54348333978fc06d46cd3867896f40878e186c01b844461970d874;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he83b085048eedbcaf1bb3c9c63200287e935bda8ba728dd945dc1af39e8ab2d2bb1f311625657654249ae23432c5eb4fea238e9310af216187c5fca3ad70d9879cda0651f86e31a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee8cd23e9b55b92997e4ab62ce356c34c856d12ed39f37c2bce2e321ec30bf4123b7ccffbabab7e3ccc7652d716a59bb77381738143042e1453c5cc15d649fbc77b833d44c9a8347;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h100cdd11d079934e2807a42978d6d98265a9abd4afb50af92e41e16e4bc31d1c4a6a744010d40f488761e32884bc026ce9896c30288f3c658fe33f0a091a136cb039ebe9ccedf3cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcb8c83b8a1895a34ddda6e630a038be6cc5725b805400ccec22145185caba56a3a97deef200b3c75425e8a0c4277a0abc0896e9c7f845a75700e67d5fd8e0e65d7c26eee37d16df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39d8cceede3e3df51f5f5bcfa27b8aaf8124d33eab9b20224a92aa53fae2b27e4661cca8c36254040594d8ec1a528c0536e0bac211a0bf50c1c369f58c95685492c797cdabe9048d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd581bb53c01f3a8632b4f1deec04e2e7c403d70419573b59e297f25cbcde72b3cc10620e2096fa0d7e83c1fbb7b552b078908d017eda8cbe1593d96a7224f746e39bfd59daf626f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6be5f4126eb2b3e3285f1730533159b4c8c3a2619cf3fe8bc359be64b0da08971c16c8c61e1f94423b434b50760190542599cb167dddb65efde2128e70940fb5ab94c3f49b22898c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6ae9786826e48831e1d9ce4a312a62bbc82575547ba54a986fb5400af6d7a0bcfbeaf83b5986a69051596a9f10396d7816570c7ef2dbf7fa2fc5c6f902a1425e99d17da9878cc48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h334cefd7ce0367d2bebefe0294823e97a813150f9e9418220987f4752e9bddba4d7e8b060caa15b27fc16f7800ac4c6ed75301116d6b8c19997c12b8ebda1ede56d3a389585bb332;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90172936cca7a9a571ce703c6967f218582edcb7c39088ed7d1161f458ad9dafc35f0faaf2d1f3d54e5a1569e4cf69f70a62042b561c1bb20cfca029d5977729d29f880435c02529;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46ff316b4eefa598a6296d277f7a0049895539f8ab77883d4443c9283ef6c16a0271e6236d9425f51fb338e81548e9ba82488cd54292d73dd0430f839fc382b51b1df396f9624332;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9488fd1bee9cdd00978e59263d75177b281692448bd6817ad25e4113810ed081cd42ba9b835132b977dd880da5f60ba32d873c638ae8a2ab27dc49638dbe05c3472b0ddf07364921;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83c61c7871d43d3dd5bad58ad7005c00b077bb3069a1404be662bf59663845c872be771b50f62565b5f57f49c4fd665b6c772f09837d5dda2edb67fecb9573a1ca3eea1dce814dc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h117e7c77e8ff75a59bb5dea91100d1b1ef413526a5d47995cbe31ff13b2c5f8c2a40ff50f22b5f0d44949048170501e4452430c31b36ef0621cdf8aee6244186d7271c881212f3f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee9f4ef1e6f45acd5dc1db3445ccb05ad71fa098ab24ab4813eb4f2e4722306025ad59d3f3c1c184d26c799ae3048c42f81d92c882f83af01c7b62389a3e2219625ad4b81de32d0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd216cde4d4f3b4a048605db70385d989a54e0ceeb8550436fd1a7a4e6e54c209e2abb802fb33e0d6d0a5d2daab9a46d9f372c7c35cf6cd7ab443e7b56bb266d8b4005c9245daf6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haae03f605258d9966c39061d35df95aa51aa428e499d9fb27c7d8a7cf7e14f4eed0afd928183258ccffbf80e76a17dad2a18222fb0ea380134acb0933c7cd2840e864dc9e38dc234;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44e52b7f2f28a5b42a7fafcbb9b9469c8cc25ae92a1b7c1536c2be00f8b4ebbc4844b5cebd7375b0e49494221175c5d73c30ae83a097f05a45fed257072c4fecd2981ebb7a2e1a55;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f3bf94a8ba581df8b2cbd69e8762022b849601e2a793bd096abe64b1050b6ec5b1bca428d55936c9f372eb5f0b2afa6d2edf5e014e637e396447b1933fd619e444cbce46017625;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d9e14dcc473f7316b82f1ae15d605f8464e3e50aad3cee5824aea3b982aba50c20ddf44c5bea9f7b7e3cb11a4ab5164f35725619ed225ff82d207a5e1726ab06b6342a68eb521bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b809ccc48597f373d1c00d4678f7da3b9d9b73b5bf10f63450411a7a93d7dafcae00e6769c770f0e3cd2b2537c495f7be7fb1db632c403dc8ad5206fbe428678ae9008222a5fdc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he072f952f1b1f3a3ab70e7566f18cd8560ac9a3c0000b17f3ee0c9acc2c74f50e6d9a735519b03d3d50c5343feb5f0cfd36cbf5cfa6b20508d7d54b9a2755064eead374c6a7e5a9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he49246f15c4fda8086d3efbd89ef3fcabea4714c8e119dd740a66e5eef807b4816868f23267b6801df1c1813cd6a60bdd897f168059adec208db7d5b17ff8711e014f6d8b94b4606;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c030d7f223cdf7eef0f4eb1bef6322f96d08cd357b884b020607d6ecf4599fdc3cd7c94bc6755d961112902c5b6690a8b45446e47e6f3e773bf3a2f7bd0a091d05cfbcffbab49b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h912978b2f4679c66e914778d33ea808b2217d78a0ca315857ce4c4b2fe4d80b16471dccc93d2e7d94ab5b1ef037481069b22919f0e69c0d176b4e6011584d292a9df05e6000d75b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20c0f9e3932e6be424383a5ddf33d24de2bf629f466c454aab08719902713c04cd85d4d5ce4dde9280e4d6f2fa390555196cc37127ac73e559c3c8dc834001b6d7a797f57b843788;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he06558e120cdb8a3d375c4c2e9d3875a842e9267be871efd517a198cf1345c9d0c3ecb57105afd586837c746cde4c2fdb6964f91f8a697978b1c3ae6faf4fc7a9ca86db8a439ff38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f0859e8881b4d81314ada2670953673ee88eb38f6385503d0f9ad153d43a09e4551114095b8de991a2b83ebaaf72e841e78076848eb16a48dcf0f078d99e69c9ed69b3d9263150;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ef8b24c874316ccd4ca8a59b8b56b84d78d680e00bb24583ff24bc4ca5fc9733139308605334e8076fd27e2e0c48a4d030947008026573216286c531cd55cb72efc5250715cb6c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cce53c081402c7c6f5f2c1e357fed0ed1ca7acc5843d94d0a52dc6d59169a0d8e57221a16be5cb636f631951bf1a91ccd88ce8945c6c0e02a6d5418bd88b1ffd145744582fb52a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf18f310d5bdbf5d65f7da3021f2ea97eec3e9c913ac5c4521655b06c099ba29c3ae7a14b80f49825e20f9242774caff8d385d0aa7d0826e6a00ed921624210e65690efc5d2b446f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ea123d91d8435b37836ba0052a20c3d4e0240597ad077b6b6e4cc572d40c338931ca9cc5b85fb65c02eb53d964a188fee763ae90720b4e02a49f47f0edc080de91532fa5299fbc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ee55a2e75111ea6a0f074a90cc623439ba12c42ce46d15061bfbb9cf5d65efab99478db2d1fec73c480d982625a43c0525c7e5983bb467ed607dc06370189ed5292272c8e989d1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e2a11d06c934f21d25a7906f273822e6e45a6f67b1b61d0d5805c8fafba774ca6002dea9fcd6ebc21a3bd76dcecdd0950ab2abded08385da0fba58e9aeef68496e63b82f0761588;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha033b873d1576ac06d12bb97c5787ba65d179ba28560e3eaf3e65ca9c48c85eef3b19b986f1a649703a349e068286f6f716bda09b48d4b1f8b9e83da63336e90c22fdae31ca85a7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4f568efa6cfc3281a1eecb79b381026f686e9b489cbe45fb9deed1d68c294885a242e8590baa00bc6f94ac43bc5cd2cd2f0d2c6e3b92eb32dc028c729fa8297228271e3f8b41922;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66c3941c423ee154daef547580b798ea256ef76944f344f4ce3fe229f3c0026a38a5baf61900ffb8570f3b675be1c3cc965f917e0b1a3a1659a86db0beef7d4b40f6f219387a22d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habc9d3800ba5551b8e052f36b5c3b498e7f1683801a8a52788d97adab720104abdcb1593b690e29d453005f3c46dcc68110ed4dc5f95b23a6733b23f752e5809dd51dbed75333267;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dd52a9cefa237c130f8cf087d7716f2cef5ae8879de73ee2178cff5125bb1d241c97d137aaddf92a4128c52fa2a738d0dda8e93307e57c958338b9978d472e0bd3b27e63317690c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b5c06981ab03e2c5a56ad942aca64547bf2639844224e28f81f185eee844f2cdffa3dc207fb3b4509652389ff6d3d462714735fd2578962658e59748d0ebf65b0e660d692463968;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45ed330434cef51c9c0cd69f25f75e5b15ca54af7b8bbe4e115542b5bebe7a120bae6795b03d7bd28db21e9400c5acbe3b8c88f2d512807b06ef7e30e1f5b70a1d275f60c21d51b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f59e80d21d842a8e4a8c53c675646d09ab6eb805476b86cc9ce1778e26bf5a4f9b28c7a22d97408d58bcd18fa700de649651e820b675091fa7f2cedae776478f1f18720e2d3bd0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1ee8b50c8b4b477b13ac5c5c655f776368c2b64c6ae10c533f34f7236d3451f770fdf85f8cbfe7de775f974f3c26bf009d61fe6067ac6f8b654d139c4864ec8126a2ba3ae6c9aec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdaeb9a6ff17a7e347f2bd347e2c2d945400d3ab86ba049a5d95b357ab6eb532d91289497af5d1d1e5420c1f55643ac25d3dd772b3c1fb3388b209b394cc1a98e691cb395aca25869;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20aa17d14d17c895b62ed8995b84dd12a1abab6fa28f04eb52488619058959c9b3786b7c4e9deb253b59c4941b8be80832eb739ec259c29ada596955c040c0f50d3c6df3985ae4f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3541a791f62742c0b8d0ab49e07132e099adcda2ccb1eb1912c0fb3b8a70f72604c8c9a53a703f0f2ba4a861a138edbf91771c1bbaa78650b7675b1f03c828c14dbd7615b8f730e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdbf8e2b21fa8c7f281577b011b68fd6e7d4c93ab2a1ffcab301f979e6794cb58905e354c354b6d5956fbd0f5383deb34b7a144abe41e1fc18cbe30829d68b846e8588280921e32e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fdca379813bceab469b91c91059d9d99eb22346817e79528daf97f601ae754cbc4c56e70dc410782220648fb52927fd7e9c787fd55d3de0d5868003d917cbabde803c4d5c483992;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3919a6efb4fb5c1d9b77dce8c6274140adce02d2480880c61fd9a903415bc4bca3a46b52034cf9ff827a392884cd2e29a5b816e0fc2544dd9a615fbfc7d66ca4fd0b3c8b56258e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6459905d155ec7c565b2923d6ac740de7f086a26b2753c36591d82b7177929b8c86885ccaa452ebd421f53a7d45767bc358c0127543c617be22b4fe8a9cdae02dcbd08b314592827;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1364da0c5315eef616194a5a79bccce3b441ccfc4eb4f742d36cb392c7b959238d9e95f45061e51219ee4753cdb1aaaf8fb584717ed088771859cd8f85ae13e1e8e602ab5a928b3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h824676702de05c30c46f993ea5007e9a5934037dfced5ae4405f55a714aba21af9ee3091651eb4dff5a205e80d570493806415e55de1c91255139393bb8c89eec190c0d407078d12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7bb483dca267c0f53f1430da550708393eeaf79e746d8ed22f00871d9ac50aa40a85e86afc61f69675f5cb48ee9385712daa402fa1f2ac2131f35e134507b51f70a7b687a7914af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha33fc39820321b76a887602eb6f47b2d6eeeeba6fc3d93efe072663ec89a2bf2e89d5ed1958280cd3c1e3ce0f582510315074659f49159564d3eea39e7f8785af11cdc2257f22313;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53cc5c3ad927300513b2fd715eff7d9bbdc08ea6bc489e0d07e87aefabfd85f01715b5a128b5a2bbb78de7b651bf9f24a6ae2c32738527cbc548d342c84e8e34c6e3470972423ac3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19edd6ef0da3919f34d3284410cb579c3bda265ed33106c40d09a6f543f3040a0d85f607aea0b92c8966b848cd342ce120f4a6b0a92dc62eb20f33617ed17cee5ce6eb3720120ebd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85f616e171ef8ecff981635daa173af28021b15eea44d05f66a506ba50f759224ec779421a6d127c8693958751120568557131a4c25409fabfe1afeb90490639fd70ab5954da32a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef0f9c16bb41907941cad8c67a23a18e31f7272cfe742332933c5af40de9c74258175fb7f00c66d051a3987f1e345ec1fca2dc96abf41070aab752bdc290d94540d492e9ee0d1184;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac8291b1d611aedb4bcf228a854317e0727d779446d0c56a133d34d54bbedcafd814fbe827f3e4b55ca474588ec8381a229703dc48876b5c43092b92aacc066ed5f27dac7a31c443;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d7297b3a421aa216de27c462da539bc16d9799a7a0dd92e39ed209bec5fbddfc81ebaebac59ef0b13bf43e3512922d681a5340b11bbb9bdcef17e0f2e19e20cd35b09d9972c54c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc43c04918285fa1cf557eb8d0479a2342b077cb7a4d862d219144f4243505255b12a1ef9f863f1f716d3445ee11bc5d80b09254ee96a1f2b1b8eaeee1c937a939e1f19b7bab77c0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20349b64ad5031cdb5660bd8a24428e5f1bc292128d5f716e60fba86a452ed2ea0845915575eb4b43f659565ecc123a1a97c61547f8589fc33272cc278dcdcb078c14e1f0e2d944a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ffaec6c61aaa7d177f440810741558ae85579ca717787914d28519c8d6429e8f2af7bf3ca8815d44c5069059db801a3d1e1874b52f6f14f7bc518c7610617e992189d33e362963;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc200af56cc8fbc956423e4d5287ee084b9ff85ea0c047ebd3101c5ed67e1306b92be5ad1783547a2759b4fe480b95f2228f2268799cdf021c6e3300804eea28ae783e722bbea4899;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90ce0eb84d2cb27484143a39bf4faae7c44f87042c5cc6c85e5842a114b755a24cafa1c23012baf065f6c067c61314f5d14958706e1091c3d1dc5c5b98d8513c5309cf0bea2cb229;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe2dca1f91e625f9206298476bfcfdf152e152179b5385032f5c3956765bbd3798d23f0b3661a95716a2fbe4ae9b152e2b9fc14801bb6ce8209333338de6452110bf7596d4ab9235;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5669e0300a4a1e4630ae58fcda7222b8d684e15d772167279356c189963a724539ed78bbed9f5b5c0a9702d7b8594a3a3156349f5efa3d90cbdc5555a7a6b0eca9e9beaa59524570;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2693e8e6edc4e12f6f5866c94fdcb8c13070e777afb7f08e13d7067c061672aa91052027fbc9c0dff07bef504dbb0746473bd0293feaf172ebd59fcf8f756285e7254f8daa3978a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc36ca0f0580c21f937d7bf3706fa31bfad8e4386bc9051d5f2515a6fe0e63ed053c8564f91569836d1fde105a6f3a433470113bbcf1838952abbe22791064424039da62518e19cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc21c5569ce564369fff202c7ba868222d9c3e1bcc91ab0f94965606c8c55a54810a4d3e07abc0c6ac9053c620931904b3c9b41e11fdd2307800001c52123b4c9cc4e2b6fb34d0d78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85c8d57adb14e515f1a8ead90729d95d45f690ef98004e335dd4fdecf596c1124183f040a132dfb74bde4be61d2e1027b697fbcfd3fefbfd3478af8a84623ffe57378d1807eeaaa6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c762f66c280f037ff4f10ebddeb2b68d89ce8b1adcec613c9801ce464a9d9b57388b1194cf93855dc15e97c2465d377bafb1fc21c518a30f5daf392364bf2b2cae6e9c7c27ad67f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19872403cdd27a92ebd16bf9f2beba091eac6ce45596eba5aa282d2167499c0b1eb0a70126f74f6db1bb142c535048f1171dd1b0665b8194e07acc293b5a855cb13bb3ea0373b09b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h334270edb6eaa99026e5a1cf657b1fa8458f11eca9a95cafc4980aac72973a16f1c19e010367d0ce3ec3329cb935d66ec96629dcefea9ec8ae909a27f36df3b6a06d249330541b47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb476b1bb2416167dda0826633de35a5a40b24fd4a20318e2760ae931603713ac859151c59633d1abf65b30933b7a08f7f4cfecaae2ab88dfcd8c3b7249621e85f32f4a699093290;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e0bd4d275515f0a5d0fa15d5e3c3446862fc171e1cb28dec9e6e5ae06066c04181333f5ea048d254ebc107f505aad00335018755f5d67cc9b530409ffd5616b85e71a9768692fdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd1e0a4e0a69b9cb3c4feb71169b039b88086c7b65d3a126a7831214dac7a40b63d359e3f143196579c3beec862cd8c932daef8a04777fd3b99bb8ba09072cc04feca2d91a5d691;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b403d791920b5c6204f7db495dc41b24c7379b0a0cf25289efbf74f3565a1550a39cf83ee9b18044954633c497adc06945642907a629b256a928169bded593fad30646f1207b3a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2d2ec2776f042a64f1bb812dd9e30a86532704d610c83a5c3b0598883568cd4aaefddf288d885042c6caf0b637da706d518c7e66ca43be78271a9b75beded6cbb0f0d18c7cc07a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc14e38058ef50c12dec0e4cfba9b0956eb2a32a09aec8f7ba8f81b5bec4dc072f3c71241d69c4e24ab3f4e10a07c67cf8b46a01bf1accf5d0671352a574c327f9f5af7e25a857648;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h977b12ee5c28b50f543292fd9d0c170b2226c54c4af8ace472f4c5c43e00c82a6d8e486d42a0bb07496eadd2935984a265cb95474c26ab02a22e0b40d99fc72e24d8bc3c8174f0e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h603056fd4c4307c057aefd107c40e3a1bd2c13d6d51f9f9381b8284c4979585942efa68298ecd794076ba912e65dd4b25b22191dee98107deb50c36e6c48815eeff2ee0cdd601130;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd5c8547abacb7bd8b760c2c7fb6253eb45b01c1967fc07651baa2bff1f5c1e5afd9a187a7203ded920a489bb7cf18a483684d8c0b4750fb792fa54185dae646c560a70425419ed9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e3412922f166aca4130a7e2d047f8cf06826660d382b7f52cc04fee6534c42a8c855ba371b924cbfd65e12d5bd63b36405a5442d5d0bdaa2fa66fb1e61f155a9e7d1add6ffa4586;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h524498d70a61c877b9dbe317d7c354342d523f3d86483fae2d299567fe58efb0d0d8f5c635adc821e40f7e0d2f6f1782b52e2a35ab3c4cc47e69cdec7383f4e5b3db74d8de04142e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he75aa4ccf0e032af5279aa4c918a58beb3a2a1654d41b0ca0e62e8159e6668e8e2d50d37d1be2f5535c7436dd717a65271036d84392266e74b9fd5783c84e3c90c1187dabe47bba8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63694d4be1dc4624c14aae387669b8768bd8aa4bd133f487666cd7c212a4090e296ad572e6810fc9e3683255431337e05a0da143bc038af708526ca3a6674f9990f7f0241457f220;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd7a7bd21551655e0fdc32b5284720038b09d54633ee17a2027befec9d5e0804981ab7b7de2e87b3d6a0541c060f7d7e4eba4689895f3db819c299871bdb99e038ac5e42da5aa324;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53ce18f9ecdd236b8f3c2b8bb759a87e4fd8929744438680470969f7bfa576e966fa2c4a5c072b32245b98d1b2fa160a2bfda56f1fb39d1d23a24c5a4d277f4a02b8cb61cc7e7f31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ed102cdeffa502a09b1aaf21f1f8087b685266a58e4dd196c801df164e58225b75f2d38bbb5dd4a77e870ef18f1e27ac141b21241e994592de56deb978faafaba1ab275c7afe846;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5384365a7dc9765d330a1054c85e0689528d9d992b38063d22c7fcada043526ba210c9b0c91fe9d34d345de96db6ef5fdb9004bbaeb75e44e78935ac750674bdfc576dcf4e98b96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8087ca5a7045202070ac44f74bbb7945a7679cfa3d416656dbd737b731b00e87f0f3957bb8e0aa3eb42d98b6ef1248602aee321f40120eefe1a7446877aaab71d56489d9cbd0f44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h385c6d6abf605d017b4cb2c6c2d5027c2223400a16925c510d1b41565ba7becb8b45416f19b980a5ff9750184e593c73c45204cd14535a28ac59cf6e91793aebb27a7304997c0b8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6e520b26249a4cb47a7a18106f2d8e36a01b52fdb8af5bb5dec5f669aa707e2627ae1e1590e683005f1d3fdf749ed462626e278e244117ae26a983a730d407e78faabf488db7b59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f9c68ae0a06287fb5a03fffd86db9e3aede553f904ac90bfc0ce1e4445b0d658e52d5675c86475c344c9dd651d8893cf23fd007f99df4d78309b741947fa082ae21c28878cfe327;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h443b43722bed63f743f3f66cf65968132a381adf54de0c02944a0c4371076ac610aa6a75c9a7b6c82868c73e5df23d1fa045ccb277f27dd21eb435cba731666e003058599c29896;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2887be1b978c4207ad24316dfeacd159a0822c51148a74fe202722d2da59032ed843f53f25522eaedd1909f44405e0bea43e4660275b0941897e48c842ca72dab0394c879ae45749;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd74a1c2484bdc23c9fbbc87bae95c71afdf6f425376ce80fa7da46cb0661533b5b2a372a6623f979a37a2f94cb1b305bc243c1bac8d05279081818c03b05e43b0ef18c6ed724ec92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cb25512107ebd5f4b1b2e56bf36b35f5c19e1729a3877743ebc4fb7299d4b31ee3caa072b315f53db4b3b08c0584f099736062057732733d64ea27c5003021511d99f40328a2adb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51082afcaf6fc838be5e139715381b93c0a063b279674a480757a2c7fe5a984365231d4ef0d65961e7349c08168de28d434ff664568f00e760f2274b7fae5b9328d6b6081264dea8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h800f010373d08a2ad4fec1a4fbeb680895ce32f90d5ef0010f5ecc289fe4c5f38de88e974d5063384deb944123ae5c7e2ed0cbba8fd87c84b181a7ea51ade9335bcb289edf262c4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h342af048ab1bf2c52314600ad676e99fe2db83c96f40539b24db8b5fc6cc451a3a0d7bfd4664b3dc662b6ee95c7e1f10eb7420e59bf4da978f350d405b8beffcd9e3a8e234387cc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1415fbbf932572df76ca5b49dd8ce8b5324362aa91f67b775c6578c1c2f048db817c3009489ea83b4066983b2a5cd863fbf4773b7113cba3487ebd030fc1095ac36697394fbff637;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1001a68a3f6e7796f0154052fc4888dd1b119d9fb5b0246cf5ea0585b38cf9b56d86026f22953ad18deab6d4bcd299572fa41cff4b26eed68149e2eac7816ea0355450cc3183531;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ceab35b24def33e9f8a3d7f7baa91461adcaa389a80b86fb2f64acab13cd1bb3ab0183cd4332b7f5089761b5bcb5006a90f2c136dedaf88f51b97e0e34d9b3f8707480e270419a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6af3805f8d229018f392aa3372f001bcfdbf71f2a576bae59209e810b051fd857a87107c72ca219fc9faccd81badbd1178d165b3b48d5ad2ea9180d86a69fb02bf08afcdfa9573a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a4c5ca937e8bfdf1f1c3c0f276995610544e970f865f820a3e88d24a770196ea2ed8f022f63224e1cb27550646134537f54b40537c45b553ae39d7fd2643d04f9f97eee985a70fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1860ee6c5df62011a2408cd00520d6946affc0cb04e6bf8fbc51cc63379f7c6e957d6f67470949a56dd901c6db1ceaeee539333017341046934aa0a83401837ab0eafcd6ba6e21d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h386a09f0e3b8a816ef22d7fcd5c878ac30ff56121aec1f6d328f41fa19997842fe9db00f2db434fb632345b16fb35fbeaeb5b60194fd7c10695b6331cf8dfa591dabe77789d7225c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2dbc9cac8044903db5e9555ff0dbb804e103a097be6fe4e468bbbb05f093ee672d6b91f8e1ed442de6961a84c030b3314664cf56bf8b7263de1da4483741babe11cd8ee8adaba096;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8ab2b0b1c56a452319624a5c7e32a47b3db30987b8e6629fd8e0313df438fa8d22ac74ce371437b0b45f348b1f1e9aa710c912113dcbbd3d29b892b892e249737caa92bcbd0931d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f74ea013ef9284de53830e114c80e47150bbf8e8ddbe08d26cd436daa5fe296c090066abb3143d291ef42cb14cf717f664470e33b738c2fc31d1a096476a845520aedf45b4e43c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18948326287f035d1f2ddcc65820a78c5e844ff85e1f1202d1e2731f5a361236d78ec7f0efc15bcd84ccb8cfbc58ba57da10164487be8c593977d78cc400ae02f4eea34f3e066b50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a3fe553b446221b5dc34750f79424ac5f8f16a23a874b6e68e075d5854989dcd5ddafcf060ad31d7e6b131969c1f61cd0dc6049d664509ae4c69f635f1526a093d5e4f8d93db661;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb2ad7ebaad34b7e354485c4176464d4489cb8649dedc74f3fdeb25f5361552d0c76ac5e67dc2f51d0e12b4f3477af57837cbac3ddd8a712fcd3d3f9286fcdb930304ef72f9009c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc51aaf29eaa3d6f119a72e6c40d2481dab5841511937b9662dff74d0dddefb88531130b453903e567bda463ca3b963408854f491605f1f8236d4473321592b96d6e91a067474984;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9c3be0a72a790307839cc78fc803ca11bbf2eadc4e15e10be2856e3a5f277bf3da14045f61e4f716fe53e1dfd629fbfa6b7092a965a51704d9248d9f0571bd0d984d7fdf00f9a4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a9001813a1b2123a23be2ea7d55c26cbbc8c9db8cbcfa6b5287f9ea50cced7f291a9cf2850c6e204d6bf7a0f0046240ee261e06bbc494d74e4be005669bc31692cc336e732c16dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a68e39ebd57f179473d6599e53b8e7dc5b8c1735164625463bd2bfacb0c169cd15a8961c1e5c79b34ec9951562e9466fd94ac1610470d01043195c7446ecb5bc2c280f41e829863;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h249ce0c5fa8e84c35912608887b61fdf42ee9c6aed7a06d8cd00eca9bdf15a3eb673857f021485f5e1f8f14ffa269aae3cf4063b74ee76b3c90f3c3c6a23a95e5827d95648e6a1b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4df0b61176d0c2062e8c1418717c92d3ef89e8f68468f3d05eab718eb9b888742e29add79951d3ed7bfb112f68d00f5d7881ac84508b9e0fefed5cd5f3635eb97579ab8a0734b860;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h421d86215f9344ed4fb8a34c3a576983a1a1211569c6383ffa1003f772908fda9544332361ea3cd73f623785ac703791c38468aae6b31049100fdc72cf93415371644cd33d1d5e4c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55fb08662a1b47d864ccb088b01f95e3785e685b4b62bfdd3c92c5f80a263d3ea60995277e8d0e063fced6acbc040e9ad37ea5b244c8cd1db3209e9278cfc5ebedfadbb431011420;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h807600907ce490b4cfdb306374e978017165e50c1a7a5e8e7a551c59add2908017edd22185b7a11c42bf4536b6293cb77887f413e0663c9ccf9e633f756775c8d77ce6bb534ff71d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84144cbabccab547417c03513fcd0fe1d89cba2de7e1eacaa23ac61c32d4565138701abea0259e728e068d77c351460e735de92e15c298b0521b3169e5dbc812367394ea8429f2cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4939ab821994b217656464daff87a1960278c9d9ed6ff065f00d4772d32926cc3bc5463b48cc051bc63d15d4d55942950fd87135a45598a178d0b8b71503017f158cc3087ada73ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha20f6fb56a0843817d401c28f713333f2f6d7c816c62e28a7592db4e15236c0cc3c6b0d8b533deb78df9f53f6d8cdc4823e7e3ac3641b0c22029af7353d6ecc397326c5d83ce8c12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc18658ad221a407ec60b40347e40c13c11aa7fc3a9012e76477d1d59311868b75bd8c38b88612bbb21c1e46ba27e32acae23a4d8ccf7ae7d0cb4204c098bfe37d177b2812618e1f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he380776c77cd99eaa1a375374b49d9c08cb9d4d7a23b8418da5dc87c831cc1bf0a2424de7cc39bb7349a04eddeae43320a871abfa59090dea754214d4eb1f324d544d73a60bcff1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f4b2a71ab1ccdeacb954efe0c78305d1c8ff79513edd9376370963c335b9c46b9525df6fb673cb2179f28a264561ffb75b2f6462d3fdfd0d1611e93b0116342c80d53699d2852ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h760978193105823c566c8538f005832f12e0337488282d85040a2c30a62a67a73a1f1d74ead8c9b4ce2b8adefe580877bffd84184615bb69dd7af06b4223c3903f54bcfd559d3597;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81201289e4c016415b23a4975c3e9e9b56d21b5f73b36730596b5dc77698660d8874b03a1194b24ecf225bb4663a2d3b5cdb181559aeac32fe4e9a5374188ceb3ee5dd900047d2fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b07c7166cc26366075a440cfcce7b20f412dba3159b3228363bc7b4be747a436a82ac1a1f196598c041fe79789df2b45e8afdad97c9c25ac3a89c04849fb46904637d29579a4df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ab4b46abbf3b47d63b959027e6e62f7cebaae10a23ab55ba6ddae8af3658563fc9e264c98cc57e2a329ef2cb5f40545c6fe42fe22e5a3f0f872951e6f8fa2c97189e4656daff213;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf307737817271241cfbe74a213cd876da592b276150085972ed72cc8635f786e6ca0855718b6a3dc20b51458a310b0943e01558775e7c63b8ec344f8b78d271290fa09e6a15b6e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2925b5e7eaa60cc0d9306846c013923a4fa4ad7f3dc3bdb253fbdec12e94382b38c14ad470f70a39f0576b82347406a1dc2850939bdf28324632330a48e21acd4c4cc4bb76c68858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31eb12c9dbd8b9fdcd2375f6896be64ac59e13dbba0fbf5e234f3aafbc25eba8756565b2b41bf86705bf7db1f9915edab5200d4faa6cd93b9db0e0502bea54aa8b5f959e3dfae5a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67ff6796bddf48bb643762fe804cd7662df5301f424787376d5b53f3cea28e99642f245ef9877af9504bd06b105aa589e463a2c719499cfc986469af0c0d6307e3392c43a2e47e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9e44b022937331d962670dd7bc26cf39d7abd85644e95d002294c0486ec83e572df3bcf917f698bb01fba2a2e653ce8c060929a449a89cd5f5e5c5f24a38b4314decbb05cb6d70d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6abb96ec43c12d124a40ff94b8291152bdc0f740ce338d9f60ee7860b4e97749e61e3ef2137189bd95f479a5ce333002cf7205a469c6ba6974396ae520470445e27894c9ef0ca88d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5f4afb7ec95d98e84fc996aea6ae16f9ce20d222d265d8cb75df2845bfbbdf5466c4ee7fa836bfe0e2d240e54ec6150ddd98850dcee3412d8ce387dabd14877d38c29cb2f4c3820;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8408de5e81ea7444112b483e0e0280cc74f5e6f268e0d199fde7b920f7d7e08dc7cc4b72fdbe576d464fddde17bb33a4e28f22014acb74c7a3059add759c75e791bef1db01f146f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a6161fd2bc7698bc012198e5e7d7e534493bd3dcc8c24a41800db576335d08ab3c518b8c89da107070e59e708663b7b5b5d441173f82d20400e919f9a5806705037e8cafb35a1b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3cc40cd8ffbd8b604be0e43f61392e11a5b4fc718964a5aec36d84f27d6aff92c662fa745c0d66c7147f9ea86aa3bbc5b1a9a9ff37ef757efee325f81c37b41aa0ac377cbd897b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d822dbf0424df57e231011a1822e238f659221a0c9b3f173112fa7462b4ef874f1280078c72ca6c00233c58d99085486b2e97423d7dee56f62ce99f396a01a049a4888831ae04e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he16f19ac675bfaa8b069d48f52d4b84039e65758db92d8619e44ffa502e8f9f06959ae49f95999d3734303506eda42ca6d45bf99b2b703a46248f7c3b942d54643e5890ce5df5f96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd00d4fa4a30e9c7659cccad4016ec92e4808a90749988ef7ffcc93d443eeda879a233633600a214021f3b4687e854eac90ba0c1de7a9e08f78b7d46d9b647fddc0886100d58c485a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7536aae6e761abb33f2a75fe3aeb8e1aef45e43456dcc9d5e88ec8e13715b3b0562c77ff679796829d77ab71ddc229de507a62c3a8991e79d94fdd1c7b1d6b2709a87ce9a9e95127;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5211324fc030683c2a4437bfdeb512b8e0eeeb08ce256bad7d7dab5536e1ba6c2a1815f8943347b79405f86563852f1270794f3acd3b3fdfb2fafdfc4df9346fc52591d83718af8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68c4180bb868fc8b2666dfc473959de8f0afd51874113b61c5951c1a6e165f4070b0a1452a1c44fa5d90ea294952c98d425569cbe8b5c95bcff2b9227b8f330edf91f1ccf55b05d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59060edee8c28c994e88780443f5f9a0b37017ad29aa8f9553b029a9a9e2a7d907b80a49819954cb123e31a5a332277b18060c7ea9c1e8eed471967b2cf344dc22202eb0d4fd8dcc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94b4e4636d62aa2f4f7595a7c533471572fcf72d70a10c2e7c2020aedb6a77724fe8cf07fc56c81d88475966d46573d3905f7554ce75ba3f99e12588bb5f4e1ca29763455785cbd0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf84fb2f0d53b877f0dab44ec7caad536080d9dc21126522e9e6da5c4b3feb2f68d7481fc3b25a9ce1fc91b82449047566c85f77a38deb0b949d57f48e3952f80a1ed84ae642609b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7d90a0570d6a682d20fbf1468f899c4452f986d465d5c5250111097da78faa6cbace5ebfaceb5a2248e91f41888900df51ac123154bebc52fb85dcc1e4d8086058467d6d1f455a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde50945e40c0ec0418a598a242dd0a9f4683b73ba2ab2f094400c1a2f48abf76570a633d04da37933d2a6e5e7a3ddee1ee41dcd0da19b155a0ce20c95701c2fcae3372837c3dcf47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h811e0938bc55330d5117facf6ec342e6df75a40b56736399effaabd0a368e34b1064ed3a4a26ccd1c159a7ca0d80da60ab100fbc1177958fe0e3ae673b4bdc8e9d9b37829a5f0718;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd9216318ea98166d451490f063c9ce616444658cb4124b9d9d20da4ae637de393be06a339c0375c872c61dcb95f97479c0e7eda304e9bba149a0b4410f06d92c14ffef6b76dbba8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19b8b69d83b11bd5d66ec72484d2f38c5e9a9e039fb44b2b7ab5535c29f274291b64cb3c251091f5c8ed7ba296ad7af17d23cc4d3690cb302b277323398b9fbd831fe866385035c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39572ec36eb466005a5493778b5a20f6af8e4f9805608bb871ce96d31bd86271d6431de9f3ac5f94724dcb8767d9745d6d4a77a85401d8e8dca6b07fd658663a090a576eebd89ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h277e438bd98adc5773904c7f05bc737a65ed475362c7147c418cce4405012935f7046ef2649af1fe5c7a702df6ea655e4aa1615373bc25fcca7c94d3105ea8a12b45933af590c33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he89e53f2af997c42e00d5d303440924af77d116a31dd80ae1ef4e69191bb612af4ff59944c3bb1669320e80b10f42dab798d567b36057b22e5ec9a192130e9de61ce79d76e30c60c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb0547b1177495adf4924192af57982c42f5097db886bb826eb02b8d4085de66ed5cd91bfde5b24ff4610f509087018598304dd1665c956ef35a74208cb91eda19a30321feebe7f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h195679bb714da6f1f008b06a9d4ace3c6085fc6071e2cd4195e93b08dab4556eb6b82b4948052e0d1c02479aadfd055f25eab98318b65b5708510b1b05d9bb17aaef6ec97066505f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77ecb3a5ea57c153a5befd6f0f2d06c6110333856a5ea0cba597832f15780e343ed448430e9c1bc9b69f5aab2ebc2bb4377ec6719c9281d2c8797735fcac33bc0177ffe05fa0b099;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h613517d8705d7f3884134bcbcad3ae778f3555ae32af36493422d7572f1a4f2c9c3ed1687e98c2428429d001eb102acc848b8f96f0274175b9fe29aa3896df53e62b47c5c490d8a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0668d3b8347bacc050265539b6d1e7e12533e0fd5ae21a51d47fbf8f92256b5b79101ae8f96f1be8b3b0027191489d8a7459a8c7c2ce139862fcf0a6d079bbfbef26c7f9f08ec6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e23c83230cc6a9fd6f089958ecb764ee575cdb57026932fc44daa5378816560bf4ec4fa9b446797bb8fae0a284c41f2d012df35c1f481b0f1fee769f69041015628554093d60b5f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h374f03d40d82767f2050f4ce7de8731f5777e05307a453ed3e4b8a15d0bdb7d565d8207e50abf741607cc98aa8e5875fc62fb924472d164c8833b2fc4d46f9a3498727676622d4d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha30456883b55497f0db284a68861ab3f956bba73629b29bf3dff838a159df8256573d9a8102424594227ad0fd68c9f0df0164dda2589f33821c7c8c727ddbb24df468a8d3fd8acc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h548acb27a7817ac1e79e70a4e78b9d77719091907a8e22d173306d582936d072ac8980c27b1ffde3b851331da004c6adf101194b74c42f98228d3d7325ef236d4a81581ddfa3bb9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ae30470bad571d5445e0ac0d23bade9c75bd3507d810fe882272d0aeb545cd5f164f84795cd9d7e32bc263958de8bc8879a8179cd49fb5ae099e1b4dd9cf4a7c74b5b768548f83f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h515adc6d017d2049f2ff27d9d8bdf82b5650c62b2d2130a95aca32d4d5923122a8ee3c9113560c6dede9de2ac76a20b1f2ec2f15b20ed303ee283b3161dd091018d5314079d073f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6b3d0c86ff8aabcc06f0b64272ee0aa23b4d0789ceffd63d8e4d597a98af5692bb4bf47d7aa27e6e4524a982dfccb55d0c6e44116773f80ae436b8ccd8b6a9e798be67f1860f8b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbc6285c6fa765f5b5f165a8528e61110a9413dc8d0088426b0a3de20e6b55888424c8ef0fcbcebf96cdaa24362c6cc694984759668cc8ef806640c13e625471a0e6e2899d93d7a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h913796b65ad4c4d009b1a21bfa81c70d4f1057058e82eab0672859176ae3f4aabac597c293f99c8b6a7cf9df80f1b429b4243ab2300c6d5226ac8361b5078142f45ccb5cdbc3fdfb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had43100952be6430b27560668a915a9310e0fba05c2a5c061bd7fd23719d9164a4932fc662e965b466b2a644b89d55a996499963a7bb8fa39df84ced04750eaed5eaa1e72b5f3257;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95795283b937312b8e9a562ad6de419ab88ccf64ae508338f0d2007c93a7ba0fbb11cf8dc54dce5d8d51081b9e9b69eea39394aad39ff196ac676bb7a33c7b4c82b701995d1cd39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd61d17d2594f444d4dde2ff54bb26ba229f794165cb5682d9e8f554ce6c692a36fe41d4b48c10b352dd6e147acf0a57e468e267e33b649ec3e1f67c1deb7216ea57ea12aa8b3b03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3c81b04969de6e76fa496d2e9e00b8c32f778a821d3ad6160f31f7a216bb0a0685ec1b7f8cdf099eac75f530b76b954fc03b9e631617076b13aa72b7d91380aa468849a9ef5e030;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfacb00c9236b0027dd6543bdc79ebff77dee5d0ac38604edde3e9be5d1d62614889cb3d3393ced8be72156fcb193051ea1a7558c0c3b006011647be7303e586f22b4f9fc07dc64d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d9a81c4a7bfa40bdfe9eb881874d0e06aa44cc51e64b19087a4862132c7b7fe6ee745827eae162fe3a743967c64753b7161238ff0f3878231318cb1129e467398ff53d3957ec703;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9494d8f90011ceab6b8169d6a4db7b4be832ff1a1ad31ae2e81562302135e9adbac8afe2ac31bb6eef9f42622b8d28e82fe936538f276b43673c8e1d938b8be0bdfbb9873af24939;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bf4307d7cf5a043b9070390da117e20bf0825e5681033374b9aed0e8cac580bbe4c0fdbc09b18f88119cebab4da4e1d3ac75272b2612b9251e2fe914aecb3f0501898e0f27aa298;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf61dadcf01e78c9cd610c7c8151484cbc4412c3eb5854f888d3f9c3eb068ad47ca2337c017c990daee8e4bde2f0b05d732a63f6074312aa67b41cc3adb90d64a1dd8c263eba66ccc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcbc96cdadd6d3c3bf5b9ce944957e58d7100ae0e7462df3c8160b263c1ade11561a70503ddb8eeefd49c2fc1267e71c6c4cffbd731dd94c7c9307aef4d32742a8d6f30aff5999c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43ef6e62c813081d49b0307f17ab4d2bc4a7c26f326095455ebb2bc4dc4b6333a228174ef3bd485f7705e2e64d2fc12ae2cbe51cf20e9b7ecc2d27c42b56c95e26c1e948c1db863d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25c1b462c79e9ceb8326917206e89235ef979e922f37d7a76095318842cc6d4027bd29e73e2479b0bddd70b90b3a118536823b06124b6779cd4f702e57201a061add5cbd0c00b4ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h340a1324bd2f4ef224f42839063c540de653648dc3f83ebd9b4ddca9a5c1095fa7adba961e8eaf767c49544aebbc380245b1ee1d60ff21be94efd2f21121ef4dcb7df0f207deabea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc26dbe1015c66fc9a54dd3a5e43ff07071e10c2ccf29c53a40ce26c66c15deab8ece71f9fbbd0b5324d4b25722820ae060b4cc6f38c4707c563fbf3fda405b5fb601f943906945c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc68795fe1083d85a47e02d8ede7a08ac9b4504588e70de0b64d0682c8d7469c675c8b6916923470d8ffd1869033c087a7482cccd178d712fb3401b11d04acdc494e4d1fd308664c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a786a290776d1b5584ef13a1936f3f01c01c6aa32575257631ab560dc58f4b168a75a953060170d0f27fee088e61fd398423a18424efd51c6e43502724ab568497a1dcec55e1c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc568cde33dfdfe67b69b4d0a1186efb360de90ed9ab6ad80045820c7ef196aa494599ee22cc4358070d838042a923f83ec227aecea86ad4b836f98ae381b4dc928e8efdaae0a9536;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fc887ecd6ee5c1b5decfa0ec7413c5c0f92138b9994768b6e1fc869df6d223728fefdefe3d66ee97007bbcb42aa2f59fcbe67ffda2f58c22c2a51dc801e427fc30da35ce6561fdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heced3261ec634dda555adc1c60e4b4056388e3d09d10cbf9777c83ea3194220499ec12be26b8d760da564f422fa70bbdc4582926f23aef9658dfb2c5bf9773fc121312053cbca0ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1296f23b798b18a4440294763fbb99d05579eaaa5fe9032d7d93e953b25860c11632e735cde9a4b84c03625393294eb03308cf106131347690c08daaa37e76260967222d0e36ee10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a81c5122ee3cc3f2d0ec5a2ab175794791980033c66c3b9474492298fb333fdf9300f8be6ddf013f5b0005af8b17c8db3ccfff02f79a81d671e8aa26d90a43265f64579654e213c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5afb9b996ddadf8de7235009af6b87a0f313830faef3a2d6b4b258ae5938b6fad96eee8da584602dafdf85b791afae792146eaa261b419840cd452ab10a7b3edd4b76a1999d52a81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ed2fcb7897af6f01ba7da9e69b9907be4f23da42968e86a366df2ff43721854c2e2e14c4fca653c5fa392cb18e30c01cd6f250aa96a92408a90b5df186c530953400d60e7cff319;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb108ab51b940471269e109aaa4e0ba4d00c39f32eff001c2f9c80fcc48d47c15a9727d1c5008d12fcb25cd2385877fcd832569635f784db7f47c499f42e1a8795d25e0aac84af9a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h432bc3c905dd860820b619640b93ee32ee7d120bf650f26749af3a314815e76c551b959254ec5b502acb59ca454f070a0c912e09a7d62fc33df6e8d8b2e4bbbbea4f72a472a76a06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e3d55a17a7dc565e23e2e622e18dcf279c6648e48546e9d2f64cee6609806d1e366f210d3614eca58aac7b6dfb9f85beebdfc6647c8be5e1b595563f692305bc167cd82e33d901d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88242468742a1dbc1fce85317b3d0204713842aacfc088ea51ecad2b198a92c7731f8b38087cae974a43cc0e0a4d9fe0923604ca142e74c8d46c697413e1747ca026b04400e8e677;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe40247c4682b514daf6af6fd8ed3274c86d44c62447c287018f3c13de9cb7b0a9f7b5fa87a8c00ac96c4afda40179bca793261672e5c5a2b9f0ccaa41adadf324df0b948d4d47f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc13d5a1f4040d868f42e2d973e83a2d78e48b6ca3404117be8d4e174296704f39564199ba46e60856192d634776380378f00b40c8776533129fa63c3d4b3ff1cee093a75b311668c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91272455298ef9ae0bba3d3c07c0ee6b5c45634f796b7ea392cac5feb4f6acb10b536577c19c4185c3adda5f4ad6891b59364efbe71d8ce97ce9cee45ecee4673b5cf0b7a948537a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94c5f33a30649b24aa9dc55ad364f7f41bb5b017fc5296121043feac18adda0726eaeaf8a4ed9f30bc6e719728605896c5b5f43c2989dc3e9f21848531a7166b635c6b9825d01051;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a81003ee3c90be76ae3385c22be98ad2470967ec3565154eac7f711edb1b36ebcaf185f219d42a35e2094ff5075ac5e3cb633619f703395dfeff1d27b522a248b6eec2b12ac1da4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb6b87ac376446b6cc5db1b033ab2f54aaec95bff670260c49a89c0baa85d1e174c8f0c9f58ebdfbd8d9874a195a21be34f8c1b07854f373e1002037be493ed96c86f83706fb5458;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25e8400dd49caa4b964abbff03ed485f1da6bac02ea9062624b37e1b75f64e459bf4b256024817307e41c6e026ed1b3a56051e382fc4e83603f886a3a56ed090bd5c7e9a1cd6efa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha167321fe4381212c201bb8efeaffa76d085116009766259bdad22f6ccaaa11dc5c8230fd3839ac191bc9e5b4e6aa32277b4b459668df2535b8fa90d7cb14b3dc3578d1fb9d800eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1b060c6dbd7f54f664d1820da77ffe03363929e7a96aab71f10d84f9925c777323df6aa99019a3bb65ec4a8dc742d8239dfcecf181acbe1abfff8ca2b2a4430f8826422a29d1678;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h407a9261ce9fbf75e0a6e61da837895f850ea08c70c82e2cf4e2bdf2e8adbb2faf6482da6c80190bd04a5dda335c433e024fd96907ea5e65fb245d2bd736ee92a28f523022987e0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e5886eff7714f2eb960abc43eb07d0e922d9ea02fb55d9e5d2c8520aa58be78acbeeab924cc1e211323a14827ae606531894905a3b18027efc469eba669e546d96660725fb731dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b4a87af34b9d1d53afeebd8932f6276af5bad75181f62271bf3e25e90b9dfad6890dfcbff02a1a3786ed128b188353b009337fec5ae77cd47780d5e0c7f1bc5f1abe8f706b59ce6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6e883c71e53884960b68a17a473cde82656a80f3fd91b0df2cd641f0813205d334ecd026cea27e4e2065cc17a97d63c91b6a455781838b63dfc6d6c2ae15e4e2f66c0ced6493f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8349cd811d873de043432095e7792dd65665ba22fc8f21eb07a87374120095c7c09a98f693baa8983ba9f07d8a219b5daf1513ff77b46073040d8d78aa28c69647d97c5becb3a64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23f3671d0e593f7e27c373be9cbc2463ac9c1332cb0f26ed49cf0a184f8f0458eac9dbcc4289b9e0bb6fca29ea3f8440e847cd6fff329632967257eeaad7187e78d52dd558a9bb1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h471dc173dfd1ec7e72f64ad9e5b68d1432f666ec042119972829663e130de43030db605f4de788e7267bcc94fb374a9bd097bae5457e99e2c3c1a9ab497da507042c8da6a9177f4c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc00a93482e2f28dbd171084e819bed073ccd158697c81d2e584bdf9f19fd21363527d2492ae6f46fa48ce2a452d38c3a790f27391930fb2a47c077a33f4bac3e2024ef050d1a0c09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18ee6ea9d120c33153f896024a591270cc2887c8995cf2a7e222313e5229af2e6a9846997a30a18f236e208d0a9a62ee931b7883a3ef40386344473569b3540e9d106c228dcc828e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7defdb04ac8fcb113a63c7f9f11aa4735ab1efe2855b55fd84de5fe1fdde381186e27058195ac8f7f5a1f311e51767b189a6d66d2dcd57a48720e2989f36f3ae79e890f80f1c70df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87d3510a2a1668e54a8585b85e738c326d9f39673f86c712c7f5d18c61bca7ac1209e3f5484174a0e3e082afbd0a9db3b0d01acdfd48441106c612580585b02889a1d54f9af69e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h332342e3027b9378c6bcc86320bfac28286e7ed4cc8c18218516553125e320aede02df3ae9663184cf1b8ae91b2bb67961c3cf9c31476214a3335bc7f3733242155ffcc3ad571bb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1308fb7197f2118cb394f60b1a8509fe622fd9f958eb72f1d0ff027d65966a977d13179dc6b3f277e66eff579a7bb0691470cf859a6ef5bdb59c7fc3b1c8d48b65eb407d0ee6e54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h335e5a8047dff53e03f0aa8ebefc5466b298db11851807420e87682d3fc904d6b89f4193462faa3109c5164824f5a123fa4a7c5480af43fd045d6e15db53866a953f9d84e81fb645;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b13a7b422146e195977f17ecaabde096611de0985dcab75dda3fc4ce562ffa933d82f2c5237f0d1e404c86401ae592c4df263a8c5b474b24877459ab7552344d79d00695af4cdd2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e4ca46559cd2cd0ad07d9e69dade438ed2c77ea12023efdd28f4b27329e735c5982727db5caef1eef385f826de464cf04083ec4229181249d5df0fa3bc940b1d4096070ce2e7b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdc78c52462de9072a5c6fdcf2424945f4f4e8a89f1c5fb6cb873f6b7c55624ae10a4fb91be427f72f7b568edfd42b1a84384dc2ae99f3c3dd51000202423987d1e501b9263b2124;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h820283b432cb3c2741ee89daff5b434861d6f1c1c21a5dd9691933294e86f2eb13df31eadd0de962f3e83478c2103e446b16b159d72ce90035e5af699fd060647e6b996160d3df98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h845355923798afdee44c28ec2cd1544c13542f487c23f075ba0d3b3bcce3f6ff2ba6048cbf01b0df7a3230203521c955018cedf9d35e0981c207e22af8eb34279a09661390178af5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1de3b857edb9bd4c203e613349062c5002c654d2e3a275f305384d969cd7c91fbc86dbb1b263017ffc9fb7937ecb417847b94408cec0eb80aa5cae09446b77e4c7bff05d563e425;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h942f21e73b1283ef326135608c3414e8682028cd6216e76ab0e5b1b348ee626a79f0f1ccc0a6ca8fe31faf4a058c86294662c706ccd6d68405a870c8d6cd7b7da5eabcc9d37260db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77daea3836a17d5b764706336f275ddf3e279d6a70d0b1f47fd7f7a0a775e2b607625ef98c8d3eb93d6671ef329eb6cc5c48f6424eae55cb35a6449d392408066a1426fa09109c33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1168986b9f1237ea8f7ffd90dd0cc19bc2e9d85b1b2651bff608f5f429e96377a87fe477f557498fef14761af4a8cf4f92470f90a12c2d50fcfe95b06294f1c8907f009ef5a1c9c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha00f73c8875179593420a6935232b975ef3c659225cfe74689dd5783836aab9256a250759cead578a1b712f480dced7fe79f8733baa75c91dddcfb6b972acfefdb3d29a65d7da5b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha625124bc5195ee29484663fcc550a3bdb3daf26f394529ffcd4db4c42ed99b406c1b2b5a4a011d5a692eb9c44d7e0f94947f8ca417f9e1fa858b70ac98ae9ece24645dc66859e75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b0fdd8640c7abbbeb2892275149ac9a517596279df67cdeff763f1b2aad9a7047840da6dfc67e1c43189979be2510d7ee21a6bae8a611b2da2501401ec83d9f6d9c3bf4a8b0b67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e03fe5dcee0a7892ce3861cb55f0cb6a86c23812fcb98e0bceb06be15e5b2d9ba4bc65ac5a3cb8e9d515af0c9779d3534d9626ca15a2432a41beb167115ed239fc8ca3f575955be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h998ea73d7964e0d980be0d9c36f7375fbb92b6de4af2deca2dd3bea37c545411e1c4c9144729a1efc142e91815aa591e9a24b458f96a083713a43b3da99f0cba6e708192561ce017;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34ec192b6721bf825e728eaf07741857b33825b81b312d22d06f424855aa19d60c63ef4181921773bb1a1493834dd1a7a5b1d1369042473bc1b0ceee002377d6cdd27820de305762;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10911d1209def5b7a3e4c197c80fa6dab2071a5ccf0a9ea30ab139731cf4e5d247521e1a9ff86642b9cdb4a865c3bfcd8e9b336ef1c6bdec12a1b4b98b236e0345d395b0feb614d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f2cefcc5cc287277153c7a4a94a5aead20dd229abc30daf054fb994247d5188bb165108cec5fae9144af775b9d5d4fd126769f16651eb5fb9e25c3b46ea6c2d250ea59d1c0765b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5417d37f55204746521ce1c4b6096f85a9ec6de0a688be60ef2f18342e3604a30f1b2be1d9e0107c578370e360cc4a8a854624c13dd566026f411a71d1defb1ce2d0440f826cec94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h430b974d93a4ec1540a8f272a6dfb2dce124edec944bf7c3e76aa27470c97e973e6a4d49ca069165e9c95057fc7f4417cede1714317b17c565828ab945126758b141155165405251;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ce35881b907e2c8cc2a4c4aa28015689257621547020cab8521e90664e590c89fe2423143ef4b75daf76606987673b7b8d2424ff6052f34cc9e19050e19f8c9f1d584897d66bd2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ea85e910f7638a957a51814e37aa9ada12e7c180105d97626db680bbcae28498772b55240787c35fb947167e02f1fb4de16ae60e601c68361f7746a856555447e8f0336e0387bbf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h730c835a1c50228ad04f43b12dcfe1a4c488ba6854666bfa3dfb7c51e7f778f3a052d330d4fbc02983fb819b2f86232931450855cc84215ef144e618e61f47dbd894908647fa4225;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb29c4f5728b49d498764fd45305af6061d97e5845ca356225a4b6f03a1a4110b2b27ec9f93c0eb181a06e2343d2f192c27d5cb0cec9aeb46156594213dd14be5f78799af646b47d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54c43984e6fb7e12810c7b0d342ffe96cd5e1798c63b03518cf7cabcd2f07fe9cc740e47b2b918cfe1e7414745b8b7c108f89bcbc34fecdb7b8ce8b4009e4da4f48d6b6a7a1d236e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5eb1f4fd96e979779ded73c711b21cde4b20bbc6b0b5e2e1c4b09a42f4a27a160bcd42f521a8905835b0b4be2847e6845dbc5463d1b209d908d67a60eb4ac4bebeb63f08cf7de31f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f358c7ee7245d28eb9937ccd23ac44899611575f539da5f65bd36c37fda3144c770f402a1ea65a8574880fa5db329b762dfab8a7e74a5567ef316a2c9f83b411b4864443bb033b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f5ffaa60ba71c43e88db20e0ef7fb3e1bd0a1703f716e5d51313d263019269742e180af72b1a3b2aab1161d10e8dbdb34af0bd03f70ee53da3629a2067c546a687a6ba05497e6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed86eac9df24d9694aa45593e0eb70f21e22361ef6707573f23eb77c23a4c2ca2bb3c790dbb121bffb08443c3b9184dfd1860b8c27c6a6f7569e2fb22f40a16a1a2e45333f7df029;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44b774258a7dc693bea4e0c42559f8cfb400d6a9bf215c3ed2f8cec0dc60e46a89801910b64d5db11677c83f1ee26fd080ebe8915503cb27356f504f1425cda179cc9594084989c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he50824328c215ea7e4d0fe40474d7dd1522bc2bda2188d56e6f76317ab1360733888733914287da413c56c03024dc0562d685124f1df9de9734085145ec670bc3f5eff1b2fd7eb52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27fe7d7704a4c17f7a37d8241a51be36d885ee097270b4cb276e3e99749cf43e1f02ebd608efb594fcee1149553cd747440b5ead13051d496c5ad798989454c69050297202344c86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf62886064877b8f5b155395db8d82f9fc3967e228358a8dba8c1ccfbf9a237329dbfcab06672b3659ca3f350aaf1b37bf00a5c080687cdd42e33771512ff5f0dce083c07cb8e122f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h841db60f37b6ef5859ed8964f768ea1794d52c58deefa9877c67e227c46616a0ea18df79e198c9cd1b03e7ff6dab7301b8f000a5f4a4e369c71a2923d058a10c5cbae92265a228f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h277387400a38ea9460abb8cdc97f2a546abd4618059878be0cc22badf4c5c576d417e463355d4edc8b2ee1d6a0038c3be3e8943dfbefd05d63625efeff87eacd07c2e064d0176411;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4be9b5c5fae77dace4511cfab45474aba7e0a104a59e0254a9f5d95023ee2795ca65c608d861083ec53a57b284eea57c209a712d6b6b01faaa8829ed1d0397691efaa865eb23f3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd472e74fa2279f4498c005974c48c350371d7e59f0d59ee28a41344a04fa9b7ccdebc39ae3ae2bfa9dbca65308b5a2d4e7b4b165a8ee1f2b567382e0e2ca98224035177dc79f730d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf241a70b5cdbcc1296cfaa0729fc03a0a97c9cb6c47ee00c05e16d8f2814f82a7b2fc9e066214d19ec4d3ae56c5a71c0c810bcf34c5cf439dc11c5465fb6c6843d6abaeee25326c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa9d367591ad29a08574f7be3677774f63d919e2487c50bc6da4ad9ecdeab55f6120a326d7fab74a74ea8e8185ee05c5881c78a7e80e9b9c6c0fd27a91b1679181c5222921658cc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff13378c3620fecf3ee63c3fc53e9d1030c00b9ee152e19b5b0ce10959fe6f96d8ff29ca6b989a59d04af68d64e44d30cf7800f227c079a44d98b86060aa0f29029e02620bfa2269;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h269e99d5be9e82edff58e9215f959a7f96e19d56b3c7c6fcee227971fbe0ec57b6e97d162811e2a912634df8789e17dcdd9c74f798e7439ccb797f95f97984099e285555d521399f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1eb1a50e2580d80176eb080d4ca7ae453437d3fffb7cfcd53655f3c5f52fc5fca00daca74d943c262c902a766775b34b94bc06d1a0b81cd483f5f72a8316d15bab5b25137862c2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56a4a4f80fa6a8ec58db176e4dd64344a3e80bbc40623d860e4bc1014c4f7873ac5fa228e4d8644260756674dece1bbcbc196c6058fca233c1db97ffcd38c6ace9709981feee70db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h259d968a6511638da6502bec1a85c36af606f74767364ef7964cf481a7b52c7a5f618e08c0e1c421df98c9699d1022902839dfe2c3b681d24d1fabef9695f878f4f052f7e7268872;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6cc219a74078a9f8117a27a0ed84145bcd14bc015240d97e89ef006e41dac07019d9ee45b600bdb4031078b35ed8fe5797c37e1a32528a6c0fcfc006008b12ce37b8281a5591ffe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd005992f2a3fe7b901722c26a2557342d13fb8017ac2f2beca250e5449d672ba41d417ee95cc3a5edb2196403b02a0a4521fd051aec7d5473b7206f8be44ea0c8f2e3c6449e45f33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98c80a77c18442ab544dc39f45784df46e2ca7d56786095669c1f45d40d16261adae449d615029e1548cd8986342374bb8cb5777d1a0c4f70f445442bf546c41c62e97e96df518a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef4132f33b18155ec99e2b346f39abf502b7b8a03f48273736d60f25a0628764f0b7af21f15f21d9ba630d163e21f82824919dd1347e2c6ff41ba7db544fbd89e987e85bb6f2911d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha78b6bd88b125b887cfb98a67c2a09a805652e0a5d8ff442c5674c06c5cf4a3d96c7df183414cf126d00965d790e31e1da013e5f251d1b2ba9b83e92d47dced5f272271aac4296e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1feea062c9d02727cfbb0bbfa3ec6eea450600f9869b77ac4d4681be0c575228a862b52b355d17f6b9abcb026c8cbad8d1bc0e0731e4359e6c6324123da1c451c4d1b056e7dfa70f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c8d644763d4d7db60338dd39f0869dc37f11176d24f11e8f925f9c209738bba10685efefb0920389d641511c38e0d5491f6bacb5bdda3148b9859c6cda08d464b7964e89687a97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66296d27b53498cd80a90a8ec4d01f720c3da2dc008eec6e59cce16df37681490b1ac777d00cbd64564b81e1aaff30c7493db1313255bee49caa76402dcdf40767aaba24024b8bce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbce44c278ea00a91e57fa89c5139bec820ce0205519e0c60d9fb973de986ea0b44fe0a14f221cdb67909f819d19408cf8e6f3a39046202b912a7abf992b0766099e02d122ba7847b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1533bfbbbdfe0581362b07bbedaf84d04e0faf12177541b12e6d7a58376d8f7c3460eaafc3a29e924d641b570eb585dac17d53cbdbc59ce7fa46d570ace14ea02e8d33f295db82b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa8223ba4b42c5c3809d45be6628b2ab52c9a200a10a313a758770d7fdc1d3b9544edb4e1ec6f9a20389f49a3a5887c9521956fcd6af15a261b87782e08afd3f480a5655970589b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h219a1de270aa013b916aa275bd4b5348272020c793b703fea18baaf452b28d789250a3bd82598cbb0c4196ee60622273303234c9d89444754ea21a0900ba49e945568155b66f0a36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3403dcb19092976d33233b3fe6cdad493af85bf4c1b8978881549b0739597657f36fe5b65b12919ac6963ec46dd43adb8654fd1674026e608698e1a088f2d76298c8eedf38aafa4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h128c82ec0da9f8f3bd553945acd5d255468b55c87045d7b1a1bf27ff4a9196f52448e0ea3ca8ae2dcc1827d10e9026450014875a71153a9b8779ea1a0a673d32397942576706d346;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24734276ca358016d737896b1b5d594f49ed19a7cc79adcab7f23384d6a5e46c1486b178c482f6a39513f28fddde7742bce693d954cf0107fd031c8e120fa459f6580b6386eaa9bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fc88e8b46b97e9907102116696420bd95de92913fe5fa33083c93138b9c486260d3ce15741361930a56161f13743ee57154a560532fe044b1fb6a3769390d76eabad9fc29a46094;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fc47367e6addeeff22f2015e3cd2e890105df0b8e463d52c1596ee158bea248255c6aef73211d4ce93525c42b6f33e493de3f5f9588c581055d0734b36fa79f1c1a4b2ee9f330a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed391ba9b607a3dbe64a5f23b5b9e2f82f709c4d722ae35dd568546835831de2e5e66f2e6162df495c0135855338634be0e23ccbd11d2463d942e617f31e29c7c43a8f503813d5c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51bbc4e26488771d4215d38bac927c7212d15634fda1bd188a743a00d4e85cd420eb7199641f715cf7a0f33bc53c2887a517dc0c4d62229899005474af9ba68446df2c99c2cafaaa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74c7c6a43c4f2731e936940810bf98e36a192563ad0d7a21a704c6a7c0910097a57ae469571ff5f3d0946148ecfe69ca585341ded96ed0d2c59ce8f980808b2285302e3470ef6c2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefa0cfed55d58b8557529f5756e709e53bbd3ca8c70bb7fe40191338528947fe30cbae8888d02483a5fb32c330ba13f00bc62a4ef40678a21c59354bf75bbd2524ffcea3d35b5c79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf34c14101c429c1d4f774cba3be6b821f0e75833d258187ba3d3f2d3a2d1734740cb9feb87168ac3a8946ddc8397f7b9aab539305cb5b04fec9f0573679e050a28a6c21edc92338a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4004ad01b99d37ad742d0ad593626ea9801eb5a6829df9c06028827e6311c5db62b3a0d3cf3bb3e05855bbffced277ed20c212678b905acbac7b52e8221de8b279bd1e98c8f889e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83d0424283f8efb22a10513e3250784e994f1829596dd385e3b54730909bcaeb4c4aaeec97b3177fd9cdc82f71d9c2af7bc128e11d738715f5e2c55dd84e51374cfea13921079838;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cd5a85f0a5c2c2cc5cd89ff67912848051edcdda6613ae090a5550e1abf6a728f850cc7e96ec92961b0f4d55ecc196d6fdd8b4475c4f74931591da3023e2a4a10e8dc84ac0cc30d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fee3d907e3a73c1278b977276b5222f7353b6345592e4bf3e8969a2c1d9953ddcc0305cea3c791356df2e882ee7981f9856cafbacb35e8defc117c979c87a7b1039e0feabcf4cc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h767672d0688c50549295f014f4ea3a7b5c5faa0d94fb6fa5e2e3f3ecf7d6ca0814295ecd1cdf884e12dda26109c069781f88a8200dab9ecae3716fdbede13ff06c01aaeb3af155f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e40a175c857fca5f67f6ebe17aa760a3c5a6f00a2c1e0712f0d42b247fa1d996313e6dc2758d845e47fe39fde3c8b80db3c4d2f60dedaa2267a3b02e9e7ecd2a2a89e950211cf3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e66c4d82374b794411a99fbe71111f4df14d5d20235b3abe4b33230266eb794a8da3fbfebba63d9ef7c99612a001c998bd2ee1eb3b0421950f6cd3a39aa55a62891dfe95df4ca0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cd9585460a392c04bb0bf673f479ba0bc8f1d70faa4ab9c2f309c98bf9a5829fcdb442d8febde87722b1f02db42cb0672340d3d3f623711210a8f5b016d3cac8e2e50104c356bb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cb7ac0a7ae9353697e3eae48718646ec0afbc18b41583f3c54ae3d24bdb8658d34eee3b3fdbcc4a84e7bee419ec04aa82850d968e4a8c47a28a9880fba91823b00cf36e810e86ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62c058afb50e37d4b6f224743ff0a4d8c2d76ad4a3e9052a5183b3352e4d842db4108f0354c966d90fbbc6c4841720fd0fdae5b98e7ed0ee121212f16e4b35d482f8e393f159ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98c88801b0e5e5d5d268afd61cd9a4931cb02edad247252f7668366a415c25d0a9ee537f57e90efa9500a74072096270db29ceb4e100924eab2f970d64a3661d9620510bdfdf0819;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h142b1dc0d8ac61693082a0005decb2fc531f3ed2aa5e7c5736ac3f7b51ed4414cb7ee47482864b1a0fbc676b5710824c02ce1917fffb37e9b695b714e553ef11fc5feceba1db3174;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1558272a460b005bcb9c9b3defd033226505c29e613bef89681bd04e5cc8f1cebc2c353370e98643b7bba0fb663a2c24a9dff3a54ea7e08c360c7ebee76fdd7897cf2207f2587d68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he758c7aa9bd436c01c15a8cad186b8f99cd23bdf648fad316a85341c45e423440828858d1efd37f9c7b260a254931860cd724ec93b1f8ba54fa2552458b2aeb6eaa5f9360af8474;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5d7f9c2dada9c2c605359c323b07426c0a14e18fe34b760701aad929e2180b540de4178e2ed01946d6ca8b97424d1f986eb7d521747fddb67b96fc95243abdd8fd6558429bb51e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7323c4a08ce84965129cd8d1c6c7237f04d4324c8c8f71f81b80815f3aa4c3c00d313ec62a4aab28123fffb51556ee694d2acc11cd6736d9ff89fd12817bf7ad740d25d02c798be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67841ffccdb601801a490c2bda766eaf2fabd6e3d4f9e38afe119e8cf030ff1f433ae30479889688758e068581db79037610d55638832cdf01e73743be70f795658e7c38b92a1c66;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf384efcbff6d6065c74b90febb752eb969baeb1e3705da3d63c58581661d9e4d2c47c863394782dc6d26ed1de94684bbfce1ef0fee3a43a196579f084ce8c180d492fd0207833c47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc574f6ec64ac1ad04387d87e0680958be0e4128b5d5726ddfb3c400082c236ff34ac570999ddf029c90a5de3fdcb2d9144068dd3291ae392b9a2892aee134693e96efdce8f8b8902;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ef0440279a5332de859f24fa4d3b199a762dbb248d3ce0ca16834d5293b3f47dc6ce9de37393bdb71bd3516242f267bc9cc8826467b59cb6680cf9380a6f347c2184e9bad2ede2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h341e345001ad2ea3566b00a1a43ff7c5bf1e8dd29107873218e06b05627cf81028307631546e9f53915137ae4b971e925d0838dd08fd694a81618899a27955acbdd83a48d69a23ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb0a3ee16a6fdb420f451b759e7dfc3d842ac79b06bd46f1a4e6cd08afa3e2f101f8af857b67f0d859520ea98ad3a8ec5ff307feb7ef65a6f44d9476466a5fbf85ce336f6d709b33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h942a9786974d087fe4d174b9158a43b8b79aa31a89fd605af402f88b9062a8aee9e66cdbb6f23d5eb16d171261e20dcdc02f76ed82c017b1632bd064e884dbaea42d6077eefd7c1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h371f79352c470f34e95edc53289ad5bc02d258d435baefcb88fafb045c419f9d986cfbe6927a9ae6f60fac70493e257c0e1986d57429459b90d415d03fc8811c0a8b8240f46683d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8f1de6a5d5242b1eff40d9f13e89c70f28b2e4eb59577c49257dc852104926687881dda56b9bf606bbb124610932234f1afc5cf3e234b2e2935cad32ee4d78a9c35778048ce7b12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2297fb30ebcdc5c7e4903cc220699761cc9cc39511dd5b1632026cbfdcffac7a4170887308c88c9cabd3be16ab6d530625ab091980c55919b8c771c963986e05d2c0f813e4cb2028;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc59e282d5184fadd017b51bbfe3260e9e03ef09afce066ae92bac7333d52a86e97b800c44a6e7ba269025db9b850ca3716fd000d9d9ea7ebb6cab1f4829989f404b9792346fd2c2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bddf058f413df80be14cce89bf98859d73ac60ce261caccf4ddfbbd4f31483a25c82e6e73ce421f11ed511338c17e2c0c4c1cc7b7e62699cf516ff8181cdc99bd53029d93348105;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7306d29a8fc7532ea973ea50ae2c00cc647a35ec8dcccca01dcf2464ccb3d1eed355d2ce5695ee1e529b1abec530e8221db6a14cce4f421508a0a0d9930769546acced35ba8fc7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6311f7081d372b17ad6cb4f68925952155b76de3988cef0993c3bab77e8f7a92248e6ccd49c2418c7d078ccb5609bae3e1140f631e3c8bef6d283909cf77fbdf1342c11ee4c5f4a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab0f33f6ec3a91dde90b414b6c434b4925141ba1c28e1c6368c3c1ac7fb7cf78a9bc6a43af01be58e1aaa1881803f02fd38ff2e7ce42af4b2ec82752a7f2bd09da8313edf4f589b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe5b94d8f9ff54ec5d610a9d63a51057c58386effd6ff8620a424edd4a2193085ba8f6dde9abdf7e57ed0537f2c2dc948d76d19dadbae00f49891f56d8f51a835dca5a39021ee0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13f0a2ef7d0a952c4690ef0e8851590aa8501232df4f601d83b01110480a574097ac85c396fd0b434cec52ff68a58572118d1dac1144a967444ee7cf801e0dd8e57789b5b4d9ae5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha27388e172a6b31c546bf4d7a4c8940c9d1c3e79b8227032c81e89371c31ac54e4adb771e5c314a1819214a7ed93c1c6bf8d58caff3d46efebe008a39eee30e56186ecb7bdbce34f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae70f1d088c4bcb4155e6a932e6921b57cb99fc8cf5794d77a17df9e9c2e59ebcdb1dc3df169f862671bafeadeb7e589e1416236d416bd8aa5ad6900be329a7efff17336c4c561cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43c9b68afdaa8f0fda4d67c8925490635d30e67bf3f156991a11ca8bc5296a1b9651f4590259876419155a3ebe9593a26424c84ace026fa505f465e1e32e0479c33145ed476f9036;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haffaf8ec59ff1bf0f7e5d71375380030a40e7ecc5f6c4e1822492f47c45b50f2028332ea68af4c2c892252ec299bcb6ece17a7e35e0b0c443742b1d85f89301243b060fb8990d6ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f0d706359f64091f42969a69838cb474bcaea7d19ce5cc30f59cc3bbf985077f19311e33aa5b73d4dfc979aae5ec0abb60304f9bd0ff8b247761b2b044e7faab0a590ce835f5cd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha72dc25320a7a0ce8424fe3bc66b80ab932d09168fa29bf9fb40687bccdb933f8496d75431bc9ca902f89a9970a30188d089f6caa79a1180bdc2704ab1818e54c70dcf3d793604c4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he941b289ac1bdb54d199abbe8f5246362de3f0b2f53d076e16d364ba4513ecdaa6a0bba081d098c01f0dbc4d3d23434a149efcc04dd80eb9b56bd72dfccca7d90028844d4b9626ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee0f6d44298fa3c16cba1e87c87f6aa47062469317cdc707b71b41b6941443a0bccc40fff32dd278e7206d6c084bf07751b689a3713fabed959442d039b92770b96652dcef7b6943;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a23cd92106d353fec5c18ce037831d86a1048c2a28e511ecbbcc5f3dc44fe41fe69fff984fb53855ca79b985d07fcc1a5635f708575abdf43a24e761156f9c4d4bae8ee39dd3237;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ff76c602f2eb13d5d66622372fef2dd1be59cae84af9080d80e33038720d61fb8a471c36f38a10006090ca9c084d84e14a840f174599a8aefc9872ad805a17e9f62a2f244b65ec8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h496cced46ea17a672c0771358222ea1a820d279bdf0d93915aa8a75bb4a10ee90d6cc1ef7506719c2fdc0c0c867a7d4f24b5809409af9a5fc25e2e093686f7323c8172f4c370ce8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79b7f902cce0605b55c120e38b8df6fe894b62742c3b54119280bf40a610b065c84960c402e276dfba3796a468b0228ee0c1df4f0a24f1ca7622eb3d5ecf3f1a2416f4d66443950a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd101de32bbdf03e0fea6ac90af2d817506b656c57eb83424acec34334ff6ba9aa5e6557bce34cd0557b67f12e72b67be927258fa9fc9dda99046522177aff1f0ae0577b408c7830c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e4ed1337811a7c5633707e48e29902c6c43da31362620bc4c68eca65c52d17c2fe198f2d1c60e328ca34630fb69ddbe0ac76da60b81645c74acf73020949b58d03db74c9eaedf7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2cf87552d2169b07ef246c6e9581837dd2f474e1074ba1e2713ba5847db7be99e77d3f64357ca5a4434d18ee2de27b63931ffe724bfae05ee98eb5e323aa7b1c2e09bf10741738c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d7d16347a523786ff20563558e19dbd9e7c189ed357de27197070e57a50a297271d357590d7750971c58964927dac622d3ea4f6417b57133c91d7c44939e12fa09172b503e804e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50c402385c24a1bab45cc848d7e84adc18e70c853876ca3be7e4f450b4504ab8382db0a8a561d70252074a907af43f7e423c22d8adfa37d994ee4da4ebd452bf87f2ff888bd93ea1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h902cf65df9a3e7a2e925c5ed989f828850f9195691e35181cf44633d132ae46a88a34379dc3b937516e4a4f64e6335e1997603d236335b371512260a7aabfa7bcc719d8ecddc7c1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49900cd1a0d341d3b753c52ac32cd822d3b65213523f95fb7fff252798ec975816fcc4d69a5616b3d1e570954b398eff022a2c419541a797067e10b9d346445d319af4e7bbd36208;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d53cd8665222b1f896ce5e05b53097c2f91c5bc575ce99957b607703e842b01dadd8bdbf11bc30786ed3365f6fd789a28832f5c72e7e8f9de404fd4bc03d73dba3ac324d7318e85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8de8a79d3ceea785fbdcafb23a3449e50cc98d76ffd0b6eb1fd97cf7d7bff2612df93969753c84ac6436ecbccc0e91fe05a5ca00a8c7dadc610908888c6b253d8b51217e6e9f165;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48f0936026aac90674de7a7c88da51125301482f9fe5ed9683cc4db62708df58edd4a1f25f670aa9d7ad8273046869a708e2ade482775a988494b385f667be53104133721a875450;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce68389d8883c0996f396bf5afd30668baa4220c79685c9633f2c2fd8e2d3ac44478a359495120458748ec7b8cfd04ea207b258a389936e02555fcccfe24969505e4680943e503be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd51174bcd8a4fbdf0f180d0b7a19399b048d66c24e0e947095737319d76885367047fafcfd68aeb79c8df709eb7737756cd6780ff1af2c8e5526961573dd2501fc0bc14b8a02d041;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e99804ae26d2a42fce8bc5997670b382a681841974c4b0411c35206e4ea00c0c182042b6856b2d467eb4b11a765d6c301215c4962ec9ac5c7a496b2eb587c2b01b47efb7c671293;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b41de607e8cd391a9c696067411e9f72325e4142a4737eb36b0cf3fe8329d81ebe2419bda66e429cdde49a154650d261c50f83fa3e3ac314624dbe505edd67b89d9fac462356571;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28038845d7469dace2e2020b56c98f3c2e24f5f34cc8ecea9dcdf9f8be9fd040a20ee41c821cab88710fd6a74ac17d4c0f96f0e49666c91532bc93b4cdeca0cb837c3d5540b56f13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1945f3e780ba5e12026502b8083fe14fbd3f33ec0528bc826de6b445c11b1cca060a109487367de382373945fdd5494dd5db11914b414b6b456ae12b5817be8d6ba4c4f6aea60898;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcaf82379ab1d0317d4a927be77a15c35a0f1e7d32b43e730b3bbfff57c3719b78c68406de74af50f1298b06eb509cba7aba51382d29a64231a4b94be43e95f5fa981d9ee856d05cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd7affcfbacc9fe6648eadb21f478c83b291917352c66ed21cd4f6450ea7199aa5b3af09a7f6a804be1f5252c107568ee4fc941cbfa8b57b32cdde61372bd736472bc087f1227955;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16543a358f667a5997f152a18681b231ef6bd2e293d2196908e781e83344e40c199e547f759ee4e3c0fa7d33ea4dbde9336ef42c9b1ffd423f289e39e4b2fba0db6a293b2fe32bdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83cea80486dff061c2414cebdd731eb72781c5746c8f59f13274debdd8b8e4da695189274678396505454bc5bf2ed6a8e89577e6d54059866b3b377ac19d4e027cde971f8a888ed2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3894919ae4a654ddbd4695ade30a396737882dfaf556767af3962d56c6ac0dfdf5ab6424234f9ee648e5cd2b9679d81871dbce39342fc3db9f3a848058181e08d16417c727aeef2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a89f551ae72b64c239ad795ccc9932ce37ab086b13e5cf776d6b61da23e318b384477282e30431ae5edfabd725ceb581c2f0e95cb26f656d8e89394b08149301b205786513c6b60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdaf417aca7017a129c2abf8b62b4737ec14f04409ea5d63930d1ad4a73f50abc52bae394c4b8bd8241e83071bd3116f51e83696cbfa6cfd43d92cda961c80a5b757f663b53dacf03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h259372f13ceacc5b50c631cc942c5983e6fdba4f5b792d233d0e236a5c966dcc5f80cde5e1a6c95324633cc06fcca0c8fac292ddf3e1e2c8c81130a204fe78d170a5acb3233e33cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1abb27af6cadcdef736e006a6942e98d122970a45afe6a8569128b567812993eb0406225d27f739b98ec81e989a050c1b658f5ee3cb733170cb5b8f7a41bc174eea6d7bec07539ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbbf833e6141b8e2bdd14e299775299c60ec564367b80974dbaff1227b63af948425efb1b34b116dcee0c6327a1fbc9370081cce7e416887961442efa15772741176096fdf361745;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7463c83b27d01f9eadfc0b064cd8e334b32483bb67ef4dcbe2ac223630bd96906bfd00035ba6bb2d3e2002ac17c86d314732de0a4708ebfd5a3980f20a7b939bc0031c49c7de3c33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76b2a50855140b8ada527cc35e6b3bed11af9857120a5d7c99232cbe60b6ea059a19e2e520ec362e68850d385c21733c5df477d3fc021eb40a9a037c935e0f7be12a36f4248fe3bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24f497661f3c3ccc69070049abf540f7daf5ae2d70d3f9971a2839630a0daf007962aac5dbce6353ffc4fea928fac3cf0f55bfae91224cb9b1539685cd1d323aacf4c1822cde68e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f45a438810eddf9e054a54ef77ffd5f1d89e300e4230a2d2fc8228d7e1a5e52159af456a4f89adc0c7327b05a5044b0017489359cd514bef2221da56ed3b176f3ef73d1a64c74cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e89646cb18e18f2ba983b9c8bbbc7549e7e2cf8cdb43a6aedbaa4f43768cc660f65a738d897c67e2afdd9d9a88cab9dc2d59ae2e188ac10efbcd534ee60edc902720710eda997b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ddac3c5417d879be79486bcc3e1c2b5eeffee96b7a73eac197043f5370c2ed08e460fda0508c51bc01a7247f9234016b98ff066254fe2d2730c3a8e35e184b3888f7faf6c2cb54d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73785fd84816e436d849e73776d63fa0c1a07bc3279d977dd8d9f2f406df81bc84ee91cb56e2560a668178ef6626c32f9abb62483a20dfe23d7f619b1d21fbb0d684f09ebe61532b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a3a7a0fce9247ce15a3245bb2bc41ed6cdad6f71d72419bf3f09877afcb3ab457dde9c2ec97c662cd61dedd2f37b13381fbc032b6916797d09c7215344fbc823b7c5608386d69cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56e551781d90fdfccf9fc9d8a842da3987af19208e3eefddc4bb1afe5e4c57f6a31a7c10fc960899a22c8c1294160aed32bedccc419160b04d805ba7f79ab7a5d5919dc6e8197c7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d1c8e61092e7f2db3d7c3915ca7f58b99d6c25c0c49f4303e603fd9be52b7ed941d846c7eaa4c08ce7118088d70f08c53fbc0a9b076a3e11388ac3d47cf989a1a09d014abd333e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd17ac42a9d3679f3cfc33a30c43997674b323c3a44cb54f7e898383912eeaf220d06867796decf6a2cc6444c3c3230b46a3243d571059ee2071b5524c06adbcd47aafdd143c2403;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbd4518a2c4001f9a2534a527f4cc0c41a293466488252bd2e17b7b52c96dd2de5a0ecd8ac9a16d9d2b080ee317b01da541dbcd782cf6cbe6184271aa35c8c06df6c396d10e3d0dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefea46935144cf916a59ec5dfaacbc88ec886b849ef19d1b792bd4939f614a18e44853f1cbd225b75c2ad62a624096cecfe0587f6e8d324197298acdcc382e4dd65fb747ff77e442;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddf60147cf422fa0c1f04e7d60ec172394f50ae2f11848b6c8ad1e0967f7264aca65b3a3a6cc728b2c0a688f9b315a8054e9304a364af9bca153cb1e7851b91bbfa7323c969fd0b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc63a2596764b96ff3f3ea48f3e909cdeee18fd1c61a13d3325d5e825fce56dd0008cc5831a9b8b9b2d0e26a488b637a1db7b9bc4bd9ef4858030725fa249906bd092f64670ed9d79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e5cd28dbbf2cea6c0ee056f044ef7f1faf69ec9c9949dc6cacbf922324b98588cc028f1c82b1f2152c939336ad457bbea4e60f58c9669f12db66c99561a29fac542c2e6f1423a5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9297e91f2cd2c571625ed43214d6be552920c93848cd930a4ae990bea020b69124514586824090be58b1688954a7c73019576a91beb148d5194c294bce7b6d60254a84bab91e0f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7ae5b770b3f2bd546ad7934619fc94b1d3628075d033352e4bfeec5d090dfe4cd9c39b579b2019a9a3cac1ff5ae628a5790412d8984ac32c755972505987df9b76bf4a705eb0293;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82110341401d373bc714a20e14c1a31ffc1cf3fdb12a131296443449810dd5322bcd91169ea275b6a130d2cb46028e9ec431bd340de79e3e2af663e296c87941cf3d407eaab602eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5b42c913693c1cf46763fcf203aec7f8b3f0e484b4c3f349767c733a58b563e8c9a73e7186603a24e7b96209df1a51469eb1e6351af3d3c41c4d87638ca998d2673236be5e746d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cb53ff6a3b966e2fe425d08afe784c5d1787a75828fadcc1c28b49b656821e9f4863c495b42f2bfbe951f6452e482b5d694f463976938666fe2461b6c23ad1260b618dd23cc8007;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab1ac0d605dbd85989b4b03b46671134420ad73ee3a17106e1e15a0aa15ad5dcfe77fb4fb4670d4b0dfb6e24a20dc4e9c9ec6efa2622f13047723519e2a24bbddf220f6789f2c8d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdb216027f82c060d8ecf6b1f0237cd3129ec4a84db01ed3a89d9bf6754c962ce6fa7ae0669f1cac1305c552259f04145a0a352dd76faad715d5c912c951aa32b6cc93bacf831099;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hece67181ca966b4091402a2aac4ec18ea07623325f35b518d678e661867759db3fd5bcc858982b442933a693a9c6a59bb92c84c624a2fcc15bf9c0a0434db9c470834b8dae6136c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbf54525741ebff218922c156058acc3eaa6b34d3efab147710f7ea79b25c084c1b62216a9baf3c6294eb2ebcb444bcb3fcb1c23605cedb43e0a4e8ba14c84379ff6275dffde5746;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d64502fc1d02a1a93c130aedbb85283f5b32e097d6451333b2fb04176b2383e393843636f5d6bff688e9adcf0af2669c1e9cb1cdba4f788f571b435992e0bc729e318312b554951;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2336bd70b42ecc26e705be9d91d212377c0218387da6115b13d6000202f4513fac7c62e3e4458e3a9249a6e51fc88e2680afa450ad4ba0284a0c8c56c1801898c5199296ec759833;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb938f7880d63380107d78673cbb0fba1273ac19bd7be228878af439b85a1c2adc9c2532f95f883f6cca936ad98ba0f9db71b7168ecfd596ede737c2c12533683d40b06a07acc4660;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ca3e1dfaa8aea48759e301334bba01fed603b5f26a88841bdcae1c1bfb1fa2d61dc4923d1a15dbd54ff7f9b300521e88587ee7e1b3a8257dc1cebecab5c7599f00240477dae9e28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4398befd373c23f85b9140b0593b1e7fe9c85462acf6ddc5385d3088d6c2030c7effea041ccc1fcd2973638fc8db5f545033e7c28cc4e730874628b24d970e402f2a34c067eb422b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f0ee30ad0f482007c062bc92fda27261c7d47768c4b55cd34a81428a172d83afb18dd8ba043d4099ee876a182e8dcce23c5456a94c9ae51de0b7b4e1db1412e8532d38621962f41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf36a31838e5d9c4740f2e1d67b9b1cec303754c891b52c92d07f6d2c4a1e20e5221c271a64bb5caeb66e05d816f883380a76f487370d4e3919a804060c8cf4bdefd83ac326eb5633;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h996cef714769458682a42b2851d707c33970df94a30b6528fa83c1a05f8656143928d3c445ab76bab72a1bfc0fcfde3523034d74caf889df1b15b6fe8f5fa8345a8f9bd45e64892d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbdfa2f3dbdd14303c515012a3d07df65110b2fd0d94023868019e63be57d2931fa7e0547b0f80df3dde348731925e80df6e74cd3391961ee2108963906dd71dbfc9198f87a0957f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4c1f3554b880c3d3f5f4e320b7c9257c22b80fbb90741a74acd26d427433fea66f0d421c673e65308f83e7042264f97b3af556d9cdf78f79bbafab7a47769187577414b9719959;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a695c778aee3a786ca1729b7d6eeb8268a73fce78cd67bbbf917d5d06e7694b0677a5ceec99e31dae103fede36dd3e2f9c3a49f3d96fb99b8f22dde2e30b64a30d19e5051bb0d7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he70b446f9611b00769b9c2db3cd734a0277e4daa4df2a29f4fcd08fbec2db649a9f067ce01c39b7c7bd523a1840ab1435b4f6e9a8d481218197454444c2da8e710a86fd7fcee5316;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h641cc5b1a39a177d421a0b3e477c292b7e2b5e198a0c7f69f2ddc6684da52c8a19c942cb79499e1a360c45e35e40b47f9f06156a60e958a1400df9864bce27dd1d3b94720785f2f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce5f4d124e15f92926fe2b759f47ca5aebc5958c3fee1ffd80c718854ce45d8886367d5525ccaba655b5054a08e4a59d8ccc5bc37c3fa03ab96b2ab2dd7eeb6d12960fb09242fa51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29e53bd11a43538bffb492957d5a8d54da22df68ab3678118f5142436deb52330b46e279b5d5313024bbab7d3a26013b858e38ba0eb17da09c1e85b70f1f2097d4963340f8e82c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c0e0aa761b49d8fc41c7947ab2c0af34eb2d1043e3489d6487f03c5c56692bdff5e5748a29899de87ad1887b95b55a46d1d097394f2ffa91651efa4e0d1e51e1425edc2ed4f504c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d8ba9d90892dd6a784f4a27fad70977de188634428b38d838e7845d4d750ab09e799101194669c31b376348cf80591df04b2b30d430d13069a32e75ed138c073c353394b9ba906;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5101393873ba6861c9001feecbfa953b0b4ac4d45988a1e73a2da7fd886d77b30fe06878ab4dc73ffe2ec8e50bea45f1ab9204c2372f52129dc125d9481c51ec1808269b201d994e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h750430c03fd238762bea217e34578453b87691f3b4e4071e06fb38f3487cf40b63dee48bea5f0092cfd36767d15ecd0887526b8bd6cb98519348742784ebd8a1bad4cb642ecd1751;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75114bab4798ca19bcf4cb4255907f403ad16d6b1d89a060682653dd40152cdc5ed781229c50766066d1018378149d13efa7d7d19dbbf7f65996c6d3828e1e75c9f937898ea185aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4579a4b62c57fff3c2cb373102106ea05a3ef26e4944f3391ae240effd65b58894daa3cb215688c695bf4451f7ecd8383f9718d4ea979b765828407785ab22d376cca9d22efaba36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dec9b12cdffd901752fecd846eeb39a02f4484b74ea8c284841da3cc1ebd4a2c3ceefe8b9b4d896343e6d1b38ac8cccb2ad6ec76c1b12d0381fbbb0aeb3c8ddedc0a1f6fad7e11d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d80023001777ecdfbea1a5c85447c10b703c38e1fb7e0ae17ef1f834996e569bbb968db74dc021b7ca64df41b7ac3db164af8301f420fc666f83f41cbf7746c47f73666258a59c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16c256f6bb94dacd3710cc13b27870990d765a23a95061ee3f5726a30bc6115f2a847ecaa1f45bc8e676bfe88fee6e356e86f4499eea3d7ffb64281b88763b49b938efeac0195693;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h617f1c77e1c414a4a27e689e88f9ccc94212b3b8e7fa1e66b553965927106e3adca23cf2e03f1c989a106232de0c7f2807933f42f437546ce663c1f766b308f49e7562a36d48a5b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8346d57930c4abfc3399c2cc0db28218081c0f0d349037fdd630f01b9ee9ace8f440dc010a49b83ac1ec17a2ed3350a7b2f839e1cd2de92c7cdf37b981eabeecebc82324fbee311b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88a6dca17151fd21662b06dc841f53e2b2284fc10ca26a37f051e1a475f3da0e25bc4aa3ea90ec4c5d0ad46b240313e047b8cbe4a4b425f7f4b009fb9acd1f62500f0a281114a7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdabed1247fcc8bee53833af5fdcca388d9381310c7d1341d8b6a1ac6992155bdbfb1bf157bf938064e516b061305f57fdfd9130451733f3f2af2c964108746306cae08b1e0c0b0d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a2a35fb031f7b60ec8aaa2a466a3b453d21709193cd4f45f0618e4b3cc5206e1bbc174472532be69a1cca0596caeac1ff08d89dc1ef22c30ab5a46570395c8fd9e85a191a0b22ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha815cb5882a1a172b32549bee97d9c2d15d97bae3036df72a20457680d9bf29a13f40829122aa5997318a2f7c495f43894eff7e55cc4745f5707c4aecb4e89381ec447c8704340d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52d0e589689a8f44a67ff17298b274a23ff3cd535da89424212b534f0f26326d85004e1bda2c81ef24705b1be9cb0fd3c87422a32beb1ac8b4ae1e358a21d778d689baa170577407;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dd123f24e835259e865812c67a39ac1df8ca71a0d62f3ea1fda5948a66c79cb00aeed0a1da482cd276d6645a36816e62b6864d14aa20bb00952fcfed79e8ff0a6e9a78a039864a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f1d1f02f13629efadbe2a28014fec916d486ec0d85941d8396a32aa0d533d788cd3a00e5a06ba3eb98d2ade15564e28b5965076088da2bf3893228c8ec1f323bb4acf7684e4ba73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h287a7668ce478b6f7e9dbb07cf27cf809f17f2ed8f68f033d9bc556a968dd85ccde14cba0f352f9d3eb2689b4855f8ad4f725588a07d5cf4a93024cd53565c9abac84e1bab4808c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f9d461b5813fd2b8d99713d2b1c07426aeb314329fb79ee4e61757173b32ef6f45ad96fbdd28d824f1b9e0d1f32df7976c36f9b87881a572c131d837909a4a6d002faf7ee34a39d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3cb0aa7473d09360c619b6cb0e44afda191ef63df8193f5a60ba8d2805a7b137e7a1627c390d9ce5d99097eb50c4971e92b49a7be184b91f5be1fbd54297d4d3c8e1f55994062e2b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1016a424fd87bd4f6e27a2e2bc4238f2e43f925e8d5d3a8b9695380d87c63ec23fe70df488ca7f482c775c395c8791704a20a8b31682ff55332ba49beca9a1bf96e137e6fe1c5eee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2815bc1f45d3d2f3558acaea02db8a953a54916579ae7a01ed9581cbcd6264f28ac75771ae5f6bdeadacd52260ad45b6972cbb1c80a7123c976be97c82c03188a54dab43db0710d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h741d92b8cc76e349a1953a221667e621158fa677a9d2fc769dd7f4dcce97ba1b1e21e6e957a01de6d5b870b136c0f1b1d8faadeba680f87f938f8a9abdd3d8294d64edc57251b0cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h483a959e53d3983a3f757df70e7da6617810a49b0b73a48198fe7d09684884663b59639d844c7c8a40d876e49b0336a8ec29c46f1b315172b8168f52b4302db7b68d4956c96cf5f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97008fc2771b8ba6e7c31f4c2dc6719b377011d891100f5ea30186324bcc7148c1f871e914d056c9bd5e283ff2270a6fa7a1f71a93bd0ab5985cad68e5b3308fe63418b082234bb5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1de96c95ac52f22b32c33e9aba6e8543a716bbc033bee446c852dfd35da2759e9fd6bb36872a7b5e36ffbe6435751b173adfefab39e196b1d3344a5cc28b35090fcdd768494be08;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43b00c217f3c726dc9567be6898faf4981549973d38fc45d1ff8d1de1a3dee9c80b330a93c907519756d441c07011b33e071b1bdadec1ad0c0764f884e339f3cef58841784b99b06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7e8b991afbd38727e08eb9c3d7cda0552da2fc9c2f4a202611fe63cdf2db13e54f8a10aa684f3d6ecb944be44e64cc41dd16585846cffd9993b7268bcad12064b8bbbf1eac93237;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3f154ae168e3840b4dfa7e3f8d14f5c7c25dc0b0ecebd4499b9139666f796c3a1180f1c4fe8deeb9fb24b997b4d584bc43ccdd50139090d2a56fbaddd8a7cad311f866699f300bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffa9db1888800740c665dc48e9327ca4f0157c59cd28b49023c155fc259562e08d83b32eb887fb9091f092007dca8dd76ffdf68b4ce10bd2f76da0aa2144994c1a3068c20ae555be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc746681dd75a54cc5f01570e2ff261fa95dfd7698088efbe23f2228c27cb8e7c3b82d88f5c80c9ab4bd714dc8cd86fd77b93016c2d2d70362de9a79374ebb4bdbd334e2f199eed4f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b054d21249c248787724cbdcd64bef983a97bf16d429a750fa4b6c6b48181af06513171340586730a5a2779049d520d69400d209e3b879a5b3b9d64a6d8a1013d9bc7e9785f409d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc54855493eea8d9a2b75ba7f84cb287417b9412e59470d98d259efa915a6bd9370fdce44c56097dde446f7064ffbced4dd3833a2db353645e15b26bf9cde201aa2e17ba0c44a8af6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58f62786da1b678b75561f28c2fd201dedc2cca728584db5501fdb062f10eb03f1a2de6dcff645f96e506dfba36c742f129a0e251a85603ef397d0355153637ec5c9fd178ed01bef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecc523a0f8106e070904df8fcef6d6c70c4e6ed86a4192259006871c63cecedb01116e9a5684d57b31a4a697e1639c49153f93bf49ff48e2adf551aeeb3edfdaeb5ed8cf9d07ff97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fb457646a532603dd43000c17e69544bf7f5ad454efe2489a28f350e5c82cc16702451b654b7152cebbbc9ac53b4b4b546d3481f68d79001ac6092ec117cc9b00fb1e2b90d00ffc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35cd5d4dcf35dbdbf96a49819bbc55d1ba88bec818ef22dc120cfd7e298915dfe3a3d72d29fb6c3f8b28bf374f55cdeec97adee85950bd208235c8ef65e282120dc5a7a237c69770;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85328af75f34b6efc035a739fadb2c42a06b721b4cc565a2b0899b2b7124407c65a6ce68c7d56ad0134a0aca7f13c60f004739553b0cb3df9e9656a5b7ed6362b115cecccc2aa28c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h914af37274f0e8fd4ede15dd39a5c38eac7ab49129b5ab288e38d4b49a5b6eef40eb7324dcb1c82477ed1edc8137548969a53c2b581ad00d9085a574743914634b758fb9cbb55a5d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a8b698dad1677a656907f4e048661ec227446969edf8aad3e51b053d7e2b287915fe939ee40f40761353355b7d7de038b7b686c450627e279a8d9b73c1b1233b96e6cc798aa3c5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f963185703c7023a52c9c3191bb94170410619b80248d35eaccf171f67de596eae9ef72037e439aaa1bdb15cc35994b00d4b376c5e9a28bc7ce4cfb0071406bf61fa7a0dd99d270;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8eb7f8e3a5e4d7b6ba01b8fd55675e02349b950e8bced517702e35f6cc0bee7c8f8408a8400271f30ff44ba6cf3cd86e4e3f9872c7e37ad71e4c462f9461593ec1e61af794acc687;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c0295234ac0e5161006c0a156fb1986434f511cede388da0a8410d0bcd101bb684892fc9ccb176270515b30b7f728d078f0d2fa83807bccf17e1b25bf68940edc0a65d303ce7f1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haffae5bf56a6816255414e0258856c35cbaa7a9b7d8bcd08dd8084273da4092ce6afc627d137cfb611ae22a73bbdd639c1acd508766d31807e615b432cd2b5c9d0e43a0a56c79722;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe8455899afac171ee5c00a4deb875e0c68f9f72ca17202e0b0e816f821680a824e75c4e77f4bb0cdf7903d03bab53db50c915c02eb00cf34280c3890d8648bfde2fec72342e7d5d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc8cb6eec81ab0233270b95bca0fc5c62c739e593377bd90a56992a9cc8562ef5865439a97b71d4d35e5637e60f637ae3f973fe05815a0e8d950320c21003c715efe06ae6c5a45be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h861525bf8aeaa436b87801c40e8e024a793c2ca5f9f44e6b0cd9204f10f1e4d688479cff0b75f063e14d2feb187e2603103f9b62a85ab438e644fcb0324e535ff07a62a46eec7a02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5762560fcd3b5ed556749b51e330e10ea5f061d19bd32d8782163928d5a028a5117fa6c91d19e73749ff867a141346b6f76f59eb2b027a8341fea3e4ed4c6f792528a71dc3ef73b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2aa302ae437fe0921f8fb2ecf6f52a7e854415012ae865d4d229794f8ae401e806376f4050f72efd34744fa53086bf6de7a549f63ce3deee3fb22c0d3188e72d6a5302f239afb3c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ce210120333990f57a9af4cf1bb3e71e1fabfa799bbf5ae49a1647c67c211285dfad3337ee872b435314b48f68ebbb38490b817f7997dafc10c6499d13b605e4367f908fdab9bae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10dba7f269761cfda8dc5d922a6df6ce93ee93463a2dd7050be80bb9744362bb9db5be05804eeb28b2c5e9ba0934fe55eedb064b737680c096d7ee1d97118228ff97b8021e6461af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha74cd3865f3321315c89c0e2162573b69d503760432163edadd2e46e55a5ab922267f9a7c2d0328a5ea253b113741ef57be19a875de9604bf8832540457ba4655af63eb8c5cee5ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdebf9de484256d736cd57f2f6177b555de610d7d7e5f8e4675897d20e43a40af1dfd5805345178e28bf7951ee357b61e7b0b8dc1d3c487739f7b89450ccef24743d192edf1ea973;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he78946b32515073a61ee02062ac1a6dccec708a0a889a77630403bc750b91ba7e3a5312e1de4383a9c5471385f787a83df12c6dec6e91024813695ac329c619357a0ec7b16c0da66;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3efb8f02b8e32ac05a1418abe40d447012d9d8bb631f61007f7beef68af0221c0f51615b9fcd9db992eceb82c4ac86438c7d09c4f7096df285115fe596de50aa43c1568b49cdeaa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7e2a073bc585ea2fc1cbd92450c8cffa3b213448a1a6c22f22d1c6ac9e2575648116fafdb7e98debad3149f7d54de9a077a42063a2f3b16ba77db522edd8a22c0e784dea9ef55e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h785e64410b4d0c060a79fc7490c4c884a2ee7ee4c744eff8cd7fc867c162773f93e746b4e1f4438f1fd376cb64ef195454077ac00ed6d2408af223fca39e8cca00ba68f0bf8c5e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9da9adb104b10675f37e82f8e27b71687dce5dfd70efd09d5686deb36256f9ab52b5213280e03934f46d89baa00be977d3b86cf1936f097f2399335bd2581e7dcc3270dd0610e44e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dc4b9b1d701f565d67e232da67525de426c99d59ae5a2077a979632f9ef9e6fc97c4f6254fc01c907118c86adf3b929d192565ac6f14141969c21dff18a91fe4fd4ca2bb5f631ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a83aac947f9c5250f134ba8942f2a71c28f2b29c11e5ae987de5e7b37f2824965f11717b11e8bfab27526a6a80b6eeed5f42170f8a67af5031acb0b8002fd321b7509f5a2aeb7ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71769dc258ac434d4f9b86371724d22c5f901d800d40875b45b4c1e584ba0c8248650e303cd9b6e0199040e2ccdc437b74d85782675d71da419012da73a27b54e185459c7702dee9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb01ad7a55caed76beeed48f5793b035423eddbb331aae2809c0bf0c4632e9759d0f254633365784c64e15c41c8c625cff0ed1f757f0f17e9afd7e93a4ded658be985deab46fcea8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4f806c7a4ed875c3110fa074fa1dc9510de9213d00d7c7d499291ec66ee99a39496a6b1123ce74d7dedc9fd834927ef9393c7aa1221d624acc305a5123a7793a4f49f74dc007bbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1908d2f4bed4eb4736cb2573537bf953ea1f1aef3be327da80daf502599bc3463de93e9f6d3d8c2724bce9691fcd3b20941dc1b620e77efdfa802966c380251adae3df5c639f82e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56ecf2ef2eaa87fa9c283e73ade2513a627850e536c0c544fde47fdc27174c9657aa51d3252a71a8eedf8d33d057ff4efc7395ffee3536da6529c0f25fafc3c6066ec1ab46b59793;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22139b76ccf2d37f54f3486f97e8c22edb7b73e8098706e7fc70711ade0d0699b9fe220f8b74d09609a987de7ae60fd0eb31d4083e3fe9e36a587d5bf77ce33d4964d8d2bc22342c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha12500e42a18376082a22a639971d706abedff154730fd3829f4f1e1de4b679eab1536d32f77539a662fe0cf9aa2da2ba28f8990ec046d6ad5102ea12345f0a9021a7400d5870fb0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc6d6fb4a4c83bf21c5cd6f6d3aca43856d69594b7f65afb746ebafef8369a50065b981df9125cb2faecf2a3c7c93e65d50b899b4c722ce7b00147af774977291bf017e5e3952a80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h666539e6c1f4581f45146ff9249c7ff0bad3812cb1841cbb10d6c940ea585b39e81776675dac9447b12f2adeb4aed0057564184888aaea33c5acf7f264217d8097c83b7ec9e68356;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h615cb3098f017379bc5ffbd5c275778a82bb3a7f35442bb30177520f77136b193f5babe8ecb77da71e2a686be9aedf93675a5efd4352367d13992237fbf25882bbcbd46c9215aa48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h760a687b3004855b94b032d9b537a00e39e97f693b1bbc594be437e40b28288c3028469956b407a7000d28a283f53911bbfe4172ae6659ce59069e5380380710c730c39aedbfbdb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8754d3e52655f4fb2c48707f8fdc7a784ddaebe4f328a48e16b84843efcc578b249757d99411f8b9ca80f0d71315d5aa48fb1936021343b5bf4b984b530477d454826f613b68cbfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80bddceaa6bb532f42f63302728b61aa62f6a4be10308f7f28e5bf1257eab312246018da32e4dbdd58c9edce90f60cf4058672b8578691b75da948efa28708e20a651e32f72f1800;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7eb0bd4c5f86d6abcb8a56a5af0cf18beecaef142ccb6a6db3a32250103f0e95a65294b9d2a9ea22e7c51bfd41342b607c6eb0f1c333faf85386cc58effa2f6058ed68b53bd758bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba0e00b796309c53e414affca1113717cff5782e37d94a289a144e9485aadaac5d509e12af5ecf0da2400ca866e1fa2b4646da0c8ff13d2f79e58d122963fe6489d302cb5e13e2ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa82710dc59bfe6db7c56cc1133a2c7fe2ce9c361f3b3b5290cc8c2cf3daf3d7933788630256592f244e2eafa1261a0c969bfeec2f51631c997114c023f32413dbe0fda356564ace;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc90be882f32732b4c85239fb56d2afab2eee2ce06cfdfd3e7eeb200678401dea9acb8a35da6363e3ddbd2fd5347dfbe25846019012d4952baf16cd352ce598deab28ae303a20ae3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31285705bbbc8237be1856286399531f4f62f897f6ada995f3627ee9a1049b2527892d99bb4a303099c70016e6afc0ff21eefa6b22ed53213de6dcb705fd17e612477dd50ab323e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51bf9f04696df87a4d0ff047473f01ad1b32a1819f769b2b1ca9c2344b84b034bd881d99acb0df0de6c6edb23561ccd8b40e87db69f394577ef94acb53d1099f1b435e9b8568a011;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1cee6ceb55db41763bef3b5355e99786fa6efd3245748c993930e8cada677658a55855e6c8023410911f74b95eb3423b7f3d4d320194340e960b420dfd2f0ac443eae16b21be0f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfa24daacdcb5f185f748af63008412a3a4eb4eb485b865191e34a074c521b46a1c818bac9fff9d8e9cac2796687e7a0034d21c6bbbcc8e00f65b37e1265acd41f61d524134b906a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323e8829e6cf59c2358430deabe970c7d43762012d8227c090fda30d0d4f12266e1d7336bfcfedcff8341750b26374ef4dbbae3f21a18b5fb6c24b8845f129dfad47b67ddd06d142;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6d97ada566e22fa07d7abc5befdaba1fcb5550180baec299a63f48e319cf8355825471ef68b1733950b855733f396d8e329fc210706583884a636ec511aee79c420b01c0961b886;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44d61fa551f7cf66e13b0ec2a3bb7c751b389bf6ebc73270955699d21d2bb496e3e1afa16d1cfc61466f39d48e8246e1560a23b7936d18443ab21fe8535cbab62fceef5f2a56a3d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88813926d6780c67b9b26a97874ac2ac435724ab99f775702ee7dbdaa1066f2eaa1afb0a04752ebd31709ec239e9d1490c0f8024657b96a6a7abeb1e221cc2c1492d10978f248441;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb482cc859cf8756e76d5ddf49d91c2ee02f815d532cd9e83a474c1bbc0e4496a8df57cc263b1acd36d20a8cb19c6dece6d52b55bf7110a173e83f59ca4de482227804e9e890cd459;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he102c6b8b33ebbd592d7bdd09a24fb39aec341616f17bda7d10dd209684e13406eb7595d552dd14e57661bf284744981c252d8c25720e16d9cbd61344af26d924e9d30dc301584e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d2a650d239f5c870a175c9394ca43095bf63d01903f5f83902a68cab54947f9e90d91661253eb1a3ab9891866d8670e8d28e6ea2c82636d5527d5b11f246849a581f25281942f04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31501129cb5477cb785babe1c06683d7196168a8fb40cba19ccea6e4ee16accf083d1a5b868f8f83c5166436ec0a7839b6c2309058d6c7fbb199454ef76b28bab123ef850be0b1ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2a327297788aaf4936abce11737fee17892835513a2fb0c69ce06a7151c69c404084ff61d2b99a16fdf76000542786d1c7fcfeb6b68bc93f2d75df4b31617e571435d0eab67370b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h382bcbfbf588e240ee0a8c5f82f582b8175a002bae6a533a921d8b0b27a75581566183093e8336ecc60784afaedbca03d16a2206c8385431791988c196afde0ce53ef1bc7db71f08;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc17ac74a55f9f83659d2362ea7da17780ab7fb4145a3b3841ac752b1cb8faa25ba631f404330c10cadb44fbefe27142251fa91f0f8be5f642700c1d53d7e91fa878dced79b8c7eea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3baff50cc08bdaf9f8463eac5d48cd3d9b633f2240525af6e9c4c7e4caf7d3dd346587e57c84ad2ab75bcfc76f7c78ff8d1472df03c540ae3a53a6ebf2cf6d9db2de5c95d434b088;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3b0979ba581cb82d600e32258714d2d5e4653b0f614f18f92cc1e3572569b6b4267d583b4a57d82ab0179f8a8f0aa71fb9762701ebecb4e48980909a4b8d9b2fd981c6e32a09994;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3b78add25edc0784765b29bb87bf7328f16f8153bedfcab45f610681498e7260331e11b20b3c5963353fa89fac9918e73f709aac1900934dda8a8aa04f094f8beee7ac5e4ebdb9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h552d240e35ab997dfa7c0f0141493e715dab16ae5ea5246df3f530053b4fa9da599d3bd8fcdc8a206b8adbbfd63848d0149e547e085b66f169f035b95b3ea8cecfa5fd034c6bd5ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4598e21568aa796d0d4f8a344502d644917819e1f838433b9f6f1516c6ca9cb569c44788b452bc561327cc9140fd8f3d5d9438781ba3f6e2ce4ba31b51b4eedfca90a0e5c0a0e53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18e744abb81eee7c8bf8c07a4a307e95231fa816b256e5d7a078e084e87e8fe04d4fbbabbd6b2702426a28fcb45e96d0a37ea06f1e43a589bdc6437adcb49a6dc5ba2f9aabb63aba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h516406ec5c9e693140fad65e685bc503293b12957b942763af003bef7a0da9570fc262eb466c287f587212491d2fd7263a0e69a28e624b22f7db5234f61629efb6d09fac9e78ab31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5d1638ad897af36380644d10903b07f89cd383cbd332cf634a5680f283fbf82f00c5f9a1009b2005366d7c98f5ddd34cf3e67070dd94e1bd7a9707cbe9b5bda599570ec9dc132e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27ed260030ba736304faafcb3905602d5e0a8872cd51faad4d1d8c4d4d4229b34bfe5a6550c55a8fc68a73e6aac5b4eaa5db6ef3013e55602fe52fdc8c5e885da78109972861214f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h307d82bb096ba8b19c1b99c4f539ffe6e5e7f91f40048b6d6ac0d65d1b31feaf9d6997ac6d4b32433e2812c123867182b4da5e8525683694187d5380dea5fe799991ceba1c523cdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fd47f49636a627cfa4e02194f93a1ce7ae04b339de86fca001c1925bd67a0cfd652f21e7f9aa74f8b85a223fcc19a7685d378aca74483f75693aebca2fa252a8c712dd28e5ef24a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69bc386714869cd4c85f59b32864ae5fbe33934dbdef9c2d95fccf071f265506b9cfd0960322224d72ba07402054da3e6667bd21ac72313cf70088f279b8ca90d846ecda6333e8e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57052f4b523ae32a1dae199f6f3a284538536b273b758a6fc1223f99c5103a7e81d5f3a002e7206ca01bb7489bdd3129cb09fddc0078743ef5d4d44f5d5b869fb116ed105b5324ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he454a56ee8eed697c7823a05eca4c6961971f3c9a502394dda33c4c949d3a79699b11283b0f685e92212f2f2236b7970948549c7839daa3a67f365c9fb0177624eb605b2bfc40a37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c37adc31442e131280d77761181376fbefe22f009ec46ffab984e8803bc769bc96d7fe0128e7f68de85ecc17581daef205d9391a3ba4689b93f7d52ab27a8ce87ef4381b2dc817d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5cb61f7371becb1d1a792c6bad7fd58c3b04cfc92ce168d448c84e1768b210dc5a643fd6b616b37db56a9020af67c8bf22d5fa9b38f47bf6a82b6794b122f88d3023677585f355f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f7b65b83b979a7c206d9fd2d4c8c945d6e92e638ce2c129642f0950da9e730a02a194d4c5e653ae332a991ed747c2cfbfc246a234ab7f33dd6985a0d91d94b55608e4f66b7aa97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26f4e65516a7eeb4899e58bba8ee7d3d90671a031b72f25aeeecba18457a6def8243aab097906d64d835419eabf6a99f42665ca1e81627cda875a54868fdc1b6046ebdcaf3d0cce8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25facbfaeebb1c566a536c89111d040210016326098f70571accf8a36f32454d3843d61e77adb6ccf981627120ed6f7135e1576dd323c96bd59d61c088ae9c38d2e83a6ce791922f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa3fcba00bda81595310f146e6e156196ea9595b62574942bd6473bc9b7aa8b158c0383e84813a4d4e1a08d95c4ff5a4f26f067241a473fb5771b4b491e5619ac12a3887bab17a16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha14d5d8e309519c5908509111eac4b00cef12199c2f2a402db2c4d4f2b94fbab5ec5def4bc5f028b6e6e41cef5050a2586119963d050aeccbfdb64127cd1afb2b593918b6db80ca3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a4fb6b80fa38472181c6027033ce1df7803c9c4b36ec5f674d59ba02b92ec30a17097ee0d5e84740f7c438133e4c8f01e3b0560caa7feda61097703aeb226ff38ea39db37e4b09f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde410ef83259f6764bf16500ad8e3e058ca784a31d29743654317712cc3e68f0c8e94d0b7456b72bd8d4f9de761aa05e3ba0284a58ab19d5bde205a9fc21d08e8f497666601d3ec5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5842193fe20e28e8b4bff5dae2fc711f63f352976f2e82184f276a1795a01b7560fab6bb0e1e5f3445143aed9984d9bd38a4f263aadc72d28ca5a09b61ad54ea1495467f99e45642;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h795242fbd0edda10eee60335243295fb28f624c73c34928fdf18805312fb031c28c95ce87efe3f87819aacb61cee67794739a245f1bc2535862daf5fad574908458000cbe00ca959;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfe60576fd8e59ee29a98b747ee765ca61484e76bfccda578d3b41323f92886a3280f427b0776aa8d58cd108f53370ed11504757341efe0905716fb3146ea5e1e2acb8f6c79fc61c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52cec5603965765219ebb67f0030a203aa3a6c6549254fedfcac310a585dda297d7d7b13d92dff92473944df33cf7b07d907f87b6c60b66db5167df4224933b5b7e924ccfd990baf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47c790cb7d501da51a730e368edbb9b872f60c0d58d28067c9dfd7991b07a6f426581c8993b196d8b6939e3730abe03fbbccd81dc602a639188eeb2abd89478679550af1941e9369;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7b1aff410c6fcb69e9a90634068772c946d959c3a9d25431160717e570ce5a7d61c7cb657873fae22c695215ae5a4cc9ab8e30dfefdc0352255489b30ab5220215beb1b9642b845;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bb458aaf0a47d262478594ddfa734a3ae1c0c97f9849fb1cd34408404c9a335c769f3ba1ea36cea7bb5528356655370c2828f4e9d9ce18051610b85940296320bb9f5c45e8650c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb782d086ed7a05895def0670d4dadfb3b3773390c147a15ec5096947e0e9ed678bb2763361a35f0f423bda6b584108f790dea72af9187d194217f1c5327d7abbbc1bcb50233abb21;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91def77c0ad6becf191e71fa1acbc0519dc002e200cf582cddbb840e34a32cb0a585c8c0af2a751a0697c383b5c589b1892bed401a703e35f9baf74bfac7d8986f91a5aa71d69728;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haefd5152e816d14da71634aa8668ec0aefca42eee003285130924191a7b0c4118971074319de6ad3f8b19799b26af9bc2ce0d2357c6cc24ad1f3742a13adafa8fb5e6bc262694c39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he616434b66f97685d6c311a27c8387150231dabbe0535bd025afad598ca5aedc76bccab3871c68d6598796194ff071f0423bf5ac4f31e83cee2533ff80126d9313c12f45b0ef1d16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b090d8952f10fd416b1ce31a8de6ed4df9ec0257b93f67119e592e2b9c192a4c75999f7900cd7176cd9de17a5c7fcc080f2459e93b1417486cd1fbd63e21142de235aa2b6cd3ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b8b18587b0d02ac3aeee7f3e9f5ff65df0dd67a17c2fe04d3af69cc4e44a73276646549029efb97332b6c4ae81590c6d83ecccc6e2cb633bf2f018bced77390efd380cc5f39027d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf49c4f2b40e38e99f121ef1a1a0bb98e20c5e4243d4ed1632e9936abeb78ecff2ef14df9875451cbd6cd79557aff01ec5f46f04a53063e84be62faec69f2b79114a16cb1f0fd478;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaa16b4ead3c07df6fd4591153290a5308363da76db36ac66fd8691564bc2a34ce2ff59b514f9e91cbf2f22be5edfe784981df604b72064536c5899e800ec90c59b12086276e4041;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78f5818f625f0c46533fde1d4a39195945143773d35a6340d1d9577961119fac1cb4691eab0603ff2cda46a5ab4c7bd6b4b46ffdbe7ccbc4af04f38ee460b27992b4af3ad624513e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h502ebed9f95d04aff67ccafaa636d1ace6054f0f2e8a97020c5437374f51c7f8261cacc67ab7f6d2dfa29223be76bc66499c914355863bbc61dcb8f2fc3e75b76212082b5aac8385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0898dc20f44c9ed7aa35443a419499e94d99a9459bac6c5a604a24a56e6377963b76bacdaf4cfe05695423eb0024729c4f8ccdfdd5f1b20166a8c02dd1dcad95ecec321fece9962;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d7e10b323517861d9ce0bcd980f0b0b80e6f301f08a8be06c63774e73a18d1443308b07fd3734ed1e0ef03ac990153705c5ee7e5ac4d359ae61d8f00e6547eedc07a05835aa066c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h321431757882dafd0ecf2eab5031f0cfdc6e558df17a24d15b4e7e3d1ac3f67663796119bbab2ec5474d437395535caa424dd28346b0c7e2314a51870ad0ed687219c87024f0b62d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4101f1b4618a46ef7eb63226dff53f162ee83be6decd5fab344c329766764b34347aa3881040527c66d4dce74cc4c39a57bef8b42fb98360c6ce33a513b72f185ed7089b00fcbac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6790d80caa2843cfaa878831f70b5fd412ceb1261b6fbee23cac7927a834907dfc5e650c9e6af8074909dfae08508abb75f21ed0987ae5d84a3fdc4706ac7bd3e16ae299aeabb6eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef97a2570898acdd1a1ce0271ae1b1467410e7dd2db5f131bf50b7c16d3f065f8f071b80579fe51b17cfc0f951dbf85a1f51833d81badca47fe0c945ecb839ccbc6a5f1e7138bad6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3472128e636338ce1efb4d6e1b727d8f440ff52bed43c066f8189ea3fa88983510d1b5ddc189540cf3ff82238f74818114d82b1807d5e0996cd835346b806883841591eda87b045b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dcc8e828280975aa309f03885b7538c99c5b394280b3544b72e2e40f0a7f1190f1d373f71185a2114088fadbbc8e918ec0138480368e8c356823eb6b2165aa519403d72b45fd4d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3ea93affa2d307e5fd6a7fa3a1f1c699638fc1bfc29f2caf74b25db8ea01d3161f1b3c7781434177effb0ef18e12fadf5db20da5a02ea88574171e1f1cf283de97a148b1017f94c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9bce6431a3808ca445f580b3c39eca81befb0d58b89cd8ec8a49ddc6ad6760d572743e632bc9b2f2944415c680d64b813badf53974f1b09615177ebd80136117b052dc3a2e709cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb4d299ecaf06f4146738a3bea5035c2f7e5723cefb99ff8eb84e5077b710562f93d2d1ee2d7f1e18e02e89d61f8bd1cf5ef175beb9a4307d21093c36504aa23902b6266ce935edb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92786c8152b12d5adc83666224ed05a04c39239933c8065f7afc881f08e92526153b25a29543a84592dc0e8af43fd2853a32eadf7e4165c7ad4abe6133ca79b8749edac8f227d5d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87902dea0110d9e459499821ad177b20e8ca15e9d03883f94a10a7dee811d828f66c5215047475a8045d19943defdd722337ffaf5c3ac4d71bf5ef048fe84c81b6dddc3a2d43931e;
        #1
        $finish();
    end
endmodule
