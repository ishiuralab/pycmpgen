module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [19:0] src21;
    reg [18:0] src22;
    reg [17:0] src23;
    reg [16:0] src24;
    reg [15:0] src25;
    reg [14:0] src26;
    reg [13:0] src27;
    reg [12:0] src28;
    reg [11:0] src29;
    reg [10:0] src30;
    reg [9:0] src31;
    reg [8:0] src32;
    reg [7:0] src33;
    reg [6:0] src34;
    reg [5:0] src35;
    reg [4:0] src36;
    reg [3:0] src37;
    reg [2:0] src38;
    reg [1:0] src39;
    reg [0:0] src40;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [41:0] srcsum;
    wire [41:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3])<<37) + ((src38[0] + src38[1] + src38[2])<<38) + ((src39[0] + src39[1])<<39) + ((src40[0])<<40);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8876c01d061fbeae02890988c496bc23f0d1758e5ebdffbb6ac966c85d2fa8c9bb9554943f7b090a69e6ef4a61845871bc032e9b069d8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h713dcfc7ba80fe3fd28615f937ee63e0f225504b7e1220cdcaf2709c9ce71273e44802e47e95ffaf1c550a99ded3f415b3c623d549f609;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6331fbae2851aee6f7e9610759d0de75e195c6b2e4899a11dab948d13c294e398e092d7d8cebc1779fd97cad8e62e8dfe5682b9c860724;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89c784641ceaa20373f745a187b33ae53c2831573f61e932c4d0d63c160c02577260a723473692afa606decd817b21f75ddf8e863fef85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeaf53ec512eae5078b318de27cfefb6aa2f076790be1f291ebd6a17e383b78629048bf4f62a4b98fd842b71d181804f17aa57d86b4bcd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a9775a4dccf86dc1d6f0b584f7cfcbd6a9b548698cc044415926f2cb678a14261256e46380efcdd79454411880c6b468330536a91c962;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cdabfe1cc9e601b0a6fce20868a3c062316619558e429b829863231d67045a625d4bd10d161238b8dc496409d2e9dac4f9e83cd2b8835;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ea65dd07df6343a20eb91be2c7c84dd5e96294f105a709e2bc0cecd08612493b0c7ce6c00e22cb186f7968b1afee91354022294a7c81e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18df62fe92ef117b5451bdca1b98002a45785cd71fdd89eaab7d60c1e99a4bfec323e968477d0bce6c3b56cadeb2cc759749356d1c317ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6fd996e14240d6a71a86d64c4359668d84b2a2640151e396b7ae8fffff5796d128154c1a8a8b6f0a7b81c737ca33f2a781e93824c5b2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12047cf9f18bf8f91f04130f15d50542909e1b79f922bdb8be18c651d02d6bdf81d88158ad18c213864a4ec07611b8a6eb02adc82aff121;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17357daede6c6b4ab4dc00ae99dc357fb45d6dbbb9e57fe2172e5aea00b129e4a0d6a42cb08e86b51f06c92203b40b526fa166dcae76d73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7c91b758e4c53bca584d59bbb4f81c0a4d84267eddd9328675f1cf616f3810f243c93e9e15868488c4a76dfd51c856883e0237aa2aad4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11dbf50885bd840481ccbd4ccc442c94f21ac64c00d1fc5ac1476b2dcc18f099eb7ed74ef8d20de4f927ec866b70bdac0c708e4b6dbaa0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120481d18e6d6b1c24e62a0aad20758b6d1c716219f2c52d06ad907afa61bba291549cf129861327ca87376725b6671cab34564284dddc7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ddd188dfa949fa7f3adfca8461dab7de683bc238450cad7264584d65bfa084b7628afb95ec79528e164c5045b05e31c006ec639e4d454;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a6414c4c35d4d03ced6985889b497bd32acb5bb6fb8691e01df43e05692840949747445fb3892339edc2a2bf01937ae3fcfd86be88ece;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h727cbbb121b123f3001ba67eace3f867e66499966819ce9212eaa2c00e90aa3176d01db1c4870a8d32336d8798f61df1e8d4eb1d9cf332;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h881d438f1415f01c4dcef1e3863e2117bfe4d25a56ecd2244561a3445dd3aadc372f5708f11d05be2e3b6cfd466699ea201965e141f9cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d15e8fa02bb44b9bfff139b0eb38373320142e6112efabe4d12cdab732243f01a021d4c11d95929212c6835d752bb4174576c5ddf3568f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42f8d9eeee79507bdd3440628105a221780faf6f2ba8088177bb9e5a031310c2c8302ce0feeff200e5a04ce969c341b777b12dd24d3889;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cb3bf47e8b15ca48bf960624229bc77a7811adb6ace49c1dfd9f9a62012af6f16cd66a9132e81f66ad73ba9e621587efe88e14d725db8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa71131002e17f545a204d5a2b00e52af4a83031bd5ce350471452f52406cbbf713af48febcd0dd6148d67b1ba12851287a3fe9d854b66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28d4ca6883103f8b7e6cbafaa9a4fa3f40190ecc672b5082923b25fd50767644725db20550d9067ea2d7f4e30ae8bcf133495b3f1c27f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3dbf5626176952a98dd23964a6ab5c1d7a55747ebcb996e7ba52945a636a7a8cfe2a4254af46f01e7ac536a0ec0fe311578caabbf6aa8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18bdc56a0478b21b8131a6b3c13db629ee22c45d24f9ae959fc561ad7c4666198a0df64034cc735ad7e3f34c952db7d876e0aff3bf7cbd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b7cf20312b25d013e6d9e062727558cf7b706e31ff2b89afc3f90f0d86ab78e3e54344795ddb976e3c7f4c1ed4492579974e77e75c8a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he19dd3c12e7a8a6e0b6bf55fcae491f8988699ecab14b63c584ec88bd14e1a500c34626326776df599bd022f3084468e5f86df6c277e96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0fc3c6015e225fd471089e9abc8d71f188f3c16a56dc2eb799e649b7e57179e0b86f27b7cf1ce34aeef78abb11acfe852128c937d48c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cd6813fce450a43a18c81e7bd3408d92e9f923d5321897e363cc749dd2f0edd8abccf983a107448febdd3e86abf9855a233dbf971899;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc16bc14c2cb5bc077ef4ae4cb685bff58b18d0cdb210d1630d2c21996688cda02e7ee7d4dbc1d4d2daafb545754eb98c1ee8afeeda329;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d20213477438c73f1f38f25118369f197de4e3e4aa8be77187c1bf4d1491662f6b443c429539db06e1b8e2681670009d3982deddc55f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ff89478edbcc4c4ade19ad1a45369e8ed274c52f6c02c5583af6b59bf074185f98b153eae00d9babd37195cbcb69c2d1088789a6a19c47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f7666d25eadaab1bbf45a4526fdfa26f38e47b358fa7e438d7cd76c4a3474013576563b1a14d858f42d22f94791a77a75b55b94f302a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1141c1c6a06804864706b47df2b8de0a06798e64ba6dc273c435b26bc510d67b8496464cd5b715a6a4a3784710e030b877020bd7c840927;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199e43f9ce5991dca5f5e353ff490ad45652274ee8de759d30e0fdfcd36a441a47569de2662d820f059eb5eb123f21e92f3bb5e04a95a1b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2730b97395bae627006261a5d9bc7002093e5a2ba317f487ffaef45199d726fe1eaaac98797da532176d4452303cab1f7149c6b89d664e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c1ad9ab72c5fcea7c6a4b7e2fc217db71cb78266eba49243a744ca23cd7eb7f184f47cbc45f00265fbce61e44241a20d632f59e33083e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h810ed4f4433f65522a366401c180c594e091b879ca2758bc72b2afe4856a3ba5ec5afb292ee467fe673e94d72a2b42f87623e4878227d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f81ddc6d61d4648bc246404119baf99baf1104437edf77fad2d6bad549e45873d7d407f49d6cee5464490e82a379330fc9fdd9d24173d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175b62ef06e68611a4af4b35d36e88b9d1b44ec77f33808679cfc07e57b19826065795fb55d9cd16b5241f91a963902d2b93b8eec173806;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a26d710be30a771c14245fbb580ea2fc75f4f396cc993d348aa99986dec6088b354a6e141ec4b84b338ffe0953165c2066c0b5f83ea62c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed9c35aec3590e5915f0b4c97d3f9e3fb5100d74229c8c9280910eecb857f9966480c9a53600e56f450578d3d085bbacf3b6285f7ab8a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b86a8f06006fe5a54053fd6a62bddced64f8817f097c4194a5d28bd900a86049b59c6c442ef51d300411d3fedcb2273098f10a4afbf10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c894393b161f841d80565496596beb10154ce331326091ea01f3f5819818d89cc804232128c2762183d73dd2a834e0119bf636b0e542;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4a7fd2a63aa480df408554ffe73148c192c78fe2e7bf56fb50133ed1ec74db98babbfc81337a162f884dc76e2ef0c56a9d96f514cbaa4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h983beb4b20fb7be15b9c05887fbd64254eebe0dab67c6c4d7d0fb65f50da77b65029f48f0ad24d98fa1ab1e2ebab8e4866d4dfd18bf6d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e170f139f1cd0bd61eb5fa6cffd5454cf21c5e080921f6d288a9db5fa58c5c01f098e52394d46f03a4b3a563e3e41fa7c1450c3e7334f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8859849aebbc8d2f30bef63afbd87dfb24c47bfe56311485695add1655d7a098e7515b1f655e32ae7fa09a836071d381fe949ad4b046b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec4e76bbe5852051af51173dbfce5674b7c8b37fd297cea2b888180c1de9cb92a22d990c9ed560611aa96598f687ad9f873b03702fc48a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4582d5eb4bb912019c91e59acd2b7f96bc4505fb504c8c144f0fde20cdbabcc36a61fcf1acf1cd527fba987207de048509db03bf5559e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbde6b1b522a18dedc20a8279d55db17dce43be7e1bae71a2694bdb915ead7aa1b5d5e450412f07fdfdf98491186b111ab393a98fae68c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ee7e3ed2c729c2fc48020251af209ed8047e5a5261037fd39cdc5352953098f50dd41bccc908c73e83d690bc34895cc2ccc10cdfdcfea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35933b878287468ab5c2ec7ce5c186894c04a0f996305e4fee2081893c38ae93c14a43b00dd36530c1d05275f20434d8964aeafb8ac941;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf3c7a9c3e7358935122325e309ecba3c43a1bfb7523e341e54f55756e56a2124be5769137e4e2bae9ffc86ed156993ef511071e0a9170;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ca4a9c03735ccd2d8cbe773a83de5e73c910b66ae3db6d18e522bf8384b353de334aa7509ca636fbda4347348fd790112c1f9b59c06ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22bb424898f9156e7d4afabe91d77254fa858dc7a9f80814dc9fe403ca3677a9a5e92c49f5f53f345b4378dac8431bce2696634900ec60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9fae26a7b3f2ff2c503088eaaa4abd116bcfe50426a4317efff52ae74e13af919a407a53b9509e80b4d23b7bf2e80148611819a8dba1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a787aec4af685c7c4ae94252c4d58e528f5adc17b30ac4780717331bd6670416df2d4bb0ee9b6a69bc3c31dc8233f13ab11d594e4d30f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32a84b12966cbaa1d90b595c2503de20e7150bf500989a6a674dfc84eafa3056c4b140647bbe835c4cbc35dfc489997f9dee204fff6c8d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c307ec25615d0d29da686329b1feb8e0e52849ccd8b1a3b89be45e5e60470b1c05985a63fcbfe9565520295acbcc77778ba60c941c3be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ee93bf398973f806578e96b33033ecd62908fb0aba742e191828663cca60a5346b1e3daedb7ca81f8cf8ec3d9a3a66f03060252339d44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4e0998c38058e0882a65d6a50d427fa59f635a48ad21fb87bdab9027082b98d5c64c3606cf80df2dfba99245a89d15ee7e1b12334d73e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76129bffc045ed21d1216fbf431938a31d978ab53fabbcb2286f7875ca8d09b93c2c10029f904a7dc43adb6a3514fc87729a713b00d79f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fe7c18c5e807eea0b8f62758de41fc0f2fd139dd38b4f1b416e6e08e79a4c3ecff779afd73b4827c3e660ee26b664c9320c32e9874502;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc59c4579f4ebdbd632ddf256f74e6b0edcffb1ec7167af96188247e1d2a0636a58b4178c04fbd6bb35e20c2277ee61a29eb6f3759983a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h50d7e19c89773f542d008873be493fc198f69cf636a479666adb8a6b8ab3080f48ac7382c12724fba6ab87519e56899e6cf6a1b84bf7b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a371d0f5fe4c4f13a0372a9838a8b89f53fb144ffbc704aa2f9ce49959a2ba89948981019543a08e63a46c4e88d9c7a9522a390b4ed2d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9641e1844bc5fd75d7fd581c678c652d32bb1913b56ea925ad1273a7529f0cfcb427eeed77fdd13f72357fe5e009c78e15862a722a2f62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d2cd2b32248317c5c3df754fd170f52b8d93f21eb9d28da8e9c8aea676e3e6b08a2ec34fe5d64664f58e64b37ed057f1151880dfaef84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hffab89922edd79f9c068f144dac52814356fd36e96335476ab817d6513571fae66ba76cb3fb01e52ceaaf05d3c428f69da13a62bf8f1fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc748b604633796511c8fe566912c3dfe850eb64a5d89641bcbf628baa13472bdc5fd5f757f520821457b6e46742962ce687a288308966a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa1a641510d0f919ed8f3a09cd494c78b18d20b6a411e2dde4ddc52c8cb95c0ec1313b31d2d275a41a86348896939c7a6143021a44899b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b315acde3db4e0a6f05c2307e431c7b64cbbd693bed34b8b69a0d8230c443d7c62e3077e30899f6f77423a5ebd02294c7fb43839df7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h605cd1314b7fbb2166bf16a80070f94950d16d9f21c88f83474aecfac62c9000e228bd950f5083d46dead4e3bbe6df889ed2bdc14b78bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7dc68d1674df065a1f0e743288fa868ff420210343c8ac6feccc4b608eb8ac2bbe872671551ee9d8511e8da449533190b463604f9aab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bbd4fc9aeee34e190ec08d16c2fbc51076a919e8c97e318784d53f4e06c084eabe0a41165286be089c32a3ab7b2d211b4a752b8efb89a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f232b03af60d7d879aaf01666dc3323d9ef5f2200a245d57b9f19f063f88cfd0d0709746973383708ab9e69dae6ec9c0cd3519e9b763f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1d0359c821ee35eda04524309fb2c4bcf7fd058acfab272e67f4fa9c6ef4c34407a51c40fead540260c54ef0fe90f2b1f5914aa9f254;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163ce22622f0eff0059cd7bc040701b152d93c3df6696cbf0178f0c0fae8a444a216be15afd16c8d28b20fbf88e39fc59e57bfdca0c9d87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h446a541ed8609ebefe396fe8ed27f59512d7123808c1344ea91309b13bb4e1f18abbc6203bb62f574768f991e57e069c3b57366b6c98f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b363b2859e84bb6fb5ed660489f04af1bd16e1cd3dae825be242bbc7d27482271f13eab661401938d376ff0f861b0eaa10077f3548c8c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179c63af4a4e01beac33df338f59dfdb5fedbf5efd42416be1cad01beec910c2aa251e261ba2f239f622c4ba3bedaa4549e65953b0486f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e92db23400a37f547a2f928e347da840d661b29de2dc33c9c3f69bbd11543ba2c813d6e12613b2fc746f39551c776cfcdcd31820efa5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h743ea0bde305d2587a42ad8be8c9851e68cf3e5b05807c5cd4739cf90efce6782832f91c7d5505995fb51cea872ffdfdf426d4b382bb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd57e4e6de7f381c8203588f28d1f3ca1fa22e32101d0cb6cd270c7c05c940457dba5a5cd8f43fc77461c365acff96a14fc50aa8f15362;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcbcad78220985e0f5570750a589118097c47bd8956af15017cd657c7c7f2bcafbc4a3f5fd72d974830b8d4beeb24f6dc3b34b3c6c5ba5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f04ea21c3edbd6f9ad27857121e01c608c8e9df0e7a12433cafc3804ef5d17e2d42898f796b8ca515000ce5f8181bedabb2f0042f806;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114d06d436c16a760ce755c344ee7aafdb526692c272852b326098dff6931e66c505bfc756efaa11dac495800051bcd9f5c710573e8ba6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18911f6db94a13a3330f01de3ade495c58c883e7711350e639b5877e06e22c5283147c443b5ff4fa90679b9026cfc1f3fa77cc8c6c4f084;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12937c8168a33c51cde6ef3f9e8501c6f085a29de82d6da85a9922e43026ec497cde41f0d3eb8601e382f1eca455d320229e5ace36499a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b91004d5be02d700dcbcedbf954dd6032481723babfe24973fea634b71889949beceb98e2d1b40dcc544cbdad1144dbe32f01a6f4a8a98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46cf64a482dbdb9eeb2eb38ee13156737ddc3b63ebbda2e35eb7f0c5d5378a85bd609df249f4a4f24e3b37a8aedae13b4f0d821e748412;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176605035e2a02ccd57551c7f2abddfabc5f7644947158e31cc5b4f587dcabe537ef7c99303677d780eec922affdaa2b3108bbdf40a9515;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117c9f5cd0c689c345d14c52655d91e0d404a35617e7eb40487df976d7e5d998b8d4a90e01c07273cf53ab76bd1914563f56bc0044691ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1569c08f7b8fe9722afd3870f1cde3c01144ea877279e5b7201a3b94893ea1e4e8122d7949fca554b4c5308d5803f59d36ee272bc7f56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59e71d3fb7d94585fa6a1822b0117ee7eac42c37ec9c03445712e8da4da382f1d86e27a8a241ed4a65897d574221cb66f9983388b4613b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8aa239c08621e9aa01475a6c3ad6911ff266ae5407631c1d9f3e62603a3355e548e803af1f523568ebb3dc9e59d9f9ffd3ed6e4406b052;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b9922c24f20ad69a01434c89e21b591ddd0d50f07b9ee54297b2b9fc29e6a3302909fecc1c886de4dc98573c1fb54295c3fe57b60f8d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6093e0f701753bbca86ac18dd070621e38cb93b7b33148d9bbfa2a190d84ecd5b3f31a830509cd8d62a5a066ab1e43cd52f27748be47e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c1164bf8ee943eeae1f0d8f98697b38725373d9bab67e4b1788820f061be82150cacbd12837eb17d044078c279131b691fe2d5a870a92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h579931647ee155e776a87c442ee7f1fd666c322fed366ef4f2d2682a57602555fda914326bf2760a904dd5d4010b5fb468decabb6b99f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df18c00ec2e765b7d0d727dd4bd6b9c06ac8148dcf11def25bfe6ee5a2df5fd1a33e693dbb66d0572b16be7b38e2a1328183c5c235caa7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ce84c6484cdeae44016efe433f627e0426b8e6017b92138563214af46d3be030c8ed0130b714896d0e54b616891b58ef4bdc6abc2159;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170b8659dfd07fb3be3549bf7da31bc1f58650ab5a1e49c2d1a26af198a3c3af6161690e09ab8abb27c735d5584cb629e24b40b3b60c82d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h626bfda6c0cb90f50e97fc63a4d33b4aec153d860f8e9273a2f6897ae3b28010b7be927e4daba7665f068e021e2da9da0e6b749f5811e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d6edc1c227eacb4b435bf0bb3c9f006011f1960a8add2876bb078d6465ae0af1a7458117d17c3a2041556c5ba9b1edfeb6a308088657d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca9d07039be6789f8d684ade667148281684e500befff20fd38bcf23fbdae50b580b32d0a1f21cb382c37b4e16eef8796dc14541cd3c29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ddcb693fa6965665adbcedad250e1107577a3db63b3f7395532f14ea4fbc59fb4e5206915636303f13bf52c10bd460d4d60fe26703256;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf192bac95fc8ed52e6c6b5b648f5cdfcabfb180a580ac7801e04c26e30cfadb4f8906df5863b18a7720147f155973e39ae67cf29f42ea7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c724c295e50848465f732687ac4dbd3909490fab68e7751c288e4de038bda667103a0496e7330d913405f1fe54ac4e83f265ff59f1c64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170a8aa28249a272e2751876dfdd2788559df0a5a5f6bf560a6023e07c0ec5c0d388bfdfc9770a76db88253cb211beaebed0bc4b0259701;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cc870566c0d5a525c3978c544bade743b3d98bfc3f3df10e2a8c85355aed2285568fd31e7ef97b0885fba0d310ca0f751ee7201fdab31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f9b00d1d84f0a35ac01e01622cddd2e8583621312d072cada2142d15fc3638bd9c1df975b8f64b5922caf20badc28e7cbb9d040b21e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14783e1a7ec721020798e529d0195ee9f02d824cab1d88496db1cbf19c622bf7bc50056b9f53881f81dbc7eeb3da25619d41198e43d1f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a3064c8d8d813913a6f639918f1eacd6c809ba9e1d5b312ab04505d6c271e81fe0d746b7de79d2208369fb6ab266d453013a4e9c986ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h707049e2a90e7654b59da44ca63c12d4e9ef002051c4fe6b22a81d497837de35708d1414c175e7a4bd22d14f1295344325ceb1ff67a761;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46a58630e10fc9efdd3fe434d5fd2c643b48b245f81a2fa27a5f09fc8a627e07036611928418a6a89094b5caf8991e66735cbc7fd4f280;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c26dffb33741436b9c5f36ae89cf7d136538467380d94ef8fe0ea4a30d8e0f522fe2bf9ae2af842d1eabf0b5fe4780afc866aa04ad104e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123083b18fdac0a360e59c094f164522edefd833133b68887fc92e2c8ecef09a32405c1dbc7276a784ed19d2f9eb056045ec009b1991963;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dd198463c3fa9cf938870f61c05bbec811ae56180f1de600a54848f7878b550eb443a43b6bd34da976950b04ce1c7689e066b22670558;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc2cb6ce91dce2d5133c6e6b7dc053b48dc9c3cdbf51cc41f82ef616801f90a3ab688a5f0f40124c3c25c68cba642de72e97cf377344a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24a4142244a72019523ec6b41470968a0fdad499ea811bc47b3f84020e1c82b16fdbb722ef782b8b5f75074761b4eb5e1996b518a33333;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f2d596396e2420e50d785c3008d155b43128fe1661dcdcdfa8d7b6cb80cc0e474b0df829ab8dab5d281779535e6460b641dd091cd16b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha80a44ce7fb3e35cc0fbc42eed50b937339766a9c60a924d795cca01c6029b9bdf2dc970233636d2f989ac760356c66bf69d584f6e417f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157f190baade2dd50c89949b7134863a68da6d4585847c5afa8a424cedd5dcbbcd7c560af812041272b03c6c8f77de131093ded4cf47aba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16947d41eb0aaf3b7fdb5d554e0cf7af4483e506b3a9b97eee8f3313399f456659b00a5e8cd16ba1e3697848214a2c62581b31d37c04350;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca25d626bfe70d315f682672cd9dc4c077994fbfcb345321e4642c6abf4b4fad690abd439a939477bd1fe9ceaa22d882e755cada40a40;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e42f5d4cecaa8771300014d5d5143a32eeb85508654478d770231c0f0cf4ad4b8d3a46b5638be340aee5a925c64a6c67ba67fca0ee1a13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee16d79a9fe44f102a6a3de668435161aa26a4cdd0180d5bef3194a02172c7351b1ad6584d9dd3cd0f27cb6f0c9095c99030f29eeac828;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139803aec44d73234c817969af891eaf5da02252e5322088da6d37e126d22bc78f6688cb46c08df72e8914a094254a99441464d96e86a56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f59a9d7276f460409742671407edc3807e831e7eb4d463232394e1fffb5755f6de704446731d4282bf147577d9e6d2a30a4e1e3b9af2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1183c8d6e34475e30c251785a919d20062a6ddc2582764723cc8e4d6201710ef20b4adfddd66205455b437a1b6d08c8a7fa1a6ff9488ebd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163d864ea41d5f13c44f831c87ed4de3384eec39d4f9bbc83734cc1f4b3b7b81e90e353f9c56817bdc527badfaab6f067b8f63401cee2f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1159135b4c3ef97cf0210a65eb85d47e975bba78deb03ab4ca4e1cda5634d15dbf82ed03f4d936789accc35e0d6337c09803ae623febe20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeba8b86df52d23a17d6576ab728748d077584f40477783dce781557552ba6d55f73fefbbbb6ba0f5f0c9bd18d655b69f319a72d39da47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he48a7f7f1e6f7c41d4e67bc14cd0efbee0c5f3021d33615f8c5dd2559e5ad38e06a39a15ea6622b070f68192794aabd0cbef5f50166162;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151f3420cddb9090ad953c82487014917e789effccd6ff776d60d64d41b6aab1e92d846ac57049e07fa998db472654c6875c1ad6e941683;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c373ed93a37d664f2524341e3abfb690e40507453d2122135f633b6560d7375a3a1cbc99520e6fd337bb33faec2d9151d7f39fbd7fee3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29f1dcd7ec44114fc9a1d164412d5b6a5a102a39b085f3cefed938231ca8b6ba7083555ee74bb929918344367c32c271a9e42f86d9e48c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90a0d40a765789ac2ef1e2149a6b51011aa4a867b911f4d8c2b56396b7aa25bdc4d341daa6886bd5650b3f5c77b4822b0460faea929c64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha18652a43010c60dd0dc0dba92d7642f69f99f5c538c71b2adbd2ba97258ebf47f1f5b8e6d891d5ee9e2e33fbf33a8f21b5c959fc5bac3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e511a84f3bba2e9bdab862d64a421f640d382a6c2f5b91761afe123dea1a7a647ba6ede54a31ae1f95b88b20b54b065bec6dcddd5bfe3d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1314dd95ef7cd7d824a8aa8de208c1015f4e20e84ae5f268169532997bd7265f14d5bc46d6b37b3b3b145a44c96f5a23eea451cf939e76d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13682af9cecc3f1974de18e059281c766c714ef64b7e536e9725e7b39e366c0436ff09e0498f85248805389233b860f5b4a42b7ababa9a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165dbaab53494d97f3780a925192f2d4e651922bd24dfe6ca8b1ad325dca55859dcc43ff43c35a4a4a484b4a94d55bce4122a5aa75e4ece;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13495509fb7b516f6d1a2a80890218b8847ca919216949822457aae677db2b7f7034e698591c1f52152de17bb7f2e3ccac89a74ba886537;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119eaf9b76f22814f2e2dd4e8b07f212780b69eff246d37367f381140b3c2ee0eca9ca222363479ed154fa5949fcf890e42d890882cf74a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he415a34a86061041cde32a0d8219b0569e36b78f021f1ced7989ca806ad9ee3f1ababb8504f68c11348aa3f0b0fa77fb80d2176609ae32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118eb636396ee8448d2f9f50158be5c2c3fa3ccfc81483258f30563c3a46ddfbcc31e4a98312396c24bb86bab51c06426951f47472c4740;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12db724e813801ab5b9bcdf41ad4ee3dd1c013ee2ebf43efa0d505868447c825eee24a089a0a3df5714f2229b8f30e1db3916fc5208f1d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e48edfb7c1a56e9f6255b26935dca0869c7a2fe97143cdd7469f33fcb236db7c6c74bad387b335a77e21b9d627dd6e35a2d83c6fc455c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb47a48b3d4b5aecb1c5c84c8a740b7f3db58635fd9e45893213cfe8b3c5613e5b3ba7c2216723ee81f379f01c5caef05cf9fbaf5c2ce3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dec565299f03316afc3a34a4f604d4a3037324cbda1f63915cdd341a693f9d8419a83d1e17c486df6501b71b37836aa9228d92598005dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af5e3a5bb1cd6fcb29758c9c4dab00e94170d9444ab2237ca9b2dea23d01a76b07c221cf785153e807fd6a75d57d25fe05377394e50a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1ebf49a7a770202cc53ed1120596682a3fa07da126c0df146a004ac5c1f761ba94eaabd9966d53a2c3dd76e37bad39eeb8a2235141597;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h857b2e435297ef5d32c0ab35c5ebeb6d44b434a09958e21bb6b7b95429aab548ce404b56edb40ce4137cacc486ae751d89078877a57be7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee23625c3fade6de0a536f9949a43a33d57e9a9171868fcf9394f64b23d4207802ae1703cf3d2a4514726d8f971d2516db50fa0370d9c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d022a2b9f80fbfe8c4337a25f1198b39b371e9ff627197cf4f6c9f3d098930297fb243ac8aa767bf041311a9c153a8fa17dd356eabe9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149fb6e56e0aa72cd97d77bfa7ba8d9554402e914a579ee98b79dfaba7fe8d05fd7186e1e608f6981d526e37d5f7cad63a86d7c384dc571;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb6b6f67fc78197da7e1fd2549afa090d0ac13a912cc4736b02fc5dac06f77d72108753acf74e00da76a5c865f4042cf1790a7b6180b4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eaad29ddb68a554a3c56b069ae8e58791cd122c6f8511ea9b7e79c3591bada432f653314b875f7d597c6b17e747c306fcc27de85bb262d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h545b11931033b4a7e62e4bc0ae194bbd953aa713fe10875c7ea5f54ae71cba9f2480c3ffd64c474cdbf738c376a081fdc82e05cf36542e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e556c6cba4ce9c6a262db4fd0ec601c916b04fdbe783390331735912f4f3dad056478698a830ce92e8cd835248addc3d3820029046666;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126ef14ab5a737ea55fef86af1e672bad1f34e67eb075a1aed37127053e6cdfb7a1ccc327775594946c972c99c977ad627fcd086fa33177;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0e3debe90dc2cfc655871773cca28d627c5b57c1d778f13056fe786daa7c25ab7333a3a9bae31aa27467c9060578d646b3c11822dc9d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb669a3a0fc0f3b66839af987c3080e502f7d00a754d8427e43a0504f633d1b54004f2b024cb46445b96e2dfef34a7500de36041083a0b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdad6ade060a0d95d73fb8f68c2a0ba2f55b3ae07368a570610ec7c13496d0a3ef67045d9f8aef06829bdce2c15050cf132e71e8cd33a50;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had6a0aaa081e7826bafb5dcfe2b9c255eda1b76bd6ccf4159e09c7797f1abd6f58d4dc974def46904e40beabc18e0567f3c264979398f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he93959d7700591838ff66e54c05410ba91ed7a81f7e7384c40d91cb13909d3066aa53fe55d30cdf09b336afde8ff3fcd3c92c3a96f0b3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0571c0e7eaaa19a8261076efa674ae350e76e9d5c2001e471b97adfc8e42ee278abcca08e5fd63e3427064176398193deb03fa203b1df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e27b036c644f4e4fe2bcf35c0478daa40713ef00d12cc3a3c117376607e058ef3aa6808c127bf81a4405f69eb13b90f5fbf9dcd8fe25d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10828b200d170a4d09c0327cb38264bef859523f4d5432a299a4af0ff7dedcfcaf8c22591a78e9a2c139cb6baa23c3dd8891a7cb6d3bf82;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c5e6306e6de19964117027321268f575a3d40cee54ca3321eeeba83861251eb74377c4ede6a31f85ea19dc4372ce8023cfa3b4ad1842b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ec1f88ae73a8a61c83e618fdb00cef9a97912c1ed75d26d56225336df5c37af880d1bcd201410b727acaef26420635605e2540a499b84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d5fc6bd615dfd17816ac31ba52c377b4398ab2bae6e7836a2f5b5128c281d6bf1bad32443072ef304f4b771c0a3e0e7be270d13e9c5dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9b0c38fd2950e5cd72372ffbca321442d5f06c25053ce6fd9d2a66f405a378a551b87ada1732d01a3bf6927fc026fcdb622eb6eb2ae22;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19099f6c50b65f80561e549d72fa498a9b50d9290a47ed54a7d740e6f6ee75bc5fe4f0e5af9a4138d6244e9eb893b6e856ccbe80c744bd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3cbd0da6c10a23e6dee7df1a164026206f15c29a3358240cf5758f907f16b07957c892ac134dced68375cf4ec9e9d3587cd405a6d4deda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ad89c6983dc9bcf0184010050332429a784b7958093b95d4bc4bf221665aa2284859720b83d9876da0faa5c43a3a373f3c2b8dce737ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ba5bc37a5e3e45d8da6822b202780b9bb7a735912c3bea1333840331ef3de418900390e86b089398a3f89e2bbf81de9b73ea4f431e372;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5e5dffde2c7c9b09ee2d16ca422e7afa7eff3a9438ea8e1fc855281f64f65aaa7aa604a4fb33ae1048c86b379b8859d926e0e50525cee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27f21ebcfa1a1f6b06910d1ca410313dcd286faa0fa07dd78e698c33ce82cf5fd17e20dcd2aac181433493762b633a0c6b7323d5e1fe20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he05d1b74a826b98aea08f92515cdb680079ad66dcd63a9cebd2118a7ba36bc43fcf87d4abd13102785e31862d7428bf43ccd3b846b67a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1384136f65cc559284f359024e6c374b0eb87f637a309b844efcdca9703fdd976118d9534c8c5e052504329ecde049da881889c1a489b5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0f4cfabf1e8544b2a7fbe1da160cfe406615c3e71f3a731646ac33e3cb670775b5aae0fd56799e9b0d82460b5cfff5cb1e6ab175f7979;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h678e15fe71dc83b2f2684e8ffd708dae8c5ec85347c89d687900fc9590a609c84bfa69e4fd92fc107ee46970a2443f03e0cfb87a8ba5bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h344778c3a148f533ca00d04ba47fa4a0b6e50e42422b4995a64612181843ee8490bb07912901fb64818fb74796960d4fa1a019eaebda1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2460720616376fe1acc902dd74c3cce73c4d083d9dfee718793b82c2cfe6cafad5283875094817cb4be5dd220204b29006c8fcb2fcbf9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33eb16fadcb84a033bfc4ce77b8c918b00825ce165405bc0c0fc4664cca2d9cc8d4e586358685a602c383ef7cef5a8811822b474649843;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac893283113ee556b91cdff54b7c8f848721e1911f0d3b5cd53a6a8bb225ed21c1d79f05c6f0fea45e6f8a756b15f1af4e298516e21db8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd5a4f05b6dfb87357ec497e4b2103ca77ac99e9380fe921f33af4288fec73838e4e222fc330b0b68fd9171b920fa7d1a0be39b3054218;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7fd9a246fc0d25ebe150a50843ad5085ac801f037c1d7bd711bc9a5dc557ad16eff3087db19b34ea6f8e552f1d36e577273b50f0767a3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb9bb5851f41adaa3616f5d62697f7244283bb3e0e6c9c2ec9f244a61638730da49345acbdcb469ff6615733f8a0b6dfeb73fc01dfef83;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15174e01d540d2646c56657da606dac62477a794663baef2a42932388826d5ce8332f12042e2f53bd23c5770218e46d0c8a54ee47673bf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c755c0d359ef382e9d0671cbc1ace34a5b84bcd5789aa292c268f7cdd2e479a0b727e90a1f62a4d43dc6d8d41e54c7e85db9783198fa2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc423d8e9bdbd64645a9253b72ed3fa4ff3bec61bacfacb51b11186707ed62df4ef189ee54e093f5ec68aafefb6de32198b0d400a4058e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc50a0be5896029638bea7f1faa676e0ba5578225a843e0f44231c6c843cc085ef4aa766da82e51f69ab029fb595faf4a30463ff6729389;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h837b479e3c6b15ccca32d37be9f70c6ed823bca7c517ab3d93377b24fc6ba09756faddfcceaf4484faafcecaf025666f7a9c9c4cd94ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf86f956995d9371d22c8ce569a103d4e5e7e69b6e3183308b03c745705ad8dfaf59556c123ab65588045c1e3fd79afff291b988639bc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1868bef315bb9e141976c4a68e6062cb2de3eebed26a57a8fcdb62d087e9f6bf506c3b4e026bcc786a948c16467acc8874faa1d76ffe03b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac65e021ac1326442c5561827a8b8ec28caefa45b640c094759a0a8d33cf98f565678fc75c999053bc2fc5581a0ea33fa20b0b658985b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d9485c188084cf79b20a56bde695b644c93151e53884ed6b8e99fd59c82f725f1e6f285b63b63a31c597a4500237b8890c512f8bbd2fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45f1d1ff9167272a29e4f980000fd80d46bd2638773b070284d4b56f63b369a77fbd2cde0a3ab5c64676dcabc13a85902aaa9c5f6cc93c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha07f96906600425a396c422fb7c2be7862925ee683618d530b5ee6414cb6c108c5eb49b41e9be76fed4dc5723460c19447642c1b7b90f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c46899ca1969925a17a35b3c938f5b7be68642a94d110087bfe8b8c8405f5cc1c81e34b9c0ea8877ddbda76ac7fda7cf12160863f5791d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3adeb73f0d2da48a886e60b58e6ee7d0516f3caa6adb8f8c2a267d4f81e5285ad55967347203857e795223856c8a5e5182724b15514886;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc395d0e2a157190d1dede512229d1b863515af0d9e480abdfbdefbb2a04b6078524597780ebcfa51a05f4fb5bb198ebb5957435d7d8f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4d7cae55d5ea50328ba4ef6f79854a2bb8303ccfb3b07d2556aa91e83329f4156ce48cda87b709b72ddc240ba8c29245e403e9eb48c4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfa73eabbf3bc577704e447f7b22abbdf19b085c3515d1b925924dca88b3cee3da9ab11bf1523a8381bd22a947ffbeab00b5ef8cecf46e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc10ec17ea60d7974e48ecee4acefa58a2d70b32dab1116f96a2906664bc3ab7233cae211fd7f3d8028330c62a794e742510bfcaf6388f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15256b1f83a9b91fe3c1e912af4a0a0a5fbb396cadd2aa34f80e4ddc34fed0c831be97fba063f2b548506d3eb98fed183c4feec0f33c10c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149912df08ade8d5714a9b457b080c3ca6683e9d9c37bde15d7790db570013a11d755e26a341b1c200009c334e122f96a41252a314d06dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b959913146672f775f10c988bcb676f7c802519fe468d74c60aeceb4908ac443acffd6ced1f836717635d37c573bdfe1e2ee86aa16cef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48bcc9d8799506e7a4e4519a8f1af2f4416cc4f3174a006bf4a0b3e27c857721339a1001485278b1da908ef6ba113c63ce4ed558bff759;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168b69403599983c6e7d9ea8db6ce09c31743a9beb288ce0ebbce53a5a56fbf770f5af1d4726f3c2f3295facf057635a1cbc8eaa3cddbc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43477ac589bc4994b2303a038295ebdb3968d3206b5cca97a3a5a2f2d0daa6fbc916ec6fff4c9ec850c774b8d42ca84757c154b1094a49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108c0808e8faade3907d054a7bb9c3599d01013e4617009b2536f5f3373f05634613e7c8170b43b2a3f3a67589694a100d745dd0f984048;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60e067f47bfed326629dbeba71f9aa5468f6e3c672823803c6934576217ad33d0269f6268d292b9677eacc8c6d757bc47fa78f858c0f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bf0202d9a0422e273341484f62aa1970bd58ec2a37bbcb72b02fc46cab2586b63e2b159ea19c693d738ff5ba6291b1408d676504cf1a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4370227119323391665cfcf65dfac297a38bc6e57362784b36b9184c436cdba9bf8fd2407852edf4111c170a5040552cfcd8a36474bd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f254542708d23c763c18a69293d84c8899b9dd50a8ab59f2f172a559fc55efb7fe426334e28a87795867aece767e84f019c473719d865a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2975705bf87eac3c2ef9f31f2f34154387e2750fb9fb86b8cf6ccdc19475679ddb3fa0271984c1c7104b6847ed5d5a56f0dc226887c8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9fddebf268801eb8324e028bfe23420911f649471b1c2d5739cf749f32b26a4a1452b0a8841c4a521f696603ccdc5178b24140c080cc2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15929f9b5f0ceaa9a760842df1481e1c781964d5cd1ee65e272bbe3fdcdd898ef75c30c89f4830cacb693e62a205c67c7d2783cf750d6a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a8baf1d2a28c063c0dce117be2c7160529e6f192ccc91924fc9bdaefea079ab519df1127e64da4a861edd7e98343f8481a0330fa2516;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a48ffa6fcfcb6c16810b825630311a4ff5bae10f2ffec51fb90f95fa5224164fdf5e3fe9e0a30a3332e06e54c6dbd43b22007322d28c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa1878ff09fb005001e9c05c2ad25f90fdda2e6b1c81f28f48fc1f9f92b8de1eb7f91489c378377c1b35826d82036bc4a7c11023ebb512;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89103627d57000b9208b7158c422bb5ece2672a7def5064a8b0fa254d39b1024dd02e9fb8a5f769d8549ea1c61f44f8c2d24c5cbcb2c1f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5cdccca7cd38bf6e3a9a1a77229886fa4a6706613b530bdb03b6438ba922d03e2add6a25476cf503c431aa4c8b1297eec4797ee53c58c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78322cb498f3c09e9f9c4cf289ca083f3534dae5ac94e3471f94b8bdf0efe515169f4e9087ee10a3f193d7cfe57a24f22d02ddfd5add8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4b6d8d4d5c7004c64b6f88181a17cb23266f4295b37b257bc1bb8201c36219a66ab5e22060e95fadbf45d9940bd277c79e3dd476c3809;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f14d330dc64ee5c21f7d5602ea6c297ece0d1a417e643b79cc384fc10a8d78c56ae11910a273aba2be285f983f24b3b0548de8269e61d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd9d665a19e04b0f49e967e32e817def4ca9db137d7dca011d228ca1c8bd60a18dd86d21a28e8c23a1e85a5a6e79e8dbd7bb3413b5b488;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92a9bf65e161e36b5c25966bcefe2d79e2ec277749dd7943fd1a36774fcfe53f31b84a324b7b5a28df56616c7f30606997c5936546a6e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb67f02e3d36d3384478b0a0fd5f7d4fc6fa18fb84e12c37c16ed29bc2785637a9c6e9b66e1f6bb70b9161e9f3cfb15fd7bad1c2acc64a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac46817b85a6db06afcca50a17ae4dc5440e143d1908c0d3fcef42b72fb250ae375f1cdd7be602391b3604136300c3859f3d09338302dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h236cf9a1dd96654818e8c1315fbad94a21a8e10ee386b801014d6530d0e005b5f2dd56eb0f0b88af6b09bc42d70905e4dbd50119ae0f93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af238c7427dc470ba75c3a52214780de517cf5a8f827a0e0c663e61237b89bb9a0897b2d4de07f63e24b2fbaaffefe790c3fb63e030bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba072a0d2b7b580f4ba16fe8fa92483a5dad0be30f5560d576e15440497220cefc1fbc64ebeabcf36505a6357b2a9b0be957b3d81b09aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151d66bac42a0a71caaecd22f671f31d294b191b2923b34b8af96ee54e45b0a881796b912b920c9f2570c0cc12d4dcfb040c43b41111799;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e563d87a182a7ee737ee847b38a5493d39347a8ec47781782cc745325ad01fb78093891ce5caf0290de7e0bb03abe3dac6734490e042de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3f09344590e0d336459d8b2203a0cc3d33df2693aaf2cd3214fbe24bed5ce49757ee55401c7e59e512ec71b18a4bb8d0ac97623186994;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ab1055594e1957b3d5512a074c65ad1fb09f7a3c9efeab2f47de1386c5be163d5159cbf6c83cd13c8559908df27a47537a95bac6d5db6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1228a5e4ec03dc849ccaa624ddd464f280af6e01806462af0de06ba3e915ed24af21ef0d7fbbef8591323493b91763e4471f181f0aa8e3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6403183617bd48df1b5d1174bde7423316b0ab07a4a456fde59cd1d8b9ee5345068b1aefcfa4c982fd9cc0f12d6fc453dc990e8c62e144;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heaa1ca38ff2d27fa274b9978601b3f6cc64c70a18092e440c9779b1db2177aa425cccefc74a96ad4d2cd0f8d3b9e1a303cdb8c3c00cfcf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ff48f38ea1f940e6984b1384ae064b6f127c4c5bab244456280b82e18e693e6b85b2f28d4dedf256a70ea37881f4eab189e99bc737289;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eaa9da63b3e24ab179b03303ec444a3105b6101c61ccd3856f074c120fac2269986389be94c521a7ba7c2114b3111580620f8323a94df9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1319b879665915720ab5c2c5f0a0236d77f75f9551f84657c01834cba6cb96e54d8acc69f43e556209922bbf238f927fab196290b858dd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156db618222295ce6f68d39087ff22a5484671c3c05a96e22337e7973cf83dd41ad58db5ec3fba12da9cc8cca9d8d07dae706a38eae8508;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10cb2ce549c84036a890386401acf832da6cd91bddacfd3bfd259102fe1f2de8cf3bc067d0ebf97beda9c3f2a6b50454025c423c48a4459;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80ccfa53a1a0869e3cbf753bffeb0634f8cc8508a720987c420d43eb7258d5c60cda951bfe157da4bb39933d0925af61dc25df0b5e1fac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4fcb5031fffbcecfa5184853ffa9b1159742e87fa150057bdaff680209e21aee15f8d79660e47a2da8984b7c0ce4bccf135e758dde560;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152ce0a86ca9f39047ae12efa65325fbe4c6943bd0363bbef64a0efe1dd08bacc4512a011f8cc91310b1462897087304c69780e1399731c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1632c973af1eddb443ff00e2e92e4fdadf74588a09806786ba60093cc5cee50d29c68c653d1378105b7f1ace47b5adabf652e7dffbe43db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91df5da47987d8d15721ea63c276c968dc941125447a364a08b0ce0c2901e3846bbc62dd3105e1e30a62600aef56934b0ee70447bd4f4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c85d26e5bcecdb4ec2d145fdf8a4be970afcbb79cc673dc3f3a1851721c9b444d142d7e565f91985faf8b5d80a83737d426e4ffd71917;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b79a3c3d2c841bc99cc5193f4e681b9ffd45c624952cb9c4cdeda920d4b48fa8f67f770c5bf86e05298dca92eab6fc4f4f79690c9ac58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ae6e7ca23febdc79aff6e41e33f65e9aa0389323606c3079d47a880d745917e149048fba063d6001182cf98a0c0c5a95f543972941dd3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147629dd6e2a648cd469feca3cfa6dc82ab8968861d8f56ebd0dc3c9edf838c29423aef9b167edb893052fcfcb6b4be952846d41ade147a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h329ffa19579898a35b56ce14b39773863b783bf8c49ca1d04b3afd1232bdafeaacf2073ad66cf6700b22431c0485fa64fdcd1cc0e910c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a5dfaa6ddad2e3dbd172057cf241e688d8e41c9b3a47b2e686da0d648c163c4e11028ee0a7fbe4b9c5d383134f795ab7f9dd81bfdb8b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc9274f66661ae46e34757fb12271a692ef58edbe8ac8ee5bcf7eac3bfd9e43a203d423c5a0ec608f6d7c7eea47ba82e507757f7c47536;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf422a648ca8a26d854d310c70324b2cd182f1b8f65ee1c3266c5c5e1644a78b5eef4773b53e132c9d4f3ce0d67d94fdf5f5e5c799e6775;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce9a634d98c2f8a59030b63ee0a60401196ccd09f984a18255e47d29cbbc2e0c2b7b69fb8e8ce12cf64348a358d0c7c54b479a77e6548b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bdd02d652913b74e03520d2b3b387f9cbab80d0f502245db1de2dead32c3f9527c22f53e25b7267ef45df0a89a6594d95991573615748;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83fb48d4501bd1ea28b4c73e1a67465d71fa1579a6b1e337dff9ca28ed7b6c9ff7044cd277f3d1f4b830986e6d389b8a3043991cff7341;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc31731f9938ee95f95c8bc326fb13cb8e564a908b4177c192be5ddb27a88dc8f64f81d40fa6dcc67296530d76ebddaa7f3b36f65eef19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab7fff4e18e91dbcb3b2095bef6e0cad5d783215c910c4ebbeccf800ae0d35d776bf8683fc6d12d4c0de49522380e1d0bf0593e6d79731;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae9b5f7184431e428930b56a2184d9f2774fd6dd77f0ffeb56de8875c75b5159fe9f84bda922e03a7c92b7c835d74df6fab817bdff5a08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf02de82db9ebecb560424a720a3a926271c94c7b038fce65f7d7c0681b69d1169b58d2c1e70f35192bd5e57515e12f9323767578c49e1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9dde5e04d091cde298ddce6b2214e676b0dc8bd8ea670950941cddeecf73a4a7c3f2be2de0f69ced75772889d6ef4202034a128577b951;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8d7bd6dbd6d7a7b28e6ab7c33f133798c8d2f6fd4b6e5bb8c0989e6d2fb3b954a04fb70a8b9f95bad35b2d8e77fe36c3c1ee014aa499b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc458138beebf49aa1bacd0a62a0a31630a38ba11db3a782520beebadbd5f83b5925c37c8dc396339253a70af666d45250f1cb53a9c5d45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1869faf2665a49c406b11572b3c3984af1d782b0e87f42240161af7e3349d186901fdd49be301160270b0b3814f4ff03aa68d58ac0eb459;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f566ee49f08683dce7e7fdc3f768cd9abcae86e93a4c13664eda94521e63d7b883003a13bdc602d90664b1e844339f688510444a3807a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd4b3dd1156d90aeb7b63ea957a0630d424021dbb2575d6321c44f8a3127b648e31192430c6c147f54a3a33fb2eb7ff75965ed92813322;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188398b6973353c994dffabc133015bba1f3901d5103a4c133994be5a3ae130d563845e9484592370e0207d0c365790f7063918439168e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bacb67ec2c8ad3aa8a0a8a47defdec329181e1e046b71c8ce6de4b25f3b53e1bf2f07862e3a9caad4a2df6b5614fef8f430b2b8e7e24f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c98e52ff5f4af5702ef4bfaf17ae6ffaf56eb71477cbe5a6436317d504d6ac2b0c12d1f18ca74a5a92ce855c6850f954b8bb15b49cdeb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h796153bfff2141bdf0c50e9a2932e376b0ebf5318337a7fc5bb53c8f8a158183472f7d97a259eb529705ef8bb3be8a5c62f42205cc0738;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15768c4565d12501737d9ceb04e82f98c460e0dedfd516c4eff915d2975d802cdbde8acddffdc0ff7292e89222b07ee237e42bbb6d0deea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heceee1571529d2673f25e887bfef04c94b1e0438652bbb4827f86ac973803234d2ffdc21e8c3208fa2611ba48070f4dfe385691ab8b42c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bbf0b196306eff6d2890de09ef13a93826e3d13e6010be31eb3d3e43bdd439365821c3acc0654aec1ae7f39fe51ea486c2b91653a5c41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af14f72d6083d959fb5c8b234e9fba4aed2be8a7d6275d0470c204988abe8ccefbd05502cc31042e66ceaf23b149cce08f452ea5d3ffea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f6747b803cdf5c3159812f2f43a6c8f37f1fc169c18079c9c04abeab696ad3faecb0597a3adda837bc3fb14563872c6afa357bfe2c72e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71e5f109b84e853d9de5c1c4760290d399596dfb37d1d244de737fe9ed7889e96c8e4fe8f6ae8e07fdf70a2307489eec4f51c6fc7c04e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdbc1901af325e60d765f122f2a57368cb36e19395fb85530799775d72578c30ce50792313f734781764d3481a5e8c28f0ee7d6878a4d9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55c782ce15b4a0c7dc953d587f09316bd8218a1b82ed019690e7b9a383aa90c676876a69511ff3c28da3f541b06f7f2342c10627fc77c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e66c5041831eff6aab71fc2d22977677dacbbc5ddf9c23d1cd32bf6ea11621eed2c95b6dafe326ec5f98b7003b5e43b6b5d10e81f66e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee39ed0400b60369ce58ec29660b9a4f43ac25995dc062075e58221e1ef04f564bd79302c5ced0276f298a0910e30d23b154a00daeea07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h409b62be18a6f69ebff6a18ea197223571578636082fc62982df67c6b4731c62837af127586a5223a13fa3e01612c50ca0f70a65a47574;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c08cc8e36a8706f5dd467cdf750715ef63e75668c4cf0e944f8c19ecc919a33e036267e1373844dd63a8de4f97c35e3c9ccda897883c1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44e36fab0ad7218f67edeea422ea52b9323a999a904ce3f77f202a11b84104428b4cfe6a05db19ef399e4498ee9eabcc35bdcdf4530b09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heda4b1177fb1516bc61270772dee76f188a1e8848499fdb1b8e2889ef5cdac9442e545e0f36f852c1e0647b149230a91d2609ac3aebc2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62715b9ba56df88efd6eb5f48d7dbaeba890a46a43fc4c9b1a2acca5b2dbe9c31a46a26819cc8a191c344ebf22106b60a48220647d18df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53f0c962f70e30e6bf48fec7709e355418999411b51b18d702efa59f49354cfa90b36ece7bfc237ff11a6f15d8c1586c2d66796dcda0b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ba492738332e8d5373025189f15b891b8998d8db38ac06b804037bd65f1e4aec2f7848dcf2b58b60bd47da1b1eef3015d4779a8656da0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1610581cf65c0798012108760ac0476d924aa9fe0b4af71b486bcb0045f014191575a4e1b168d8ceeefb0d83f710b85d2dfb75486c52e77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b99be10132122e059c86e23af67ed93bcff59534761f132bb13bba0151ebadc3a54b1564390be2ecb42c6eff5ef311d9feca96264926f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ea2a76b40ca4f1f19b52c561091c834f7234e0a77f8c23e944164770524ed86269f132d9ce5d00529e2159a06557ca20febc7fd817ea1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73353d8434192f568e74dc8a48f13949da5f5ab59a0c50db0bf205ba713b6c6c25bb796f0acdcc3b02be4b84bd56d8e5abba1b6ed77e04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d6b9602904a2853c4b4632ffa8252f1a91b81b023889da2848f136140da63f6941c34f6c5bd300fc5d5c113b7d7f1d608a036a5e0adf8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63ff6db3e53f4d2ede9c227e48f279d8e76eaa55185358a31493f5bae2f1dc0ec535676e3414198a096790a91d28ea9260cbde6b76af3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a6d305d2ae66faf9c375152585ca05c203d3758390acc283bb706e35d3cf1489b783e952b27a25da5c35d48886076aa3c23fc94e6eb70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0078dcbef5cac687bdbf9a1882e00a18b0c4397d3ff471943f5c07c6b99ba8e8e7f4d92886519c67018c4c33fafee33b0ed25a074f1ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb9c080c6d5f16abc1a704e981f252a6fa714df5c5246a7b7488b1f2d4a8e8585516849826742f6d9c880324299dd78af3a5b0faf7ca8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h244fbf038d907f9732ce0b3cfd02f92c643dae822d0d0b74cef43b4eb7e7de0d20c6432f1c609b523b8a811aa6e502478f33e7b17b105c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11dd4330455df0663d5397024ac77e85ddcfec2eca0f0d78b3c23413ad6c71cf34e473b16686a2319da80e9cedf59ffc2a892b6ea9d8baa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c9bb405aba62374a794b4b3056575b6fa2f12ec0dad4cc7a889464b6cd0406411175ad31a8e83be2e24aad7f3622ac6b8f69886547699;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc120dde99544814665b455bfa29692d53b30fb74098411419b9e48eab37b30d62a802021182f39affcb74cca2df665ed0fd7e6adde7a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34ee4442db29ae5b72f1303a2a0625d94d65f531f51beb565f6d2e807014da7ddbd7409b4352478d1b487b4e4b6eec9ba0e962c35bd6fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd81a620477ff56908a09c4ebe96e9f89e5f7b4f4f0e1eeca3471687e6405ec333a5f9e9756ff7859dd64a317a7917aaf2e883c915a3ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb7852aae1309c45acaacb6d8c51319635ee53c4050cd2df26ba8fb95718ec6f23646e5b5a97802d214da9542588377594514c9d8c0a94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14749910de3d1a89830f3c28b60aa9bcb3bad0c6c558de975245361740eb1b91ec0a3687398e617a21c05aa3b33660179f64a6a00fb9b3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1133b2d83484c4f758af5989e633ec06dcb059ca4f59ddb57b51a1b77a04427292207815485f9ccf54cf2943ab4f5dca497f62d76da2e9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e031347e27d372a836508a59cec69941abdeef0d926508071adc13f0b02b827669ca02aeab399412c33291609ba043f1688889751464c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9f423745141e67d7b723b841a6b9985cd43dd49931901cf00b82e0bacbf883e46a7e02f83c4da2bd6f59d9c9020b85652ccd8d2188106;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d89f27f0b2b43d91ec26fce8e11a60b94d458fb206a4bd9066cc4242311363b7784ef804a4bf67ce114cbcc0b97d1dc957bac4eb0b9f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b264865935be4758bb5b4d2e3c90a76bb815a1a5761d8f2e1289cbd3330ef5a2d2e368ef355b864acaab817030a680a393437aef1b33d3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bfbe38f8a608cc0dd32f516a2959b9f02c43fb053d465b47388562ad7b042721c92099fb3e1d39e9e02831c409f2932bd54913299f331;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18577fbd32fc97091a7b3247c2d810d0c558b7257f45d2b3778f5a25591973babf1760a11b8ae42e7feb004ca48ca2102e3b13258d07f26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80bc4d8e29dc0e10d413de5ed6c0bd1abeebb2a2cfb267de792717989dfa79ae0a97f1b18a772d0e14ac7254dbb65c35a1626e1a103ea8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65caece45562c2df9c4c2b78a789298e37909a674211d1e3082753121d67b87164219ca979b7b49d0b8d3ba3f5cc9559817d29a4dfddcf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178395f4ce9a706843082804729f35375bfbdc09c1aa0f9cf25219df307654b38ea421f698d1077d063d312d39cb377169617a1e405671a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ffb242c965e23196805c7feced2a8bad5ef5d01a2b9a2ec9b490d0e9132c2e548111d4cca09dd403f42203211def17946554750499170;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h72b7364dd40dbeedd327fa67df64c83cb6ac07db19906646e10d24e39938832ed14f5bff310314aa3b790f91ac1d5044d9dbc6c695b0e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b011455f000ea3ab9d8e50c26eea53e41ae0db94f03def397331c669ceda785196889dc6b77d06fdd426a4801ae5c14e4735ee1b6a8768;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ae289df5d862dc7774b03b51b4aa0b006acfda644332c85c8b0617e7e5a92b14639f360150782ca75913d473745e78b638abfb7ca13d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8977214e11ffa63e462b7a4a970dc3a7c0878550b930a1acfe033e4092963d6984d63fd111cb6bc8ff562b05860c6463467126026a1bd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b134e6b2f47092e90fc3ffc3fbf879f5bcad74ebe04899b50bf705e6dbd796b2fb7a54b9dd9e299fde036871aff8422494bc81387d861;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca3e20875045cfbb4c93358ae6d3ef759e474d9d228a8fac06286ac3aa0ea9d416db8d70b262ca2a6e2dab5adb9aca222454ccb4d6d3ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a76351c12d0059ad18d725bc9aaeb4d3fac85050930c0fce65550281aead3b3ed8b021464bf2fc6e9f6796feba4110db719bcb4a495dda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b743b62a7cf98bd8017cc57bda75ba0793a67890e9cb93eee2b7c9b8fc76e0febfffb7882ac7fae553cb62373bb2c0ce34940f32df9f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1735b2ff14c5d17cc556a5ab3b8a0082601862a7afc94f1d2d93b7e39ddf4c8976b86039b0be5e38bdbb4bf28f49af24d2a501e254069;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ede429f6a1de43e3cd520fae364efb8272623ec5012c017c9a059240ac472b92a7a01170af0273de1561f8bb84ffd50c4c561951df328;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7e3f1ed1eb145e88d2677b0da5401ffc92970ca24d961bd07c70695f54f9813fe32555baa7b5982c608e96476027fb10ecc3c619899a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb055078a2c904c7959fa6ab3e70edcb15f55c20d73c1370d822b88fecff05396ceb440b78f66774ca03e683ef4f827bfa315d7ab5b7783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9389814647ba5444b7863d3deb9d7a2428e80ab70d57d76f5f2bbeccacd153daf8d6c458c46f54dd78afea030c7205e60d0a446f83a244;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124f64836900c03bfa0510506bb7f1b22ff57c99675bbcdbbb74923252614719815180e9b4507db35ddce9596807d5a74de14bb16b08578;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73915fb51c7e27cf85f7f074f7ec5a3bb6799693d4554b67ba29fceddac6c4db2d114948c138791e28fd4ecceefea8259a934f2d3ef441;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cc60b2d4b88e81f841916c20491ff55f2fba8455eb9951fafe2352df531029d1a1af99cfa5e29061f9c77fdc6b691bcc3250d4e14e53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a692a940d4264ee9ce4315637de40d61ffa56efe56309493a40c212ab0063bb557906921681e25cc870bb28ef37e0c091f8c5831720933;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16931cba4082f37f7cac55de81844e19061a3f3b68ab4c2f0e88996f0f1696c3ca2fb6829425a934b48222d098c9404953a93d52a59e82a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a1c6b1aecdfe1dd06d8a3686d6c5ed0d60ab5ea774595086cdbadd0664f7118054751c47255cb0864a0f23a75d0e68b49124af1356f3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34527dd40505fff41a9ffeae5894eb861baa0bf0fb63481e18f1edf9abaf82c6d3a0b1db2dc18223f033bdbbc1b046158a85f8b73f1081;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde7a43f8ff87b8627e6002658e0e8367650df4228a6aa5e238d2668016015eeda558e98e7509a04ea15d2ef19181d37bf4bcda53fd87c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha51e42127a6a730cf3317e3107f278c28b48c74fbc33725b8e8c44d49ad40b10df68e845531e759bb6205f253b9b8967e017390805f35c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f7885900dd4b7fcbcd17ea80ef1b44dfda57b1f583c23dd530934dc06946254d64fd39d79bd59dd89e5e9e5eb8621fe7a1091af72a61f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1897d4669027783a8128ab7bbf22160e997ec7394a3526de2a3567214e20e275ea86b9ce9f3b5ace572a351f10fecd2de704d62ee38ef79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79042d67ac0287297d94530458f68cdbd5a5694fdaa14f4c1398cfb4525573ba97c61abdeabaf52324dd33abba55bb3e1da9c62e30feca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1736a97459e940a9c23ec1b40e111ba836bcf6350df223e3801a4c789c7e6255cddb7e63e334ae609430904309b0c61deeb6d76f88237f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e9b8b2259f1dff896d04794cf1578e81d34f312f534b31e75b578537922a40d28cc8e200c77a5c3be3aed2f2b5201c3502f4cd53fd788;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ac5550765ce71652a61828a31e5c7cd84f5c95158628cc9185c0ade0cdddade013585b591461d52180e489c48e5ac22c60ac58ab16c9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ca607eb37d88ea8dbf40d9dbb98adef6d7d4f73add73bf31cf02e2db7ee737967d035c41f2bb882fa0d6f8afde4573965475ba369f581;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a7df8761ad65c09d5d9ecc3bd7bb054104d6f5d71332428a0c1466cc12bcc5667a5ae69e6f9cbef97ae4b235bb0f6edb8110fb408d250;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b114ebbe12aed84ee1d6ee859b4c9f6ee8c46533d44725cd4ff69075e9e5062c3c900b79f90a2fcf8c2cf57441953b531534a7d811d03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91876f4cc1bdb644c41e58d59991d75e224117ffd1f229488e1323eb951997c879d9c967617d32a8b70b78bb5edd5166c58154214aa453;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d591d3d8d726d74fb3be4e8a2e7ea83e56cb34918a17bf2087ce01e815f16509e1a095af186517ec79be88f9b43895332a1819c117ad9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192a408a6bfb626f2520873570d2192fd0a031f8737d0a5ca393f3baa0071c36cfac874009894e3820ce433cc705a7299c25b77a364ea5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8fd846789bdf7f883c8f4e032648177bb729620aebe449e239e62296f73926a351ff46b7eb6bfa4aff0797d463a35a14a40c4adf4f2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfe6f72c968c9e5ef0f7d2bc1ac03be4b5eeed554e26b2c2d024534be68bf440f9d57c42b649c48531328b957b1530ed0d1afb5ffabe29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5bdf6bd4ce2f2d273fbe0af6aa6c7ed2174e954e6ae0044b421c18827939f87e12b7b694ab2cab06d2ae2621fbe159d74e3ebf7d29724;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109a4b1351e40d554b5416190b5f3d0c19a96bfe5b84135c0b4214c060ea69adfdf1f58026f3411c4abe06caf2ab58ae1b71dcb3c6082e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b714ce74f2268428f4dff1bda08cd10aa1b02baf80e29ca0255dfecc0bb22706489662ac9aca012b730ef2d0cde4dd712b61690cf8a534;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180864ff114711a68c5d68a902e786e2d4bef4466a1482ae75f5242cc131c89f9d2a654afdf1f86018a27a6872842d7195c625223950eb2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14266c2efd2ac33306d0bd1218cc337505376a1edae62bd839ec4eb275a1361b3880cd61fe6ce6864d4b4086197e4915dfdb480caa9e9c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2c65cb2f4df65df97db02bb6efe14b1e0d5c4fd3ce767febf5c950f8647740b17b271e09fdf9d945ae12137d12fbe1d9a781fd5e6a1bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d260ff75e19f502f81f40d4e39fbfe89a7e8df923e6d89791ab220e1edc416cd5675f9b86cdab964e3320ba3d2b553bb3d0265fb1dc73f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16932ab9065525daf7002c07295e9b693bc1d3aaa238ca44caffc021141d787e149ddf74dd866cf1d5bde6cc85b1e41c875362839f821d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179b9953e40cc39902b533b543bfba423945ee34049c18f06848cc17bc6582827451e42ff317b47869597d266d9b054426e57a0b474420e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1747294f68c6fd2ebebb04338518389eecd9a1e154f91b0bb661ae25fa3ad705a99250ec062870f96f2fb5b495493cba31fa6b54783b386;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e59112201d2ae992021af47ce461e427f0e6ff4d964ee96157fc32c503046a433839c840d98762ddf3727e5147b8312e0130264ed5440;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dba182fcc6f5cd0e63ebcf7bec20a3cd1f42d0735dd7a249a50cd373b6c03cac835634d43725da2e9d75de33079864b3925c16db1d461d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d188e2ac477dd08f0ce333d19bb97b41fb5eb6b28a89fb7fb9af6ea0124c5f418c1bbe0d55bfa60e05fd3bff8ef2a31dfc746620e2187;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18300d70fc6b41fd8ed42fcace8eef49daf1b68cea94465051fd3f3256012aab2d1fddc862aeedf1c27367a16289be6da85abde887b66da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae737405431cc445b858323245b8f7f197ef4cb2d11276e4ef1e99174e9e9d3b27a6621bd30f8a8effb27aa5beb16ec61ef93ac85f6440;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcf05a2597c9882d4e63afaaf15d544be150b54e31475f0ed8352b77521b781e97975696e302461b1274cda5ab4fb04b2790b85528858f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8c24d0fbf79579805dd30b8895cd6880c0cd695d0ee53bdfa225609ff5ad3162e0ea7a3e00a9069134593e682fa6e0dd1504505d47d60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19613eccc7414d31443f0cb088d54f3298c055ee926289c6ae98346fa3d443dc00e18164c9764629d8c247a24d67b7e0fdfa67b15024062;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10beb00af2512e265b504e5b895562c460318973a4435d29cbf5243f252a037ab32b89e1547759819c01c66c6c061fd87c6b73cfea8818c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc290b8ce1a4235141816be13a92cb1670dd2c1739f65a529447dd36a0e9ba66381efdfca631fdebe1bc28e6d57f4442db311d2d4158bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66298140f75c9afd6f008d57fbbd3233a15565ce086f21bc0664a9a26e7cee996f406845f48926c8a40cddc31d73390fd43ea01a2fd372;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1244dea4622d99f36ec73c6d76b2236caef54d622ab819377ac8a0c21a3bea652f77994a8fcc9063e49802bd1f328295c643e87fe3e5376;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b42ee0d7c7f804c85f7d2faede9f5bd82181bcadf431b01e28ed8bdc536b99d2ff964e23411a6c0e135c34c4a8f55d909649cc59e4bc69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9e741a7e629eb4ae7c3618255126fb1aeed82409ac4fd471f5d9e31102bd4c9eb77968950f87bbdd7d395635cc53af2ac4d1b28c59fd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1643b3c8ddf1e8f55fecc6c861fee374f4632d8bce32dc124ab2fd119019fa93650073abf96e245af49e05c9f282c4cea95b8805f4b04be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173b109108cfedc3176e7bff503f49f6a036ecfbb9e064c2d81d8c172cc720d18ebb9136a542dd2227b6e67357751de0be05ead688ec6e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138ed64fff07c31b4e8d31cc2ae48b18ec70efc1e9c2ec90b171c9ec7a0983b2aa88e9e27c490fb45dcafc084738585a26dece2df396989;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7cdf3f05cb7e9d8210efb7953b8afe26041359688ca3117a7cb87fb331c62dfa0da9a2af1e75ca8b1fb4d9f196b4e6d512f346a90ee8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac20cf711d4f528f0ac1ef15416165655a46ec48c16c4a2f12199ede32d411d875325be7ed9d0e63c3316eaceb0f14bdd2e09bb18b64c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c557af5879183775edbd49e7b5c0a356d2dde03b8e101bee6d40bad1b0da7f5cc1999499aa5fe34fe49e6881df55952f3e1d4962ce0f26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee281b9f6692d69eb70748f5b0be473bcb1b1c0668ce97da9d50e9e4c1abbc0cc179ac825cc4327738baa80e38f1e9778b5c013ee1d015;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had24516fc1d28e822aa60dcf40a8806106a138730c64570ea9e8ff974e5699bc11f0d6352cdc9ad9e6266d813df0b8e2e17d480e69cd82;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h592625a78d1e9942c9d641a7d79e30881a43e8aaa73b3da7e246b5d4a6173b636058b6e7da5017a804a2369537b1fed5ab3269e394cf66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1efc801ff5d7281869725f391176ae51b2277f41d6c193578033090c856edda2a17955fd9de3515e8b2373dc93cd98c6453c8e53deb5aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54c1fef3640e8b62db8f0eac3a2aad663e05094f63a319509219ff1279f0a146217aeefac1936b58f4d24cdf72a3175fc0a5ce50de46f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1747b71f7d37acc1d858ac7a542ced79356691fece5f79639dedb9f6e6e2d144b8200a64fa1f28eed5ce04ebd5d9af6b95b60cd5bd80503;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1553bf0ebe6892d902726126e38a8322fd9a6bba101aa1362b80f82b84a60bb4b9f036024d134bd5d3be2088dd5cf18d68df03c8b14e19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71cf502bc886c33e071cf1fd7c7673c4de66956825a54d762e372d4a109c15399430b1c98f124a9e81b3cf3f8683560235e9a81a1d2020;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8c0544d969b561c1160badae46d6907ed7b54d167584d097db99f73a874078f44627a94c5f1196c9f840c953cea2e88724e09b0c04241;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba5315f551defca450879051058c0f81f7f771341c0a74dee3f7804bbffa7b977cd30b50c16857966998385898627346ffc4eb61d6fa45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bc3e3f17ffb1613a8802434954503b7efff42270687191196c203a8b88d21cc525af82663dc9e4e9c61628769e1624a127a79e0afafd8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8da8ba4240f255cfd971fbd0eb5b0cec102a41c9b4a8334fc1233d999bc6f45e0f2bd3d5002ecfa1d901678e8caeab77bfe4e9537fa0cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17737239e8d874ef9f9f23666bb4ac9bcb4078584fe060cfc06943ce6e4a252f400c51c398c7a6aabe39b783668c0bb02c4f2948c572d54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef7259a8f6d53b39362161fbb8cf06698522744e8456a9dadbcd50e0a774bd93512520be56be1e2f0b756d6c9dbcdfce7b931236776e16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbb8170c46760382d3c4d8ed3b48fc867ee5db645961a67308f4094fda0fd1b60706b02b508ea3a365b2f63d10c7a27b533aa265297427;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb20b8ffa176cac44c94a882ddbefce131a3109e547b1c45b8454f31e3c29446af9e8bbe8a9811607ddc406d23bc2347dc5e88fd1e7622;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb50546ff1adab743133bc708f12b170b0b765a7a94c4fc517b1f08eadaa26a240939274bb290bff94929acdd4b0ebb52a720f7a8fa97f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fdb65cb2994e53dd98f31131978d306aeb3f6abd77adea4234d5379d1b57c3dd4a721b20e8fa6ecaa450d0e8ead2b33aafa47ddf97eb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5f2b6d8efa3fc4c1cdf8cfea1a2e2fe97112e16941bbea845a0d4aa381e12206b64d51f3c4f429b873b301ecb02fc1add4e4f79a7f517;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3096ac9785eee10edd94d9e5926a12507d7f17c1700e00124595f5d0a5f00e36a58e4f2569063d48d9bc7fc81275fdd8568672f8c58d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b04284d556647682cf1584126e19c4b4dcbfd8464d8dc15353250eba5db8a6a24c76c5576bc01884139f5b91b80d55efc842e9e52eb45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f36f433130536151d3506cb0e91cb28211c918fb53cb1d6c527c6f61f55b9a085af1b7e7a994ae821eb1f609c879b8f7761154c621bc03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d2a08654f6ef19c0b173bd5cd088928b40258b03d9527e418b5b475bb56b432bc12fb100009fc67904929e5d300cd7be772a1f0a058ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c209fb51b04aae14264068e97f66409ff579a5e4776f7e8e4360b5cba753af61a4b394f917ea6266652ab0f706677b263598ca4c6127fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d394540e62951ec824660c53ba241f20a17e86b07ae71b092cd3b14d160bccb1f6a155d3abbaccfe8391e92a1d745e0f27a8f7936d5854;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a925b5c8674d76324047b34878c5c9da1cbefe42286bf26db52842551f0091d375e8d7201e045c2034fbcf4f768772d1f41d2a701df5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162907aaae153ec1bded2956886757a3d235ab66d0cefaad8cc68e8a0d3ad3f1c528acdd3c8197f00a1b3d418180f183235521f8684fedf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfb1045d47203bbe45c53f946f389ae382c91bf5fa0d27001a94270e1853cb06631a1ddc16e2f3d27ebddf7260f413eea9791919a3a569;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc125bb4703e076330521433d2bd2d7a0c3a709e1e456b45a1352510780b219b2bd6feda1d6d27402421bff6e497dfc465107aedc52c8d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b18b494403c305da52cccd05c0aa22c42386895fd74a4b6b6edab906c9b5a78cf492dff3662378804db146cd877ddc9aca8161fbe3186;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4482ad10b8bbd38e467b90e3069ca65179b907d392849d8eb4da5494c579aee21b94e0b38e1543f93f35cffcff6e5a7e0d3567087d1ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0177d3d6410076c1a53edf8c91415c0dceb7ed7d5d64a281bf9a78a752ac3e0ddccb593d5f945d03f0c25f4883146a27f330b4f336c63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1633e50e192ae34f28071903bf2144ddcc2d1685df3b4122a4664ea5442f30bdafa6b32333448de51a6b4bec6d19685249828bf54022ce5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce4750cd5467958f9ee1737defdf55974979c57d732afe84505261500df4a1b58de9b8c7f1c8cd1d8ce77e1b4e5c2ca5fb07878fc0f470;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2778ab0076a1e2381e3723ae9e110f56daca2c4e1458f13c0a15d32358c0d03e65199e21d5fc99b63ceff645e625e931cc8e0cfe80f4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h262ae88aaba2d296a9fa245026e9979932650187e8e842d070a03a0a3d2d48e41b1d56047cd3b550df2acd7f9febea6e82c6320c510a78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3368431e0ca9f6f2833e3ec3c50081b1fabdd3e85582bb4846e3fcad9f72b5414012bbf52e816512b7a54719d5225a43d6a44ec9ab30c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8c5b1d559bd92712cb67bf2ea0544135e6c0b4bed71878f62a4f0e712c9871999d6fb975c477cf560e515817672feddad1ac5c7140e17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a75d1a1342298debf965837628bd8d645da929b5fad5cbba9d8b0ed2dc9ec6110821438bbe34ebd2d5e0cb8002e12eb3db3a13cacbf97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14841e92e3d01104f707e7b0fa978b07e28494c65e9fce99f4c011fe6413191236cd9af3107dfb101e51de0a17bb05fbd0022d331f7892f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h203b76497cc499930ca3ce1d06dee0884297b4e8d0b003e82615df535bb6e6f9c66391ca44f064da016f9a3a2aaab9bdc3dbc28588a96f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fb7bc6c6748f16026ada316ee6277a4e59d1c0b5358137201655fbd2dcda2bfc273f9e921cac42214b3712852727692fbfc265427982c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1daa2184853060e11a60e1cf76d7ac7312b4c2803bd3ab33609a54df289f6ad21de1e815e013540dfc8d7475103bb638ce1dd7de3983bb2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8aa2d549dfdcf5128988351557a68daea9ee5ed06392402262712e13f45e747797b8383b6a628368bd297ce958aa37f3ba89b81538f522;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfad798379d5bb7a87e83cffce9a3e00f1f534274a6fdf818b6b5ea5b6f5e7b0c4b2581665ef54b2893feb0e2d8b33617c290566518666;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee0b3348c5bd89df664ddb6a8e40719cb3239472f28d9cbb4ac38000cda5acfccb8b2606d59414a7715d95d5d57705f85536c3e1aa61a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e88d9279a8ceb98ec8ba9eba5e9de9aee8dc7e15aa261c8c1d446775f8cc364556efc3d429aa5de7a19baa0f728f99c1042193597fe6e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192603a5ff4f31775d224839f8abc25c00e19aa88c44b54f3c7932d5535fd2629e5d1eaea1f16f69ed2b59243e8456da524ef83dccb8f04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a5762bf206486508908418a861739dbde133d5360fff27f19b19f9b43df304abc1287fff6cf7a473fd28955b4efca84bf8a9a4a88190e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146bfe5e8bccb6a443f4d86ffc038416835d7f03fa855e3f497d9c1505941c2f21a858d8af301d77c19c682eac1bec1b80031781c860666;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b6963df9fdd5c7e33f2b89c05d7ddbbd8d3219bcb49c5d85fa9e17fe1613cbb5e29109443782ac569241b75d9452880c2ef9206daa33d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbea2d0028d1e194a4cb3c17a429c7886d4436117ac5fcf7fc51e04748b40b3f0be4f23f31be087a08e70a1a2193d2cf0ce21a01db1cc2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111a62e7adfa0a7a2827381a519e1f85656ac6b8562cb6692959248cd87ea195c1b29da8c888881516a72445a3210b927d62588595bb22b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he293d0b323f3a970a6a7614f168c1754a9e92236c7e72ed5d687120006e5517f2f74e99dca60fbf8f95b680615ac0612020de40122d1ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5eb92893f0540cd7f94a98f698edee820664101727d40afd5358448dd5dfa84032131e16ef7f2044ae8e434208b8b0a56f0c4539f4cbe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ea5ca9ca5dbca13b28e339b83eb3d8b6b0f50f756dcc447a233d5ed48131adf7a9c4d83625a153c924811647501f5f9f6dd5dca9195b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6cc65e2bd05234e97e7512938b96868fc7977608723913eb07b6b7061ef79076a5a331c725753175ead111c691f787415dd48d106aa3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198f906039b5d96294bd5f9dde2f951e31115eec2cdc7e5367418fe6142b5ab3267510873519bbbec4d3c57a1b5d22dcf8fc2a2baeec045;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h721d79bd4acb35d767385aa9bbc88ba590e3ec8e970422c63f6e0acb28dcfb42002fd46ca003e9a5b29562dd850ad1f8a93f725c854f39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d4b35ccaf325444f98905e70ac986b53b0c1f0732155e900d63e10775f8159aa64b72c48889a21b0b44e82d7ec8550bb62b97a3910f2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b307b95dde1b81bb15c9fbdb3a080677031cfa75ad4878733f9bdd67ac7b0cd1257a6b7a34d8b12c4f671807b2c8f401dddd5efc15d495;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b483cc4245423b94aa387bea3af92a3e141f07d36e3aa278808486b74950b529fadf36aef40c25034e62a0889a00f1ba5ee20a1d875d7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac7ccbc57fe8fd208822b94491711fdb1e729c8e03c93c70c430c4b83413d73d3fe65c7a641626212bcbb55f5b1d91b4c2ba442c2031aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85376cec193daf163b18b4ae7caab1700b1a0242bb3d0981c9a58fdf70cbfbaca03e757d654b478a59f7e967453b485bdc0400d4832783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4182377c2998ab7b11352105b4ce680db675b0587ac592964f7433825bd4be4845cbbab89763a509c05b3100c5d82ee65a665b972e323e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1016b4119f9dd59c11f94c72fdea9cd391016b3cb291265b28a5daf4b7f566937943daf7427550c0eb064ad724444a0c8634d857c9a70f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1836ae15a7df3ff34f9775ba9be281cad98d60895e574d9a051a5ed851e53d9683851ea8a9373a00aa7d6ca6a5eae41ced7e866baa2e03d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55e128a34b1bf720a2bbcb4cc1a297fd45c68e4f7d02824edee69bfe65d948d7025babe0f29fe93373df8ace34af03a9d8ca6fc851503a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108510c6cc8db16eb8c21697c7882520a9e5b8425c2abb664adf52d188a6de7198353da3401c01576bba71395509b83011d8472834430e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha99a910f838eb55e58dcc61c80da5d6af9eda764f1a94d764b5e2b8c5859140c9effb46b09817a768fd12904f698821bc70e47ec83eae3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa53ca0beda013c59a8c87f7c447576e0349d89e839ca2047fdcd98eea97749198b2aad77d63b6ac84308be2fd60c88b4e76f51d309986;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc105dbd0786b1957e704a84e8bfc74a13091013fb4e4215ac4b8bc2d8749ee0644ad226bf35f3c17cf6587e0d7268da2d8e337b4b6e36;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10420593a29213c7b1e0d16481e4815427cfe6eb57d970d6b835ad80ea5557f123e53e3ab8d19d08c3ef4c3a5209218aab72453794c98fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9c5241b6963bc57635e6bbba24f2c71de89ca5512c60bed04527e31c41b52080c1dbae2030a4484249ab99e670aa9608916125b184649;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f819843566234ac9d3a0964dab44ec53b0643bb4de0ef1313ea11f8557d277f414f7867d5063fc29eab00e58e0415e31ef5a7e8d93f87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed8ad9964b78e5a16850736dbcbb101b4387c1f0753eb9901950c016e049556fbab2640fb25910968d3ebe9c63314abb059e5f1f92e212;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e511449482e60a6b924acdabc3268252132df1e8d16f6647f1fd4fac3a9ea5c4ce429127e451bcd7f07423f28ba6961825c14ffeb81d65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12662055cdf0312314cee1eb202f520c491644b235ea28117f51ff5301ba7ce307c0424141ccb636df1a14b77de5d07dc6e8ff69676e986;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cda7cb06ca1b27a0f582af2571f280d4ed23b12d599470113ff98677bc5ed4a924cb7f3ac01b5e6822fa3fd254f2d441bdf5fcc67f44a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d240a95343d6c7bff5afa80c5623682350e5c5320d38cbae781946932d035ca3e4b458c8c09bdbeb8026541c3fec2f5bcb7f2435be0868;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hecfaa30f3cee55f19f5ebac16c40abf23ebf8f9f233235cac567adf5004be299ac4409cdd288ae845ec4e7c28cbb61b79eab839f47e7c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159f641c56c7c8e1262a4bab069814337adbb1c22120bb137d983f483676e78179310a46f8be3164be57e6a2ae779be329b9240489a57ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2eb61ca9444d9ef5d02adcc035ebe97f9851765b675655e0ef1c1cce708d0b02a4b724cbbc2bc4393c397aefb329c223cf8f1cd438d321;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1452fb522ba74bfd4ad447f58fd86885c0ccf65281baf22d37fbc985df2a909907633ca7ac50ca717ccfc878bf69fcb01631cbb0dcb21ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6993c904b610ed7ee1d534889a9112bf1820b7018d439ec4d4bdcc0e7462e82d1b758593c8343ffb4079db33c344c97753b078400378;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a69722e024230dbf50848ffef0b988e521a634378a77d175e9828612acd4fc4edf16737497cf174fd3dae7c6911b8b893ce998f89b11b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0147207d377619a288b84b0a224c521dd427aa5373e453f8264e2b9588ac7e50d3dbce6d13d6ae02f3299493ac8900da5a276ad1b2424;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h661a1e7c54e9963e88650dc90601277e213c0ff5183a792028cc9f06803479ab09b0b1dd437a4fd58cb172df18b283bbd844672e2feeae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91336ff8ef8e78dd3dd06732e306cd66fdaef9c0713d31066c2a76f1c17fa8abaa94b4c40a6424b5f845e4ba10c8ad3d0182c66a4ff7c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbaf2585061d15e1edaae818a49304dbeade4ae9014b06dab90ab8d63d00ea1ebb604e06b6c5168bf2b5a73a72b27f053da247affb97944;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f084a5a03c5b7b7994031f39c53ae9eea5936ae8e9449071ae7cc357453b9fd18ad99ae2ba166033739bdedeebf3c3089e26647f2ee43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1230882e65361f6b41476c71ed60d07fffce3b8895eab23cd0bdbb95194884a4c2290acbb9f2c3368160a7a30951050d768d9f40dc9da34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11632230012c3fcc76047646422f09292ad783ab68175f39c6f54dd6f52b4a4bc169c0b01e738c00650ceab8b639acdd00698c66d22244b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110a33421396677b10cacd08ac51e1241278bc9a489b2a3c3a247e59c68d0ea6f254a1bd957e4ca3ff31760b2300757c7bd5f8aea2858ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dc79f5a6dde22982ffc5bcecd5c13178ef1faf8250592d72a4775c250a98cec722778310271fae3f1c60686953bc9c702ced47234e7b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c290630b0729b9019d9c81f1c3b292e0fa5feadd54a14cbf65203f2e3d3d8a2aeb84be521489e76a9352efef4fa5645419a19b68405ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h679ef75ef49f27e7c8d550a1ff60362b723bbf9a8920604e3ec626a30aad57b91311bdcb51fa2b4dadf1d5f10fd5fafb3bba5cac4bc199;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17cf83eff7ad9c9631fddc1a876a196b3b47a66dac13acd2c365f8e6f897e35c84fbf5090e12c4bd79a076ac86fca2d2792097bf451b6ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1935ab84f52254578be213cbc808bdb03930ac9c6024abb1d26db7e6d971d741e92208b8d04c6d07396c0f6eed208a8da44adb2a39b3557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de622745cea8aac87c3b265ab0718ffd21cb0694476b78d2fa2c0940d724c954103211ae0e85a13f79f4b18b2ab95e9529a0a7862205bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae6afa957c650c9881ca5addeede22126515d02387f866e34ade8ef2d231535b007bcd3795a0f05c3b89af00e4d34afe6013243acd65fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e6c85ce7b9d55296e3b7117a791a201b250147455760b450b3e4086096ec5cda121896edf5c8d22d0d825bcb81f5dcb9ed1e7f14c4793;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1903d1e1dd87e0c6d8e755e65041a31a4582f2cb6b36d10bdc2ee587067ef76fc32b3771e5ac1777a80c1e17a1cf61a3bb7059dc58a72c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce45ddf7473343a4a67a14ee5da4e5597f7be39b7e73c9689c3cd177c7542c0d31b560db7511364a42c46b514d3c0e498077ae5d3645bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8dbd410dfd9a7e6a3ae1c21555c029452ba3d09b0479cdece5326db7756a22c832755ee36722eb21506e42dcbeaf8be42916286df26c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb397c36a23e1d2d97c412065f8a518752240336f5b50b16233a4858cb3726dfbefc05811398d69b957d0dc0392b9e7c3ffb126104b5be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89098d1756f3449604e1d37fc0ba96f84deadc52259bdd290ebda6da50b99ad42ce2ad3d33202bc7161df20dcef0f36a590591e3cfd864;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181fda377e5e37f7831c9ece1246db8976a2699fe98aa30c013448ec944b0188ade313e4529cdc6fc87dae31e1c1dc4f184c4f0f5782a98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e004090290fef5c0d759485225772151a00447aa26e2f06bb46cf2d44d60832f07371ba125b6daa0c22e665986681d8933957d06185bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f4864aef2a7a0c5c1ad28de2dbb5ee16bb499bfbf064cf2b89f226101245a3bf55dd44f139e8bcc788431270db129a3e621254e6e44ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h564e92c8faf1a86682ac4e6bf32ae00741f5e9c2ee7a65279201d393cb07956b6a94afb12345a1f0646d4ef5f973201c2c797d2d2182ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75875de66046b402ff1714fd2306453fcb28155943a7f45fd1f89126f145a43c39e5eed01d2221116621fa827b1d82958df8b5f27a7a62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3f9e7c436ed7b686f9f7d8b4c228c8e5c61fdf39d6d15f3bfc74e27a7d2d9ca37fbb62323c9de696961c0797a2a96fd6a1d11c1af19f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha41102116e7444c5b18a23ccc65d7283d815299c75c8e2b41fbf01aab1ec71ed99a834d67c4e131f4c7b0acdb1dddb16b4957f034d0166;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3cce0f8cb3baa94aa6e5fa5d2377a91a35ad0dae0ac7ff9f8aeb7bdc80582908bba26bdc6aae7069adfb3cb35549527b1076574f0631d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110e6b51ae6edd4b271a176bac8861700d1c4cb8456625e49bcca4196a68cccf0867f3f5460b298a15bb2db0d7d0ce62dc3b98eb10ae237;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1f27ea45a5f1d75209eb9ea94654e610d722bc5eb8997d3c053d316caa0e3a4f9b97a3a2258f1e8b8625bf8aabdcaf95aee05f31e52b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e492adf4db649bf124b0b89b31745cc44a9fa883106c62a7346e3b8a000cb0db4e2f5e9696c6c460b7e06cf31f180cd2c204959fcc5c16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h148abf2bd99ea900f672ae94f176f89f754a4baec98ff9cba8737e9098e30b5027ee967e3ca074c40a200bda6c1f07d70b410bd8478300c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5d02fae3d60c571747469d266b33f364e42c77de258310666e83c3adf740038aa0a6265fbd9de294804e0a72776ad7f90b5e9dbba8ead;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a71ad2b4559326c1acf3380e9fc297bcd62b78ec63f56c493012aea760c0c072b74211f76d3864a4585b5eef7f19d19e782c688a828c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1900c78f0815de6a83c71666ddb761a291b4c5f508b37910a7180fbfe4c8957f355db7041fd8ee010d9c0da24c7020577588817accee8ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb9c801dd7e57f73f73e78766c323538dc63b2e67c687e36487678b7a9229f75074fbb1502ef4815e54387b0110712a9a782d4c50b26ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heef9711ca3a1f8d97e4a210c90271260eef99162007a84be48987e8a1264e02fa772bddd275053abd5b4a6bd4284c87127eedb3bafd2ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7bfae7ec01289e262fee6647c0fd7380a08f8acdba90de7cc31022828c516a685c72b804b6b7e54c020681e2b212e5fe7665f0ae4e9ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17654d026d7c71c5d6d602b7d8f147222902f0b4fe6141659becc757b0248cc63a0c989dd0b86476df7847714cd5b950be511691dbe8a05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b66e924fbee676b71c6bc4501fb26e5871c8c603c0b1b2619fe85a0d99f9d6cac07358c812cc66dc4d86da500398c238b349781e8ba2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a613bc3bd45764417a3e3aa0a23ca5536d40344c8e72cd0ff8a3236c412934aff8771bfe74a5755ccc6ad02e5bd2858e46b9d61ecc015;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec4052e198dc48d694cbb49976628897f2cf0e1ec2b5481c4939cd18e3dcdda4ed00dfe1d903ec94fa0e44ff44a06d2d0e25528e68a688;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba7b5d79d07f455791f1ca6073fde6f95ce10e1b06712de42c33267ad4d4c52e819e01e2b4cf819147b153b178d964b856eeeef939b439;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b44409244c2f98602408c65128ed0f01425b436d8bb3a09268f77349c8a0f7c29e3757b724be830715273bee30643c92b146f4f3a4a15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h732d23874ca760f06f2d1fdacba6626a6119feb1428062605e72d647109ac142836de982e872bdaba799aaa1442a807353dc9fd1c7926;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1958621fd544ae9518f90b76240e879f98dbf95f8a81240d2036d84aef88ceb34f1ac0a55798681c171e9dfd64a0d3ed88c7284f3cc2c2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0f5b5c52e9d1aed0eddc52b05437c7375f75d31d4fa289fb19a1c74c2b766f7b10f014ad40e83d8461665dea6f78b4e19ffdbeac0b328;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc46ae2631cd34dc394304d3e008829539a0074c6044460e2db6da4a8cd9b420a93204ba7e8ae621807a5137732990b1eac64dd4b68477f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e12102e94dcf369017c62eefdbd5d96c88224a069671abed6ebff60d64c5e7409fb079d847e7d2f9d234b20ec736111b964b83349719c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6308b1b3709fb4a18a902096746e50901dc91ed58346769da41b8fab044baf2e0843f831328280f7e6b679d09d1d0a668c5134d8320f64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b4bf07cad6c64d28a448790b9d624d62e1a7afc3998d7b27dd4817e551d1cec8f9132d3b38a7bb6e17bcd36869f5629191a19d3b84c43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a18df211d26a382cb833fa96e06f6d4c7396acbc1573733eca669f512dc4b29e7133e1f7a3431a632835ac3a4370b37e7aad3b6fc52d9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e20425d1a44e25876aca893a014e6e51d2718891da889ef62387fa195f36b57aa7f146f84fc890ba5d136dd1c5391b651ce55155228a3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9710a4a9860f4e73419fe44e2bdc1defcb5f33990e189425525d3bdf768dc1c8a16fa47a9ce9f4d1a182526b1bac6f2af93dce1363b51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159b8fbfaa4f1d0016534804bdfa32f104469c285a474de5ee3df3e71f1bf3a5f1a3c60168fa509c142d4d307b28e7c00cb9a6f05df013a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b96badbcfdf50642344bb480e0ee100c1d2273f0568276ec25c967451f2c3a0e155699ff307e0d6b099276bc215af257cdf9bccc08154;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d17362b2b9198d5fd413b90404326455f55238bdc26adde5ca9ff35aa8939088a6d62fb843bd5bf0121632881e02848deab7c93e7c976;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9f522adfee30cbcf3fe9f00bdfcb030480a2c5b79c0fe2641cb0690d3753f7655f22702165465e0cbb5531596dcae4211fd77706fdb1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cc4840bc9f8f5c4be7a5bebb21e9ddd640aac31cca839da3b2bb8c2a51266c06b152c14397148be6ebd24987f5753b51b5fefa2c77d50;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef6c6d56fac1ce241b4421babe59fa3ff8b1ee281c6bea0b966c762156400bb2371d60be5bc44d3d5cf49934b6ac9b829152278f4dbf5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21949f0383e67db6c847b93d86f94b274be431088b58d0db9daaff6395615658a32d1616297577618577e08cbaf57c368ebd94380053d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8601502e3059adcc285777adf3b4294cf2947a13cabacdf21ae91fd13c34086f4d43522ab9fe49966f2282e5588a8f7a6cc544dc095a6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9c4655d5ee55e0e8a227dc42ae3bab1abca033913ae4b7cf0773c2daa3098f7473eb1c707177c88daf95e21c2f1cb8308870f5ce5e872;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4568225b02d7844ace664f0c4ac6a5f6391fec42462c77eb14fa2769933050b0a5b5fe8bbd655950414b5f6b6503545c88833773e7012;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a01749459b03f9e0c8fabcf3b64d27397454610d4998292eb6aed5a8416c3a07328811993f82114d28225934c1f0eaaa19a9d9c9068c4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e91bd6a949edab1f117e6fbdc52b80973d5b15fd2d159f7e7268bdd6abdf3fb73ef95fd7de3efaf1cc8b8afe8b2d95da587ecc49966b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cea44e281868c94323f44561aa640e0ea91e6921b1b0726ce330e84300343a291f77b3c82ed4fe8cce04f0dd1e8ca8bb2538a798b90af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0224f4ed962507198f085d94aa2a9c10e35de85bb8ebf91a12e6b20dc816b89c30a663312c322b6fdef502072fad8d8ed76757be15dd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1549acea80acaf53580eaaebcaa9a3748fb75a6705eca43c6f02595c7d4baa1f5556f89a706e86b1b01be12dc3cb5abdf6e72cace71523c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9dba71478dfa29db73969a87bf13f01586a9bcbffb348e7412d819a635cde5b06169b24e3578ab413747d421c61f5f9593e79a064afac6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0bed951424e76d0c05bc587ff7b9989ecf22cf59fdee696ae738c4cbcb2419661bdbcb87c89d1ac0db3c0d7f398dc064b1cd11079c09e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f74dcaffbd3622056cebcb7e081a4ad0620c9c55ded21722ec356aaa24ba4de39ab260acd608cc24e9b04878d3f8bcd2204e74a24af3d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96723013d5dcd98501434431b8fdfaf526f7765f1c2d3ded74f85f8a67939b0129cfed95da0717f54d4f7c1d01c00ed056d698fc888c27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6982b3be6cb8be3507b27dfc1b0f753b0e43104274ec50bf5eaa5c87e3b6cbec9e9a58febbb0c1f74c32c297d99a1e090a6d320b7c0d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde05e59dcea9744683cb5cc9d2a4d2d3e98523e5bff290d01a82baaaa26be9c98b51f053925c4c42b19ad7712a4c8ae17cfc9381d5c9c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd97d7031a5fe676fcf1c165e92a8e13ace80b2ec7cb5a50292c31a5bce004721b204beef92a27f453146f4ab72ee1dcdadb48731adfb2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0f24f682c52e83fedbd93bcda418f2d49ddb9f07a72cd037ec95a021d998396face5951e38a957fcc47c5a19717bef415877c9a87dfe8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c93a202e189c0bcf9a9661927a0108a85710269f4acb03740c57fd83d088e72303b108204116ce99bf8d947c116a1f580698bf9376d85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8d67226b830e67fd2f66848a60ae13b36badc71a3cf1e325bcb0a5d94f6b0d3234dc3ea06fcb59f23d58cc41c6343837f3e962e12a1c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17daa569e214ea27aebc06cee0a92605dd4310ff35112d39d6098e28f62f7fb6c7beeb1cec88ffd7683bd1c772e406e728dca730c66a37a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ccc31e81ade80edb22434f01c6b930427903d8b40bf39db863c100ad6f5eb1ee501b81fc83b78f21f2524d8b362d29c94eb91b3cf559;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7fa1f8faa0f9c21d0b9608a1075e47746a5f00feb277ae34a83a205cab8bec5a581c1dcb8a8052a36b581ae8714862980620041ed9d31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17adcab8067544000c03d3333cac3eb786313317839dbfdf944ac9d40528c56283d494dc418bb6dbb853a258053f2a18599ce9ee7bec16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d917afd4810747ae65abe32addec436356c11fc31d0a3560b2a92e458f6a65f1e985ce0b2e107d1d04d39dd81f55fb9a85297d5c0fd48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h558c3499b90e11be7f21f5aa8d05d6580c4acd5918298533161221e5b6444cd111a773807e85aef5ec14cb7562ec5e674e1ae4eba90ae3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f5d829ca5b046eb4d7fc38882620a4934b258b6f1db025b4ac511c71cecc3c09a09caf064b4d6783958f873e44c232bb598c64db2d8a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h148f6bd837e3bcdeba065e7f7daf2571627e438c7982e4faa0a2a2173eda1b31e547ea36bdaa69c8542358054b0193eed7fe7e38bdfe1a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde91540e5c89397a0b69825ab8b1d429cb73554fd0be41a03d475829cf798fc922d8893c57d571d6fb387a86385a154843d81f0f802464;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5245de88ffdb2cce29525a1327367190ce9baa9c4502d7fabace2d12f943b996a157a95a4f354cc3afd6aa1427cd5345054e7a2cce6a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90076b1cad4d4259958db4422319d51f652ca39e0f306d440ffa528edc001c7dac0aebb733146be943fc68f1f98aae74d35da8ec6571c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1983e80d696e0b4ec31e2bae70d644edc384fc619d3dc8c994abf966a75f91850e7f7031216bb0715a0b5f4dc657f3dbf9231955ba31dd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8634c9c5ed64ca64bc23ba87c5e2efddf1ea48e4c2b3b177390b874cf39e5ae149111465416e4b8665a17ccb4537d3c3ae62039e79d38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf649477a116250ebcffd00b22edae3e3e5d0c5d827f90bff9279b2f7f8cf0ca63ebbcb3f857ab1a8c8328e1dcdc749ffbc6f586e7fd04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b4dabad3c8c188884e93cbe3abbef58bb6de18a8e2aca79671f0e3857a1ec73852068e0cd599b704925265356b509f7cfb8e8aca816f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f67460265f61451eb316b2fb051ab4c3110a215e3d2bfea3f59b6e458a63f13e94676ce80e0e90b91503ebbdfef9a3bff5b21e0540b3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dee470321e4eecd04bb811792baf7dd1dc56874b18c4c9ed07a491a1c37203cacf66c6d5f41660789ecaa0bd2d288dc64896ba635d2b98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125245329ca241993544b9b4a09fcbc25488a02215216ec7e6f972fb229753c9bf1b0958590ddbb4d9662010ea12e7bd6cd6681ad06165e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af487c824f1ccfc400fcd971b24625e4ad5c6f20405e55d1b234af66521f121b591e35d154bad7ce7a49b95657bfd137cf41e4aa6ef1fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fa450c9d15283b0f8252db3930bd01395bbefe887c59bceb290a562f11d132b6ee0adca96959471f50a7f12a2290eea83cd20d4d6cf2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194ef84beedbcf732afd922c2b394e73e8befafe7999ef48fdecb242d0f788bcf6e6870c8dd5bd33c5ce0786ab39e4c19438183534b5bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1705658f7134a9977d17eeebb5efb82b861c66fecd2daffc2f980e492c6788b99e6991afd9bf0ebc6402d10fe235560e57e9608d53dded;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96ad63ae84d637aefa4d0c8e535ed28fd03f00c8aee2926e618d8261da173c6d87f1130e24850a3bf410afc7c161699661066e09ebd94d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h897a2ac4d37d70436712290344af72bde19bdac58f90d6dd65ba555b70b0d1979dfc087a28acbde101c12c35458dc0918ad8740ba077b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd000439d7da39f0ca77607c9eb796819e173d1c5c7a51213e6c0849319a1f9a03600c556eaed7f02b546df2d3d3a2a436193323bed968f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13dc9a08fb1672c29fefd94f14cfa879a484acfbfc41c6809b8e8718495124cc7e79dd1639d79b5980f808dfce0c389f5b37532ce682bd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1860ef73ecc54a4fdac4bb40f7760b8650ae391df3aff9217e900bcf30602f0a8da5e80619d9cb393768c08d4cf9295e08fa408d3575a23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd0e609a3e7d5719005799c9254ae21aba46f32bcaa73be2a392d6ccc84bb593a266d0690dbd9ac3df136eecef04270571c4efe8465517;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3abaf6ada0f3c3c9fa43152eeb4819e91c1a1c2b5121779e7d2ff93bd7f624f7d26c79da549f53de5ab78ce668d1b24de59a70abdc5cc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1941587a941329a44ae0bf2f273c472892bde8be9857193e74f6525ea14a4da67a0e75c5e0e930e8ee8245caaa45e8b95391c1c8ef406ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e7ba0173e718b3ecaad967c89790007e2ff525e82286d225bb6141e2991194a140972c297cba80ef119d9f52bfa32e5ed1d84c885cecd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9e5b233da9b1c12c2bafc2c4d02844354869399c4ae38392cc8fc99853e0a0c0d6bbe76edf48d30fbf73989f39d63a1328a26493efdd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde01df7c65e22b3e1df4b4689495f32b6d15b6872868b86a512afcec754775d223e8f51c8fddf679b299f104c64f4dcdf55483efca6b32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2711e23762df73b5deade36fcc2be402f71dbe730e91efff63e4495097bd995dfad8cc6fc49d535d59a3c28c8c9c2f2e0d7dec5590cf1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45ce2cc51b1a7a80d4dc321b3dc74e40b077e35e0a5a05dc821f68030f649ffa87594cb3df607a81e784bf898b0f2bfe2551b20e79edb5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0e0beee96017df2ecd702e1cd670d2160e45fb42b353e94df0369e1877eff811c20695d43fd35770c366083efc89f34e0835bbb098eab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e4af25f76189848165a5df598b145a143c717b68b58f5ebd84f4d0da1fe344bc475e94a59c811f27c7974d5bf7f8c555f69b1cfa1e3d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h493b79b9d930012cce3aaa37847c691179738c50f8cf99d324321fa72e6d20c47c58673d47bf5047806887bea4ffe022e1039bcde5dd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd3a1b8d2e16db68712be314471b4ebbe4b840a682cb69d9c43212ebcbaa3ae81e6a796a5d9d7bb1ef183c195a781b44c0f3eb89d6a479;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161d0eba57877b27ba3eb5abceadc2edc64b41e8c96f646da2ac34a0ef63f3440aa8a05fab42d8dd90d37eb4e270b1cafd5cc393f9d178a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4953f2afd886d80e0e773e27256f4ef31f6dc628a22aea97a08ec5308621d02165b00bc79a42ac2e0fa259bc3302c6ed9ed2181ab3298;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103e85141c5671275d26e0226f2fe042e72bcab912e31759e913d5f18b3b16f34c653837cc28e3a18624c362ebf0ec48e1689797b0c2cc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9268244df17da0255e12017f73a600e20b3072dd3acf226dc6f42733d8fd54878906e9d72202da8e1f82a4112e8c22b34674c68d3b9d16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3e1b22c35f51a24bbea9542de0131740a002a8ce15bb04598811f4dbaeba460fc68a1acea97e2ad26bac8aafd6512c964c25dbbc0a24a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f12fd50a59e0fa9a8e6ae2d436a9f835c49833715495d79857141ce80c832d478338c23fab6a18234bfa666be5920e84881edb95e9b18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fadf46302523b04f2ddccfe29008d7349cbdf122d8dcd8abfa8ad18299dd00700a3eb76b49222039d543cb9a8b492202771d0f17145de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1dba8acfe4f4aac73a837ae4fed8507a9ce61dc78b83c526e3d00a75c02b952f777c45d764f17993d7e5cc1ff40c102cb101e0a425105;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39cf465d57a5f487123142a3bf1eba22fbfdde2d2ae9b522dbc43f972c0c92105b7b1988d522178a6f7a307062127109e3ba5b01b3fbf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7cfcbeaa2df5c85158e3764b908d28b01c8b23603f480973387f9bd7885c6b5b041cfe903618c9971dc911fd6086f1c8b138ae8043249;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183864cda948b632c4b383e71e1b99cf4a96acdd39c2bdef06b78a7aec91b1326f551cd6129017bd2e74b53e027ce2f01ee9b6272a232b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a5953a45bc4c1c6c88f0c1c28baaa4db8d4566fef0b42f845d379c1f8a35994b4828564bf9afe8afcf482ed3e630d7a3afdebc2eb572;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h809f3e203d551c080c3349b263fed6ef987577da3bc847c5c33ff73e73745dcb89d817155f118cfeb6c6c97011a2eeb635eaec692f74ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bfb08ef2773a34d0d43a88bb4a5d21ff6c0c936133e0a1c917da46c03a1d61eb7b02d81d88ea0618bbd820b3eba454c70c0187ef86aa2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1450ee7132c06ecb9baae7d7e77afb475385d935f61626033664089126b11d67797cc60d6f211071e4cd817fb68a75165ca06955b03481d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e8fed02c5a1567f079763c1ce31cef6bcb971c9ab33798fc67cff40d3844002246f2487aba3203d537e3d7fa54806d89e87376d2dce46;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f66b54130f114c31eca128fffbb8d2913ef7f82a05ad873ff3af03f79a726990b6b4a1a1aba76c8caf4e1469911ab90f52f60ba9e95fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7173d3a8718c4dee7134ab9bac05a8de07959f75a9b2c1d1654adfd00efe0daba7372bbffb40f747ef5bbacfbeaf6346aeb7324a298f89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce57d7f35f72a73b70f90ccc8a84952f84bd8e2bde1518f3d9be725260bc7ec24d25c8a5eae4267199049fa71bc44508e9925823fbd4e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6450385bc21277d4ee9467c26276780ce57e64f90aa6be3bacdc9c20b8057052f4061a6bb8b47784024f368bd383797112c50807324a44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12cc08d6a98cfecf4abf9d9728b79940e255873ea945a52b47df4c7e2e2d627d212c0c09d9c7312d2938f785e9ee93b843339090bb521aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c96992de6a0f26edd2297f421652b45ff64200e9d1f3cf39a76654cac26df61a8f99bc524427642fe6c6e2cbb502b11cb6f6d7ccf7796;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a4c489ef01d11caa503a544affe588a23d613bb8e524dd447b733f41fa571edf544a3645dad7d3c6e3131b93d4fc0bea0e8dd5dc322b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e85ba68840169fdc2c226c6d3b21425e1eb7f6c0a7c4bdaa939bf88663f2c1fb712ebe87cd18b5a9bc9aa12fdcb3fe20beda28d1a1ce2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162d37e999e469818c8c491fd33915f5778920450d96913eea31a78a77b93a27b3106a6e5f1ba7bd458c63d6fedd9b7d65353ced67555b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e8e6a0bb37680601adcce18e53db635c461433012a178b99f3441d93978df5e990fe8f93f7acdf0378b6c1e59c8e31b050fae54c9a616;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h948cbc6a5c3f11c741758c1fc55f3b9b7c1e0e020eedb75f1f1c87c3d4492bd801bf891c48a0737fe940493458727a404723f515b6f7ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131b132a6ad733f049f267d1fc4f2d3d51e199ec697233dc7eeb40539ddc19485a65a2f889b4677c3a4122272849d35c4657f73bba07395;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0d3bf5bc666da6dad25e4d351f441883de40662f1b4bf7355ff45d9fecf87620d47331820a5d5ff906f713cad66d6b8f379beeca9b0af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h789bbdebb79d1ccf88a02837cb55df378d42ee40aa6bfd3ef6b71f889528b3f1e3b9234fdbfa7f5807aa8963e25f66b00c3bf503f64fdb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6073e82eca953514b7c5506d39bdeb1a2e857b82c2b65c02bbb2fc7ba55bfa310f531f7e24881cd01a27809a706ba4654dbada86c7152b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0b063566fdc734552261ea5385b975c45689273502db3a0effe1853e57dfe5a856e4919dcde376763d03aa7401c0e10df529acca6edd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heccf763b980c5d8b3e3811075d6448c57c030b600ffd8697c1cbb5c14c5d42eab99cad61ad6fcaa8beb5eacdabed34934f74966346112e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7a5a53c347af494f47fa9db2c4737f825c1edc9834c6c1cea5c6f2abebd33ae30f662a93c88f44375d577e4be8971e138545ec6bc2aa5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e2b4eca1102e39f5586d94f978783e824e04fa0526a9e42e353ad96ea8b62755c46295d0dfb887f86598e16f5ffd704c4cd7ddd6db1e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0da634276cfb1da20ec5f23d0dcc4e37c693fb1886b28732cb743797c7a22fd17f260c4ab6b7f225ba0e18a33e2ea145a9138691efb5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1031f18d4bbcb7c63940d84689d6a01133a73eb74141ad1a61e11c32fdb3e8d84f310b2d42fa51e0f549eabbbc8129f93bec94247cec9b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f5e2ed224bfaf4dc3811d58acef7429d295a0caa7069599bdade0e3c031972d68dfb0cf1e172925692cc7b6f7ce2bba7a9f9ccb673eb3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109bb9359d888b9d2e51bd9f744657eef9cc08f360cdbd6b2b2be53711f895c973d1f4a5cdb9a840c7b8685d427d0bfac0c5a51afd98234;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd912632e0b66bc5d158e7207f31be97c667d177b3e346c72891f70bc164b50505325f6eb1c8ab6c82d5c2d53265faadf5967171271db5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2c05c17990300845b61b949f1bbda78329c0843c2e656bc7bebcabe845248cffc2b47d66353de5bcdab9940621e282003d2c19b92565f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd44d1437bd590b57f974a06011fa07ec0082855b2c5f809d4675a8734a92625009a1dfd919e4577159ff6571116974cac26a70dd4ad2d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4b991eb57a6d0d75a0f020ddd30c3cb6f81bc4eda711220c15964f3ac8673c1e2c5e0d80531aa0f87a37a88020aadc697d82060c01189;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a8412324523e61a85354729cd37b552721cc79a53291650e1f52264dd43a6ed9aea80a3720409c412cf6c1cee77acc02251ebca24d501;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3b27a43259791adbdedc6001c5a4aebd120769ce8dcc3808b9347c3ec0dd928f1186013e5ee72c7a192a79ea6eb91b94d5590017d2a7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbea0dcb4e6398c6632ad91df3ae16bb70ab2cda913df469312b94b759586f847499c20c65a45b0f2cbb88efb267ec4d97d54c18ec2c12c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16334e7355c4d5f99c5a06caedb19f8739dbfec59780bb5e4e4d9c5c66b9a725d126639317d1ff884c23ff64fcd9fb415664ba914f532d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2ce06388693ecb509b5d57cbd3541556584953956a6ab6f60b5c4381a326cc4d47f0e044b642bc2c5aaef5107ec8c720af85b6a57d567;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h225cb769669750af87814db5fb568f9a756a1ffa55bcd02a432adc85cc4595e9499d065bd4eef479103c6fdc6d4311a2e5b30ea83ece47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c355bcebb4adbbccf20e8cc7e47757c222e1dd9752ab988c08e5c4f1d4c41522afb3f55daef61de7f16c9daf0b587c4bf7907d26fef43d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112d23140f9d2ef76d0d56492a8e9fe4928846a8c7e4fd841925d67aa54e85880f3ca631b7b7a04ab2ef4436081bafb24a9395ceff52972;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h514b8465ef9d07541abc40d6f6a5a9010e10b5728e9ecc7af5ea4e0915ece35402efe7f230df3ebd083e0bdacbab6a5bdc549c26a19cf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1215e223fd3a3614a053f2a1f16546d156a7c76ba6aafd96a809d5a58ed832d5d9ae5be5f08cbb8ea6aa12c1a8019317769609011242821;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c420b20920d1c491f5bb67faa2f6dbe5bc9fc7ca32d5acb45ffb7f9fec46eece463a233f8d5d24b77087181c7c71483810fa2e873d646b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a01fb5a6bdcfff9e1f4514d923bf18109206727c1af52aedb469e02f140ad447c62ac30ee17caf8a628a44cfb41d39f9c21787f01728f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b2a3b5f4b1f61d547602721d6237a2e26ad0956af98633fbe61f645342b0c99fce5fba1d5a92c7c8a10aaa055bff98eadeaffa3f74514;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111647838611f1702c33bf69315bbaec24311e9bf6a83829310cd9844c71365f15a13a6fe261d4e28fc34155450fc5b78c002fab3b1505e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8603959c356804a8d49fb41296feeccd2049037cc9e6b6c39a86bac6cc964cd1d3fa78bb170608a9f79ed94faf54d916729003cc6794a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1f57e784781ec3605723a90d577e2adc9675e533277f9ddb3a88318ad3d2c81166c067b75adb8d6d7d3586b25985670bb2995e1bff2a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d473558222991f6b22ef6770cfba4af47352e28c4dac2e19e1cae4dd3aeaea0536c2810edc2d02796f8b9744e37d98e3407876a7f5dabb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb4313d6cbae4c19525b4f5183c2bd98f68d5cb9ed6d0e9d9a0634ca27c6bd828763b136bf22b446ec98d623c6243ef733edd57e925697;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcabe7d6f82075808e47bdf0e234f300aee6e17a298e4310f3e37b7cb6902ed295d8d4c215f3002b0d19e4d656c01ff5d263565e716038;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1063a49c8bd509500b18ecef392e080ae29f9091f15ac7052585342f2f4557def071afd45324e3d199085652c9d63d2fb92f7d99b1d70a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb01023ca7d3431bcf87ef8801319f1acedda58d6cd540f8cc0f44b28856deb31ee4afa0a1165d565c0d6d02a3334e91f45306d63d6bf70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151abc6b56b25c91de811215bd3c1dfcdd4416338501bec7994e81923b617131fb6c3920ec6f1620aeab075ca7654794e60ca390cd15bc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he624149bf218d3a3b5f3b075f19f4949453b28995a8da06a2d65b48a2b2fa5193cb5d0a41f2a65a930ed0040033e2bb001cf5fd862e98d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h759ccc39ec7975433dc5db08cc1d1df8702a1c24e45c7dd011bb5a3cfdb06655e8513663cafcc3c7e494aa6df7b29192ee0da6db7a097c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1edfa3acc01bca3d3e3c759843767d1739526bb9cd78694cf54efc7b2d17622ce32f5adc1e4fa6432664f1c33eb2e2a5891ba713d96e2e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5330457f734a7a6b0371657cd20256030f16db7c79e8edd7a08dad4e51834441a7f6e322641922c63246be07397cfc60202cb1627ade95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197b11de5beddfcffa9acedee9657b0cb7ef0828748a9fa959c596ab424a377364e8536c1930782654f7ee4518d4bc28e76b34bbb5b51a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1546ee8faa4d78beffda89b39a36068b4ab2e5425e6fb17de9411501aefbcab609687d83364e97c53e20f8dd2b53160bf2209d4db9edef1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ece1089c00bf83f2995f40e726eb5bb7474f5bb892844e1a229ac55b961bc3c6fc3ff5eef85dc096961cd3b2d68b1e25a7265948eb4220;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9822c32ef23b43719d97b4a57b774415c7cbc94f57866d754802ab2b8147579ce7229b8ef34e2000ac1b579a6ccd7e90d3b7a5330ce46e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198ac3186e7ef706880f1aa3dccf5f3f882ebc4f316262225652751c58453ccaebaae44daf85f91a83d2bb19be5364c4967c50d20717e4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc45f767ff21192c6f7fa980ef97458a7eaea3a4501251178f6ca6b6563c87bb239196ff4f444688aab49dcaf3f42efa0b6da3afc4bdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151b07cc929b66420b1f4824d5ee7293448037d4380f164d94bfbb2e70cb15fdc8afcb5aa3b4af81d665dacf7bfc13439c3659d92e274b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4768a6b5206b4076799bee46720648703822103848b0175a9cf861d213ba587fa17f7d816cc4b01e1b881dc9e410ab78581c332083cd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0b69cff180d3fc1973889d9f61dcf2f847d0e1e9a532bea3827aab6b9651eafd9fd9457a2d9939b0005c98a6c5f762a91133a871d7ae6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1395545fca74969183cc2fc87199370f17440367f562febf68b449601f201a5758f4b18588cd13c8e8fb9f8e0784ee8a119ae8414c4f4d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb92c010f6fef924ff294f2e34db32cc95974d72dd3e206d8b10f08871105e51ce5c98aa4007e8fd1382344704536ea3e546b86eaf403a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b25186bd96b6291264e895157642af70335d285c4816972cf7ab6df22ce19490194e962fec365ebd68bc8524fb9440e51df3f44fde5c0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62a339842262358fac64ef478d486587f4bae6c6d4c25271d8b28117472991ba3fb91f993d361a10a5c32a225e49479d01cb45db94f91f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1812ae8c6c221eece50d1d524491f5eb9a69c514bca4100f8634edaa7786f31a44b334ab28698d219f4741195a0c592d21efcda11da0c2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1650b675cf82ad7d866ff9e432670ea9a651fe07e431f3722ec874cf0b9ca5b9beee1e17269134348592d3333b00126fdb1531878a598b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c421959d6942c0923fad7706971ddbb2711567cd64d1de346633e230ebc452178fe6c693d523e7dea6ae5422d89a967e910e7bf1fa52e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e9c67b6f56af2295c1ad493d0e9ed5198d81e12eb132ee21ae7112f1875586be50f0a8aef6d2188e9c298fbda789844aa6ddaacbe2783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44df4a2cef2ca0612125807acd4dc4dcc267ba4bc426c2b9b85a49ac86c7f33dd1d38e1198f127bb390a6aa3a13d9dc43a1a9dc3aa8f49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h873548c1cbb3888393f46a87b9a15ab9e2d35fcf1cb5fed9fd3fdd1c82e0ae4bf2afa0d29e40cfe3d1cdce525d2137ba9806b0bb08d2eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fe8f47e4ea7f48d12d8e2042a383ee2a2b53f443408c073ee1b0932651a3d9c57e53336455c3da6a6f16d1f75acf60bb3025036c3af7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c93a7ef0ae963633dc3558b3523deacf9dc41468cbc5bc403f8182fba8a9e7ae647f4827776c64bb4460d5f2b548528aedab53cfcd6a1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cde80849d67be8d7117d81416a2c90b46ee37420493a322bcb404f0a494b1cb1947a8893c3b97144da750d44a8a80a253ec818e2cff215;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfc2e076d84ce36636c2c34c8dc82a75b740804faefe8d4cea374c572b96320d43011ea479b17000e4d240b690208b6ea79c29effb200b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b45244a991bd1913f8de169541f4c43dfd300b2dc5c1855a3f470c83d717327eb102f49c6914118a79f154cf5ff1afa39f0f69306d4e31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf472847a16aa07694aa8ddd0081de258a80b87ed66ead633276fa2bf453e36761a177926a11364606672b608b1ac011e722707ceb8b76e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d41ae559efad2181f4a07a9a268ee4a2c5cfc1bc658e583ed1e7af55a753536f937bd9709884b2f69934b65d2dcf0c5229bced18a1d969;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8528384b289838c6e63c65cee037715b5b9716311f63cea80aa8a8012dd574cfb5d1f492c8cae5f1b1e484705fc9968b11de1d50b9b89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59b9d047095cf768b88c8a00a96d18cf05cb9b3797e8b4eb3adece7008a246e4309a0538be8265e5331c897106d868186b5bf8d8eb394;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1215ac496d5e73e9f93ccfec9aa9c9c553fd696d7dff0b678daa33b53f44fd1ecd4dc4612b5076c136e1ab2818a53455012fc683ff6f3d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44c880299e5723d6beba3649897e5baca59d865b3156f90825d5a501c671332f30509fdcf349c3252a2eff0e7df848b8fef940ff04d46a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135026b65792b9522f90b4934c269c1d6bdbc269835829d254a3acb70b42c70c5cd76c84e45b618b80789a0f22ee4c88ce2b00de0d97437;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58b7b6c9b4e8090b2623b1572b50dd34c0c18618fe4db2a117772999b465617420d3a288e77bd39f5d26e6dddcf31a6cccd073fdbb4e2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e74c47bc66b0c2dd3a6bd28acd732b01a9e8c70b2c4806ac605a3fdc82d41c24184ae1694778691c341fb6e4b57b2fba186231b2cf3be4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0d81173b840deb384a6e2f4836b4612e526bff275297b295bc90a127f878de99fba27caf1a2579c31f920c80bbda7008c4cd356c1d68c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he786a928f176c9b97f6a0e5287723069ab467009b81226d46fe689a4d702f52547347f335fb5cfc6c14664f0ff893e84d67dc7403e24e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b15b91e2c6bf187f524c42c3540f366eadd3ba677e9b61b620f227266b12b00ed767229658b76fdea445310a6d46883ca51f36b48a9cca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe153f04df77f67b0f2325ae79fa387ed0caad2fdb7b974cd2e8557cf28a341d3e4c2297b4e6c16a0175f85827d580caf4334da43ad8fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cc28f601f24e69906194e50af681d7f6254b207c23fe1ac141f27d28d9554e587eba53d6469f1f45d903905d2fdcd10cd46a1385e5574;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1914c80e05e95548773bea6a63e0dd42591850f1844337ff7158f4729a600c3897c3cbbd15901e1b3f0afb2c0b7bf830f902c8c9ff8de1a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc0247eb5bc5c074478e49a15eadd9b877707e6dadb1809ef5bade428b81a209b46dfd1c200d18c6af01b01424285f55d570d49315a2ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106bb4f70452ef35eada7a126daee100edacfb16065a20924897134c55e8a238905badd75de33a51f5d4a5d91ec7861a89c5fc0b8492235;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d7adcf50853eab8cbdfe8c7c5d9d2f311f637f83a3e2268054b14c7b738fc6e6058c49b3c8544aa13475296a4ad5353320a81a87b4b7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198973165ad018426b8c5a9231acf30769176faa77ca376146f611ef4b6da62ab157d9c0cce8a57f5546565716be6241840af4b1a6dd939;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161c630ce915324563d05a03ed1f088a770875526e15821243c8c98b6017a1d2952c08ecdeffbe5dab12b23dd7b4fc52d3a52361e3a5daa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1f5bddff71be53e37d9fcb5e4d9686ac962a75fddd9eed7803475cbad707453ecbfc97cb7a0dc09ee23bf7f0546639adeba909944e6fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1770f8640270fd3406c1ba9d8f4a09d9c685897010ca53af227befb41b03103ef6c92be39c194e8c5c0ebd4a695fcaf5498ecce99c1e8b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7161dc234d06e105e364f11cc6c9352ec67b594f35967b07225e63b5d6718db6218800b1c8a9b49f7c6fde99311126d5d85349335bd339;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7bcf656d34e637d790b129549e6dfe24a44e3d6cbdef0b73e5ce888486b92e77408b1a7f352b7bdf535370243f034f8e25d446a2b93bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173e0db17491b357a4a6742209df0e910f86266bbe820e6efced3c20e24e7f8429071f33d0f3604c0066904fc7f626b5391b385db28e08d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b9676f98adb6dc503926c804ff5071f3ef76c54651bbe70b36d0f8cdc62299d745a071c12abf5151122bb4c85daace6824c545210d53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3d3669d4aeac99d58210c9ab515c9007f94eceb4c6f7f45e9023babab7c8ba51dad097b3a01552381605591663ab2386d20722058c5ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1def710fa4bd80f568a8b36bee6bbf534a66ff8e8e0248e991d46a81772951a5be7c2ef92bc33905c398d1dcc5772d1d5ea0f4c4a9d8e20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134808aeeb75dc1c2e97724a2a84da2fe1283ba07e6191cc6b5e558de73a2ba891355dfdf35f1fe0b0c311bd7957eab5e696bf33537e2b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4b723190dd0f9204931de87df71b4d103c25c09b63665ab551c20a4a5aaa87f9dd6f73ce7cfa883a43adac03a53e434e24fafc08a549b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adf002afdba45305f8023cac6be5692afb461a0e2c1c98287f273de88fefcb755f7e623aa6b41629ace7472a29b8d83aab8f45ec447a6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ac3416307b76c17a3a56d1293b5896aa9601e2504ba5c8d0bc00d46f92f84e2283ff8753e0a59a825c2be4a2a8cff06ee22401bdb05e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbdfb762222053b190e3406e43d73f570d5452d8f8ef4a56cc4e4879551c8e14f323489cef00684ad1cfbc7b36f9fe6d46cd9b283e34aad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4203ea85a68696293c17759067b558f019da3e1033663439b87c145cb8b3cc12ecd8fec3af18dde6c0b720cdcc3ecdaed569142c960735;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60c5ec5b3eea1ea1db30e69b9faa958b8402990caa2b0ac50e771c00b71820410443dfe9d1cf60c8d40c0cc4cc3ec22a991cb0dc10dfc4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b3366cc312c4a2459ecca5c9b0667e107b0d02f91955333cba9e80fc1ea3522e1217f93dcb5f29b6d7f82e7d6a1519efafd31dd84ca0d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78dec1cdf2c7d8918a49e2d1b72983620937b8e3282f247cf2f0ea5e912587382e6e893719c4dc452d5df18da1c83029dff62e66caedfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2672a10e6d02b77ab8dd63287b532882b69d58ab3b08e8cc06410b109123de141989a15617f0dc72b81381e459402277e7fa7418b86a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0f400f2706ccafdcdee1e34cc6f2744f201fc0de6c8a6ac7864dcc54d8cff42bb417592430faeb96f757ef6cb69c51fc56f879347a3ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d76d781952cd0b89e19d1ef28548fb8ed6c086b9b3a6d0bf5bfcbab13ae06df769f32f711a02ece1e00ff54761bd82d302f46f76f9e91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d9f625191c61b3e01aa23153ffcf7725301fe4c06addba873e8bd6dfce841c003793d3ba083e8a9520ce1c434bc5ca5fbafa19ab5365;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h828c99860d439c652a8d7c53b8bc802367671bf7f9674d48d4f1ff29f253f0c47c93be464005c5b89355d6811a789636d89aef88674263;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9be8e7a3808f8329a83cea76a5ed06076a6b8078e588c7103a3db0709f469fc040f68e39d8276c1c8c3e9da192cff481a581f7a43044fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8eac4d3be0e71512e5b7cbbe6c927ad981ca05d398d8803945d6b678fbee3f49e916809eb985e073a178dd56771a34a3ec6346a8a4425;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f8ed20a33222ed6048655a2b64e231a3df0afa14f713ed3df1b9cc06d1d9300b75bc6f474e4bf7cc65eedbe5e3b7c225459ee37fe2ca7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1d674a0d283ec18b1746d47d00bde990674b6dfa0d2cbb51764fbb599d2c56820f46e93d9a78a67ebed0dd894dcd2c1d39e02cd078624;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109d8bfe1028d91d5a66088135f2999af2d095dccfd50f81148f4fb85affa3c72a201983cb50435102d8a47ead5b5714bbd40a299e5d091;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2fb31721e9eb3155586504b7f97dd7783149ae228e4695237d790fb5f08f4117883ae31535ab6ca93c650a3b20c58ea6ea2458669d986;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6285fb900090ec34a8eb4a170310232627e8da2f67fa95658c341424a50f34de839c06ade890e0e31d07bdb14cd11a1a8d54f1e1ef4ee5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1b5d8b049b6a0b0f915a7ca196d7a401540ecf8f16b5ffc807ceebdfb4d54e73c28b1c8152eed22103d716b2b8b444c35feda50f88309;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a7573d384983a718ee906fb201c0d054ac222720bcd64f3afc8abcc3e029605a6b6d1368039ddf4c90b6d8ea4b51c25e243d8b783f3e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c60ee2da1cb12caf74a4ce66829874511392f3ca6357a08a8cc7b1be052ebf0830656c632596e91700ead27f866e45f627b201e70407;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1291a5a9a8166b553e930aa94d6ced7082e8c23e19557604799c69a45c685a53704127a588ff9d2a71a31f86a9fe3c3ce92f49a7be30ed4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118f998f76b6ac00259a9832f98098619b4d18a61a6f92377083b9cee176f80abc194d5467eb3a571dc999537136eaf1f2eb9a25328af14;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcce7982c590d33d827f3213261efe926c7b2fd6cf7c91deb2d0a220f3a79f455a8c723be2a6690ff87ac8185ca995728b3b8748cd68fc2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9ac63cb3f04083c4631a07130f293dddfa5f2aa1f9b026ebf8070713248e68bbe792cdd326daeadd218c45ba4c71d27f53b9679f2470b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8690685e1a028ee4c40f413772130b0c8c4245f9b83bd3fe7b231f31c5ffafe4fc3307bb4bea315a5163401c6a59f8487e2effe3ef681;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9244f5537997e80f2f0892bfaa3ef2e8ba42103a088a1e8bd8e30ef5152395976954742bdc5d71ad709637d86b672f288e9dd2f04de16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4a2b8a69164b82329e9143b0f5bdd4ac9972930155650987185bedde3b3318ba48e06b26460192718fb79c62413ae9101d5bb9c04c089;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ab3068a2a3352814551c415085fdab2fa19ae11f359bed80cc2f7f8739b3b585b5eaea310daee17dac418a781556f335795ce252f5379;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h212b5b2a38bae9e7226da58a3af2fcefeb10ae1aa8f47b9d2020d92dca3d0a3b0948c7e35e82e8465d0e4b1fef3220af0b19a678809f19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2c818a8b69018b8a7e68d4c9bffb94a92fdd49c5948a73d92791b596553e9423f72009fb47fea3e825d39b618a2b0de64ed7a6f12c65a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c469a8df287e33f931f46687e695e902f510d2fe953e20361bd1d97a69019e0d5fc2fe9726ed3596bebc71e7276ec894fa6145005048d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0d2ee9cc6dd5d2c0acf772908ade38ddea8650182342785cb60a82a886385dc1fe601ec3151d646246242ac46b0276bb37abf79645f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12be14fdda81af44af6f3a2da1701903d6d18831799e66077fe02dcc93fb98cb20a8206e7a67dc9c674d53a22f90abbb12f0d5e62d86543;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c3fd70b23b46b061672d8655f43be55293d8ff91a61fa1ac74db90e6db6f47569cfe8003abec0d375480bd7c767b6b19b0a0899658a1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7dd4fffec13801cd725e6fa5ddecd3b967150a64d3ce56574bfa58961f8e8a9bac07b0752b88faf82694239c44febafd0c00b2d60d06a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137abf6465db16a45892f8ff38a5e1618c92f2a7f67a02ef6592b1081e9223d968666446559205919ee9f19af325768772eee3c64617101;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbef27f4f9bbc9e92a8fea47be1dd5134986546aa308d0d0b6baf718dc87e3b7ccb2fa00ab0fb174eea0a847d32e7145e347b4db268222;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ac5c007e7ea7b75b4bf445973e473b4467357220c9e62237f0d4ab7aeba09b39df0c2070a6526ae0911ce22e6bbce0c13ef81770bfd79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86da4cae163dfb51bb2171b2f79e12f9426a82a6b5ffb9ad0811a9538277124dba8ad04d450b5ece80594ee6625cb80ab6d11ec52da0a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1926d80e1c42d1de514b59fdcca9628972b4711e735250832fc6f70f259cfa411a9402ae90fe9030e195fdb16dfb424bc5c575944e44d09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c28da32eda73175b9a6d928438541e7a8b38b9c1771ffd474e8aa0e9037898fe70440f7ea399629cb0ff270f34e3a6811f5f389c46ba23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd31d24adf780f6d1ac3be9dda93e3d8e2473e764180a2b49b4c882f05d570e985b68090ebc82780a102839ea537c9d2d15ff1bb3e1e538;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1352b8bd1ebfe3cf69a07c24664077a1faef2fa413aa88eb484408e67eca2a884065e326fc7db79c7143a9c7b76801f039459196dc96c28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194a3e0986e9b456d7ef63ce6662a9fa611df4ab088cf0ad08407f43aa3fd149e295280dd820413a04321dcca656d05bc9d5d6662da07b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfdcfc070c264f4e4c17ba48b4a4f2e24257d317c9d541fbe8717a5e77ebdf7144faea31b0f9225750ec44b4de13e18645a505e2c6cf452;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacc4d29a11ed0919a54ba9db688eb351be5032ad42b0ac56b516eff118abcada80d0cd3be27aadbbc8e963538ff573073519c48a80736f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b38bdecb06450821f956be3cbe0fb5855c5e998597dfaf168e35c33c530f2b43b825cdc9d1b2a683136916fd9bc4a84b2e2f8bef452f46;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h158dfd832b786a3f880c0582e3daa11c6c16c41f642d486c4705065b452bebb3ab2d7627d02b0a3b0c628630435a8506a352cd6ef7a086e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c91c54491db97444e18278aa934bd4a112105960bc03700ae5759ed4552ea14e21ef9e2f7ea67b9f8ffb612c40973ba50ea7d712d3b93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16fa022b6f9be06a57ae5eb068938b18e8673405edbbc051e0bb49c84543d35cb2ce96cd98763937d1ef1c9587067344e800f42e7a20588;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d173022367e52dda93e3b8683dbc831a908c9938bccf3851db504c1b8dc042adf22186223d59102ef8eafa88d95c14b9272806110c5f3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fffae3f662a8c1858086a2d8f41eef3d1b7eefeb082a99518dae5ebc0665e8497fff7848fff60d3f0030d2e491265f673487150e5d18b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f73cfd67a2315db5d39dd63875a21e918387f7b2bd90581589c207078353012291f2dee1c22e90736118b9f9f95de1863232c0b1656f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h467cb30aca259385c19fdde80861cb64a889ac98eebad5ef9dfe4eea7d5e084ac23086fedc0fed5eeaf29ba589f15f21f800a851d39e11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed4ca04cce894fd46e3c47b21032a11dcc3aef101e0e53ca424355dd2b3aec6ded66a9213ae950953fb5668c41fb4223dbceade7574473;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4dabf0fcf80fae654897f900011ecbbccee18a02c8788c5bafbfc11acff006df1bb4b6a25e6bc11eda8e24f1441813cdc44bbf96a1bcd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0a0fc9fc90871e1a6e753c26812c03e4117be7cecc7d5c41755eb07d32014d1f48c60e89b639d28a8c51c4c02089605b3b1056bd56764;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he45eaa62fdddd4869838526cc8fe2b96f628e8632c2127da45d362814d129da3c23be11e2da8a9f29a987073e64e820a9947d760006f9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ecb5436a2bc71d388d082cabefbf18943e91e2c450c3e1c8d524593c635d92027903caf858f2a348b57908724f87cdc7472a655d008bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b6807a0db8b374995e8997edeb2a7ef4d2730900bb12945ee731d569044f3958feb8e5a44facc8c725b6431d23a0e8cadea003bb860bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbaa86832a03d14b54e0330b27b7b2bc83c7d6b560a56f850b82228c0456743e2503a7d75f9bf62b402deeb13e919c0d93fc4ad4e13de06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127253cb8e9885eecc65d0fc2a5f7f1b6dfa7b1e121b543e764c0bf79d9afcd633e61be58e1a711d5faadde9639d6b4ab0b710f338f4944;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14332ee05414f9c2acc2b1833fbeaa52a8eadbe839f63236152bb75a26dc60e2050313620accbe144b43633255d814467fe809337fa9eb3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b5da8a9cf116693a4c8efb21f7a5560ba92ae85af43480efe8b42f81374f0d3ba48399ae39f9764d7d7d7b85dfa5f38c31908cace0a8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e80d325c25537cc1bb1beb1d54b5ea809965a3958cc31c39d0357c20859a6f3428fcfbb41ab6a946f142151eaefb71d00119a68f0c5d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43fde67e81d1854b24400d156e186a0d5be8c347bc7de788eb290d4b6c9c4314e9c4e34a2d8a7a014bb2ed605f1438dd0ea9de5cbe8c12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d771cf3d75a554a5db2468d9ce3863694d820a09d2d87b6adabe217593ba9976eb95dc217dec77dfa8933df18af45957389be8ccc56a6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91405e3eb435eea8ebb41a3693b12d73d584dea593185913b5d5413aa87570e22d11fcc7ff68fe36a90715f3a14b8f413eca0ae8a47015;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d8d245bdad578acc7c0bb616473a15b0accc152b541ca64b68c8adb342817678d325e2232f82bed35d39bfbd50c4cc20581a6965647cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5966683cf358808a7b8f544dcd68b2739a43954fa95f6065a33c6fd1f18f0d647478e9c80a663101c51abbd0ff0e9d834037589bc7c39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184be732db565a2902abe2ae6878050648e36e80344dd51e961d0a97ab0daf0751f4b983912502df506ea250b07aae64bfa21105742ffda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5c68b1ebd920fa8c77d1d3c46b2f1b7459f8c4fbbb8d46b34a1f84e6998b845a8bef27220dda66c678bcc4c5e00193872e26e3912857b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11061d51f80060b312172a8863f3c8de7161eabddaaf703c59d75f0eb98b7096edee0352260445b3e9c0c0b9591e35517d0fb82baab7e47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccf7d214af247c9b3f09588600dd514afb45deeb1f10a5ebce24e4a81991b3c2d71c1ff1bb88692eb8afbb2910a195cbb70825527c3cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h600b952529a1f9f79dc123bdacb49c88503954e5d916c0ab3eb2f61cf53a003b1b41f53d9fbdd641f5239bc5bac319705c748842a6b6a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bc0a0b54724f0b5c253be86346338ce5e4547661c84fce719ff134cc21973b82a88bd421517f29382bb6b882555546f25405d52cf528b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145b47a8a260896222304ecc36eaa459d807bb6c90e0b24af7420e574f6e661c0d559cae442d7c30f6bec3f828e22f73d24dfc59caef875;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100a7b97dd6b3e0d4bfe2706614a8e40f3c9d9948648326f97a389f54e1bde274e7b0b870c4208a24cda82f1fd6d85064688716c55208a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82bdb0138d66c56530923adced68885f93d3ed799dc673e571d282add5512354250821388b376d745ac151e71d4af22f37c21ae1e44d0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d30835eab1c2d1375d49e94f54e8d069dff2a8988f805ea3d9c6338f9f8c4cab117aca4d383f26802c4b55a144156a29975585360d9f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb376dcb168a5c78af431bebb25adcb126c12a196f9b1880b8587e289f27dcb5040899b76856771e1bc88e0b16b27355fac90fe4cd2aed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5aaa40c7945699003f9c19dca33f5a2b21707c0cc0c105fef9ca85b1bf50296b0b0a8ee02e36bc72b91f92c37a41a2e8e81b7b8b3ce0e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195ccd5722ad21b04ce1e1676c27698e1a208e751c6f9faf9d83ebb0386ecb0521126d675815f748c02dfc63096820615010d480d28c250;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbfb634636b4a459dd23081eb6958f5d4e6c9978f6c30c03c75962e742e11fca7e3d703b4910b342f265fc98cf3fa8e3c1afa0e50063e8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2594c39960b3420e4b7e76f4117ed6f7a11339dad4f0342fb32cdcedefa89b98b8a8b7f3382d9296c142e29bf94dd51e532376e47fc43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h392008054c5475780ff86128e25407837050f04989b6b1c29b9038b212518b0f0181d17e4df876943f5a3a329acf4354151a791f3e03d3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a6e6ad84c8f61d9e66f1688af0c74d0d82c4d3d503f3a512c57008d43c8c1db4196c21723946893f9482b0a52e8aec9367489655c4a12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f80ef5de250e33e820f8ba891b9cd651e4b6d658002852d447f9e1c3c4f87d2bc03b4a91cafd2bfdd4fcee9a8093f9be79bcbf2b6584d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adae55c45366e40499f6a35da41acc5a21824add5a4fa33706b8e2d9abbe7a160216951cf70bc6ebbd70bb837fe6ddd95ed961c695248d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h514cb987a7343c768e1731cfd1f71143280b07dbd7946cef4be095323d921375e4e4c6da3800896c67329a1d50e86afc15a3e5ab9e9c83;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he48aa7edcb6c7b525af99760be0ca93add76a9819ca971c71d426a8dce31c2c5d4ef0c39d208d40a8baf7f79eaa92ca0a85a224e9e50cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff755ceadbe604a40de4b840e1b28f8a0d8c37426dba03c1b05a6ed3b2ecba2f32d93f8b9366dd0e8e9287cf6af6c121e779914a569a12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6be2e78f4ab2f746ebb9e22b3fd15b6ab61df06b6355ae63315a08832f898a6b7ef4d7184c36e3efdaf20a6f41478685f6b7208abc4e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb090b60a2befc7d5b384cd216457c463b07cc1d4dc7367478f93b9cae2af7a4eb887f28b8895fd4b2a17e711a42bca2f592d0b69cb585;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb1c01bbdc4f112be1380aec6547b5b445f8d7cf736e7ed56a9890dbc690c40496419eaac707da4de4226899a9263c117366a7fc408f47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198b6129f3934dc649e183de4cf66718043d6a0704ffc3c975cbc3f8d75155fda5a1b4ac9f344e7977e2e444477c457ae4e205c212f38ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15469afa392bb4ec9364129910fe7d35a5ca143599184f80677214390e16f9fdc8bcdf04f60094c8caeb7b6e3c60f888d493155266e6197;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea005913f29c4d7e5d392e80d726e6e7bc1199f6c5f96f40f059e5eb80ceb1568cfef0620b2dbb57359c62be12c2733c0521782e6e7a16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61a13a68ef125033e699bf98f5197900f621112ede0d8ffd0da18aff7985eff35ff0d9eedc0793c58e448e1049d6032757713710b893f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bdbdc8b6c69655bfc68a69543eedb0db74dc6bdc0c486716c90293b64c0091f594fd068634c26fbba428f1550212ee499aa9aaf06c013;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175839811d189396cdbab32fb97a5650945ba5f57f3a245df3e407277755d61d794ea141c10d19fb7692638edf4077bd7277169b2af5bb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121fcc5914f8723609305a1cc391ce055547cdb71f3af81310c90ff49eedb2c4c3261d0c0b682e335f514d70f177060717c941ebb9ddc63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159051c6f84fddc5c9367e908d89227c8234301f87ada7e4586b81d7ef9df43ae8d889df15326d83c30170eb84ca180251a0eb4eef21762;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105ec8faf7fb034b190480bf5ba96a88217428854f6e5351b50a1a801fc9e89cc057d161887b4c8e05e8a58ba2a1510d0b23b180e8cdc73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2075eec08f1e07f155af2b3ddd315a6c2b33df1bb7a28de8ea2b552e93eb263f03da3c4e4a50447e0ecd9433af9691e610cc78ec8e688a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc1eb5400862384dd50f062d009bce377caeba15b08d7398ff77cdd25da78462d3f6aa68d64392384a806a59c10af439e1b37b02c6bd1f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145bcb4475c201be95db6e3b9a725a55cc27fb8d388dbd605fb774bf54f3b1703053b4e07d9cc72788ba95902b667b669ee34e31bfff842;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c41a081c0f6f4df46dfb7fe9cf05e50431b1c65f9fa2101b19eceada966d5286d1d7fa8df4f597c0b768f25629ba96ccd285a671487cc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d65667ea410bfbdfcaacc8d5e3dd68ce7461738125fb529c4a59c8f03c094a131bbf1f42632b3780e7bd5d7f811060ce1d00a22cbc51d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13bea68650d891d2aeb34e7b7a40c1df12d4a36330f4c739ed52d64520cda987a1c977e74896c66938abc93d636927aa2a573594324d703;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1007bd7f70b13c41ee9f4b67bf5e675e1c2c67364fe16b11dd3e94c5ed264d4dd156a4cda1e75dafe8562839984fa8ff6bf45446500b68;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf19bad0d4dde19c0c71c872b470fcdf12eae5af4351a8d8a06c8324259df5243f51be9762edfdc1464b16512713220761dc9fbceca0d30;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14852b818f0ecbfa48f0f3c2aa15b8f08c3acd66235076055622aa070b7c9a72d5d104f1ca3a3f665e12bf6c0ecd5d7e35184cd3183c402;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1689d6b20f519159f687a9c7dacabeeeaf572b7780fd972ae4f6ca14578047669a07e3487f310258f8df5e515bda75753ea228d6a58dc7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec2b15b45ada362ec7495ca8bdbac08c92d7b0c7936ee8daceca9616631753402b9856ca7d4b0ce9270e30e6a419b89cacf132feee2f78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h304598d1aef5cccafc8e39637c5ff7a9c9efe2d09145208b03b637759a9c4ead903faa16d4e0a691b2d782d5f2995f46eff298005f108d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddebc995e36323ead581961e3ac9b6ca6be97f8505b5db4bb69683f57169863dde198a0c704a4ecae6250ac0ee2f0d745302b071e749ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1d652c410f1a971693e3dc3939979ea78023e98ffc415c16b3e896108518484c26c74d46c28435cba14236dd00bb43322e0fe711a30e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d8c98fc21a8a23e49eb4f919131607335b9798fb36f3dfcf0ec8ede54d9c6ce03e9adbbaea3ff4d1d493e05555eb2044e6059bf23c6f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca8548793dcbb6942ea679155617343b3ced9a75fc3ae102b9142662ca041a5acbc4ea66fb0f8cec9abdb1ffca52f6f2130e6371b09185;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdb1b19b233f611d42a0962f329e7c787ab97d5cc4bef349793e27f3ebc92ee2a6a85b2e9e6425cb7e8b8a3d32063b3ea1b3cd997aa0ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156bf2799ef812fcc51b4589c4e2da5e8b4150b0ff24b00c23b93d85341c8cc8dafcab824492d8314ce2b63383b0045575e6751b5c6c4a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145412dccc47cf044c67610c69d5c77d6dd17fcbd82948d840632bf06f7043e405bae55fd6f91c977b7293a0fa815a6e61303ac72f486c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc60febb27704dae994c3794170fd2a10110203c4eb86c7884377b17cf07cae56af12ce3f018442a8fe5fa04ebf34b67819c7c6aac95d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h337a320123235f6820a9fb6b063abd6bfb5d5a036d5132a0ed4ff03a3fe6fad98182f466853420a1906236d0c4387781bcf690ffdcd05c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5ef17a2d25b5abc6822e0857371f936e2ea36e0d39fad81da4b1f4861f93fa54b389eabf177464d904d50c9fe2077e00554ed34b4c14e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5086bb785c253ea3d941192c6cd4cfd9a7609043ee3b5bba2b059beaaadc96d4e69052514e1aac5ca54ded04afbf59eb62b92030f9f48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8e9c992e52401415ce99f4f4db06976e7d96ef779c7b1b11fedefcdc15b3b1b73fc85204bdf690389b9e8850eca4b5ce9bcbce9c506e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fdf99a3d7b55d13d90420ac12aa0084fc13726a813638b3a3034f7814c545dd416a77029449d818be39004a48dd0adfcce49a4c729581;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5a158d3d097db702e755c60e8627c9cd92de776f5c819788f4dfeb74ea04a951c8e0c3d26fec9422bf1587f6b01b099e5474b91a17fc0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dea7527140ba85b66ffd2be77bb8422a3721729ac0e8a39cd126b1201ad71e7a572b287bb153eb559926072c7ea72ab101f14cd2b751ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d609f32ba38e450bb5821530da58e7b71386896c16f1bf12dd52373840144c52b4514a1dd29f13cd417250365719d367926c77327755e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4ecdf7dcdf1fbb22c89e7a2899ed85ef591aad68bacda3078c991e83dd45df80011de9af4dc06fad4097c26db89438bd00c97a31ecc6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76feb0ad46334311fb8ac537de4190482ea150e75c696d0f24f4795bf9ae8192b98ba208f87a914b721627fa3c7d14ec87994b75d31ce8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ed9c47c0e982d1f08d7890265f525f83260277ab25d063285cba8492e23b07a74a5e88a657fb7e2ea7e9439aa159186d4c46fc6ec64d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195dc5b134a2ad0c7c0a4cf7853cdba1816e6d4724a225bd25540d75101280ba5e378881f7f7973876b9574829ee59381e786db37aefdbb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f392df8c05808f99fa44ac51375a8a6d2d084ddf6f70703905525349e114285689b3cbeb340159c89acb3505ee015d07c440e4af8a9f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81b8f1512af7b32fb3e86627a822c18d3b96196253c436f2a8452d0163ac5815f1d16cf802ccb654815b4653aa4c38e97b15920f7dd59c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45c9e0d5201e17d1f7d31b965c5738de948660949a2411956d8586a7c3266fe8f2d373d4e88614b0dfc444821afade2bd940ff0b30c154;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149536516d1339eb5c1f9e17b33425e3ac534f0bfa4e8cbca94b63084d2e3a975a69b4b5f0254e4ee277d44e4f6ee884d481bbcefdd4521;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb956c2ddf0e6351e37e732b6e49ae8ade32e2efbdad8f7c02537bfc5bdde22726d2be2ca57f92d3e90ead14040cc8fd00813f650e368a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd628c1430d89ffb8f32c6d679931238b82616ad8d7bc7c7183eb5425db72099bb727d674a6336fcbb13bc02dc6840f54065b77eeabe2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2536bc1c56c2c4bf086432f8abfe85cc2f04884a6ba46e409bf5c6d79e2272d4b308a828e9db7f183e7771be7efa266f372466efae0dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc8539207cb666f0eb01979d14d65b0346c5759b4057fb16a6240ae1be29ac571d8ef93fd250b5a78fb00289166bb3671bfefccf847d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161230f97ce414832eb1891aff8024151d41e65574783ad614fd4de6c901b638f67bfc19ca76c022d6dc35e420dc998ab73cad7242dc1c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ec3597c2891c8ffbbc3c6ca8f982aee5e5b14262bada0175810ba8773300915a80f991a7292dc262e67f6cc4c9aef36d9278fb880ccc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141378c95be6c92e4c3f34d71e2031e3e2c4a60bdd0dbfdc7674c8afae29ac728dfa40c8831d7d846d122d9eabe43aa433ae71764e0f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be3e3556bc163c37807f4f5ea5177b2d6edeb916b4a4bf9e13e5706075f7cf28612249e98cdbeb3ccd706cf6d27b063318f6db34315db6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d1f99f543816f0feda3580fa0d89eebdc6134a2cd92685ba8c793b66ea3e3de109cbbdde34b5c578bab971c57c15af84220ca34fd387e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b289f53747adac462fa55a6f841d2128883e2b2383ed30ef24d21c17654ec19e4e0ccca309de39899d2522a0264f0a00d8aed1ef09240;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135de9b076a107c7979519bfebd461ddcaa03fe8d0b8206554ce4a3d043711d11725d7c6ac87c5aa103236e1ccad23f8610ead03233a96f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8329a67277d5cab2e0f8476174db0b96db16b607179ce302e215dc21a2781fc4a728f742daa413df676a5ee76425cb2722ae5072fbfef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h902b54ea06c60972b59c11c8902cf924e14ed099ce1ea102136fba08e359664447ef53a59dcdb9dff58d5cf57b313b4660f081b882d75c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145c8669aacfec983ce9d9160437d3abe1394dd19062d380c3d5553ddce616e603c2ef1f464b0ee5ff4789bf5ab441fbe1d024d2693e29a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dea2842000b58fbe2220aec44e66237a5ba1764e00b2f2faac57647766bd061039874c08d11ca1825756e44312cc2442ee0e20801e3be3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3791e1e9cf3cb51524fcc11ccdd022e5ab905cba5ad73f018646028b6d92c986d7337f6f1e73ee2dda83871ec97a7e225ad9a23566eb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ce4779540746f7de3a2e85764db0bfce891c22f978f411cb46362a52f65c50412d4e1da07aed02501988af2ca757768510bbeb8def769;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f685498542564b1304901203863ae54d29334ae1d9a8e333948fc3d2d2ef657f713c2900edac931621eee0057d94ddd605ac8ddddb6b61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b612a1bd8cdef0a968b5f161b46e79b4d94d8acd08d931a3b73d9191855a73200c75a5404338aa884dc05350b40c7a0a03d53eb78b78a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18acbbabf5545d2459a6b1c05449806129c95798e63dc0312dd01e5ffd8220534907ef2de09bc57bc1806fce48f6b0a9aa482ca81d2617c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1035614ca2d3a7912c554c050fbf233ec8addb527a9ca5e8afadd581c7f236afd763bc8c030777cbcaa1b4ca133b3abb91cf1e875f12202;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117693bbabf359d14820dcb694f6312623f25f068734fb1c1e11369f29c40ec98cb8c11d243145a4666e1093af5a88ff07ad30ed8051ef7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1921a3af01c3c5445f78d554400f66d33714c994de6ba64beeb831451eb4e23d1501fe0f0a991a0d1775dc424957cdbb606def23581f708;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5dd22862afa8c6b62bb621318021f24326849ed51ff4764f26f1eac27ea1bcfc03d626fe9c00dfffe60a4c1fc425772915d94a4b6eef28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf27bf9a9c36a5588f1fcabe6c0370a2c3454e43ca0e56aa7a9bb8fe91ad43c02c2c4b48520c24cee580f9aa1fbd9cf84877cc1c4c90f5d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d9f81fe080a716b6b6b1ef45454869f2fafa012765c4a3831fa8e8616b4f39f24c2fe47cb885088f166f07f323ffd2698b989a2479dee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2906e2a7063f200d547a0b7358be9f058f2b2bc9560249ea12a126e6fb407423c6b1f6b2bfbc6883e0432c0328881008e6383a20495eef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be096b3983734fa6c1eec8e90c7c37915850a46920a6f0802f5c35067ec4829692b6f2c65cc71890ae98b1117f28cd98de3a016580877d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc2f99094b3dfce57ea76f42c7532ced39bee2a5fecdedbc6e7096ccfdfc5b7cbdf265f699a342615f3a2909aedf4ed389db7d59bb455b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h531e52bdb17242a76d5929124d0bbf8076c1594b7d0d1c0450e2f32d588d523e5dbb02d0bf39292e52e142408e3222c9d17784037e66ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35dbee9a4b5ffc2eea5ae2fb694b369eff633ef0a044748e0acfe800fb7303d78d2d3563ef01875fd0b26dd2a86d9caaeb8f69d66ed8cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170ad4ce231333fa75036dbf53d8d30951776927344d530e204c79195e6247b090ed34c95111c331f7c7507b22e242661eca917efed8f26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3aef98ec016d4e9b756fd7d55acddbe667a1992f357461342f8cedeabb5b40aa16dcf89f8feb5a52988f5d23e065e8dd6848d050c926e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c70f05cfed8355914cef381e4586910774854e01f92e31391b62b00bb15da6bf3af8e9f4a66d1142f9cba3dae8c460f08745e1984c7c0d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df127c30572f2dd11542e564480aaaf81e5500e1e4e0f0a7a687b5bef375c3d7f7f9070f69b57b4147a7811289386761144a6f5a7f989e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7912ee1a579980485f62a85eb793aac598433f49e5b1c00163bc5248df690f92874110a8503ff476767d3a862278537ccae3f432989403;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea0261a08679a1a9a6fbff864af7d8e2785afb56f831080bade9d3f81d02d0695181cc150faf5b7391d2eaa6d9103be15aeade4b1bfdfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9a68489e8487709eaf44e1b968c78d14c910cb0a9d5ac62f072af817bd756108a181ecda1f0c5d8522fe5c930eed8c39b85802c23a7bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140825c2ed8556b3d050c48d2d441c7fbef6bb9825e17e1a74c3377d57e60c8fe0743c41e017a67c58e9876d65317d37dcddd7d663fa8e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45f8322f5844a0c0f21afc3e74ea930723fa966c091161b7cdbc57db1eb03b77a16067265c04cc96ccd3bad6b251dffbb59d108b6a2959;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c8a5989561c105b1344dad592814dde0bb6f04c268aeb28ccf28559f5d18090b069d3f7fb313a08d589e682382c81a7d4ba987c5ab188;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6d582460d16f2f600fed4d29233c068df317f307a162585c7bc77e3efd653bf019ef7b2ab9eca0a833400bcb5e487cc5a626acb112401;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0c34b940c501820ee1731de4afec4cf10d54a6b0f064c97093921fbf078648c63201c362e4bf02de9d407f5f529d96083a18b6198bd62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc42a65c36223dd74838be6acaad8e90268360c02abac8130b0b034e8c05acff6c4641cce40e92951c2de6373e6ec5352883ff31c811b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he00fee36de6e83bb8f9edf0c10cd1c0b764b2e9314e24064cb1f78c32a62a6e9473cc76804b86e4747403fd91dee63b5888d7e8bb94eb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f81bfa1f1985a8efc78b19739cd456bd06759ac1b43c059b87e499b789bc44faf6becadd60d094b5111ca019ff50234f2fff7999d9e3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ef6478d83303efc7d726fc02d7e393917b1598a285551002b472b5de4dedbe3a0af9507986dcfed3d05558418c1762bc002e3218f0acf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b6b4b48d7a166717ac62c244df28e86e327936d8805420e7057b4f951575f15b4754ed1815e61e1d02a5e44e0716615cf6d7123e1fe39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc030be1683dd130ba1ccc58a16b8566ee5e7d022eb7fd6465c32134dd361f539157d53faa1fc6d20da1043a381f8fa1b72850f36cf1a55;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d507498e0e4da6efcf56eb0e301c5b2e7eadf27a9708e61919e5683f32b64b3835e5aa231aac31caff85c6a9710c42392672fb2cee233;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125428a7782a6a281c2057c448a642eb05a5d9927c473f0be137861339c2945b91d5e7d92ddc32d9b5c5a76f4e36b926b5d65b1209ffb51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h955c03ccd35ac33433c27bc3e70b3315e59e9964b4442cac3814c11c68d776be932be0238353cb19288fbf388b5675d979af7c216a1fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d656fac59b08f822f591d08d751034113936cc53f2ee3c9cb74e17333252d78e181da849fba3d0956f360360cba251bb09256572dce96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87a59a481ac823805fdf4cd7ea6cbe8f7a928a6dfcbfa3daed46dd8e72a483eb16bfacd3b1f50bad741e6ad8883afcc637b030c7ef1d94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155e767615e03ef9e66c4f3ae478a3774401dd4dc4489cf37031207542b0ebdf6825f36823cabd73f9e49fb65ac2722cb6fbd38c2d90405;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha83576cc44359637736df8c54013f1e248b04a1be4247f491abf932740406490909204926589ed560897266e285dacff87df4950dfbc15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b4dd9a1fb89fbfbc897cad8f112c713d555f08d0271d1eb276c4211b3a3a6c2748563c9bc24f194433601e64d1c22d328202c79c89b3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9daeca1a30779efb22221c09c85c98a3f9cd2c24e2b50e715102139e64c9701670b90aed574732c4c156beda3d505dda0983e084efcd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe90ea070382295382dda60d44e0157459df5a28c5a146b77017beea3b4c2a6ffee30bdaf69e581dc8f9c31f09da9170f81498f48a0532;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc85998d731870466c93bd5cbffc5b4fcc2136ad95b65724a06c065c6ac0ee1b17966794f3a856030d847cb5a8e41668dd284a837e2f98f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d305a443ea11805a9ec06a2a8062d057992b257b93c6015b90ea3eb712ed74ddf7e1c830ea4f17762dd0f8f54d7231ecb306d2d4b55f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78d57ace79d0a4decae92eaea50b234a2ba63ecdce0c663b360ff525c00ec81eab4b27a7ec11cececb4ff2b90b6f639911e72e7bddc6b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5dce99c9426524c521fdcded22d341db812ae3fb32a8a5df36a66ec3b99770dd54dda4d5c51d601ead5abd0b4aea29a2d4986322ffa1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92cff618481bbeaff4c2f39c1f002ef8f0190ae8dfa57c427f392a4a4815a058d24d7361aea03465701173d36ac50eb00b628a2f2d97b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad611c730b80a8b06e1ce3d7b828d64f67a370de8dec3d87d8c38746b3a4624a6baec0f4aed5b5fee457ac1daf5b134b9d9a0eabed496c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2d999dc2bbf5d88dcb0698640e99216e58383430f3cf9c4cd078c12b1dc72eff930d82b15bf845f6f9038be978804b7bb94e114886f6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14af70bcaa88a46a996f4a04b48f53dcebd491f7f2131b2976e7c56b5a3d8f17cc243d6c1f54672025a6f2cb5b14cea975734f24d5d8b77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157c4457a8c0d5e090d1fa8994ba54ea23c672e4dada6e2071b9621e06054371ac35f2feb807c86c07ad634179f9e7b0bd43608f3e0bd06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24f4d7569f014cd84a48f5881ab11ac8b3970a262c63d76421a466847272f266ab16f6c85e94beea0980a32a89432e5f6d04092ce6819a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1499577089c4bd4c2c3e599e4a1a94ed29da81fb0ccb7c51cac7a74886dc1312bf7cea2cae5df04c313d360455bbadec5f8909247f69f2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc231946d59d9912b6ba93f43ef9c98664b24b321f9f42eb7e3c9f74cb25cf835288b5b7a4378315c0ce4638565b3790602a15453f27b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f4e2a01c86c9a93a6392dec2c6b41c994eb01259b00f99762b7d5ad630938588567fb3474f8b4e417204e478b6083ff78f20ba74caff2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c176efa9667850b84928faf8938952c1a1cca71765cdb7f439975e2190ebeebabb113275239d5b6792c304a4faaa4547ca8d9e234c871;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d4e9f7ec491dee97432e1d6aab9dba6f41abd3ded4268d6282aa80e96fadf05495e9236cc6fa2e3604ea4a31c83e8624f55474b852225;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3cbc61ecc07cbf426dd9f4e4e986d5cdf2d2f06819953e3fab2ce8e16b67aceb51d805c43775489a179764754bfae2418bc9ce1b6982f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee333daf19becb7ca08861ba8100768190e612ef54eaad4d461fe0b8b3840f80131bd42240bf071df240f09bdd9f15a6c5745b5e977259;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0ba61ed07b5621b0277ac0841b3f917a446a2d7bef34178171bb3c5b9756e2039d7c096824f797186e03d193a08d2b843f1923926a476;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19aa1a794eb44ad1cc862aebd4780ef2508d5b9284506bd57062e9743fd80d1bed4c93cae1718866cb7a79b36e9ca4b359322f1468b5fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e339b4fd491acee10aa5e9e94770362e740862bd1e31275447d96b1d98959f755a39330d273bdbef96944fbbed97a58abb1dfdf594490;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1ba366e6ea2db4877e06c22f196048510107557bfce145d92c47aeb33cb688cba10ad34ed72f32ed2d4c167dee79394a21ccb2b21dfaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heffdf99fa82c6a8f278fb823278913569db695fffc7f5a01a0cd819dbcd5e57afaa80eef387dec8f12ca73acd2da146e623d834a65af39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5f3fab061ae6e3e15c2d4be740c47c3cc274bf15d6f7925029848c87db130d2d7f14dc5d0a966e11b0ac9a7388869883df18f9adea2c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4469889123ce6cffb791f62aae8c547dc1a9ec2408746c10be00eb1cd8c06fe7c88fbf7d6de027580d4dd5cda39b0361915dccdae2d7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f78a9c226420a7d98e4e7329462bb367edbbbae07a83e35dab680d0064bda03dc70c638bcde89b0f4fdd8d45456fdce2b6134a578e064;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c2a330b7a4c88bfadd8f39d10d95fa6ef65210edfaea07a4e6969fc288f1572463d127ad9431afb383bd9e6b99a2b6fc1b395eaf2a5af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h394628baab995e145357bc19ae3b004914ba5e38036cc3a75d956971c87658e103af424572f47b8a9a99074baad2080a356e7659990333;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82dbce0c9ff27d89e9ce744eaa4cda9b4fa9f5868a7f62f236100d0354db1970a3b3e0da861c9dc9fdacd47c0987d1c4d5dbd83e93f241;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105e28e0d4697decd885fd863047910cf903fd538a8f6c14ac18cfe33f993b5758bdb4de76d13469403e0ce084884893fc98c3ad17b26b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ddac538ad4177d8748e8a173af1e1238baf2b9ebc9b3bfce97bd3ab572906825d314736c9b375ccdbaec320814d2323d4c3beb6093719;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dacde4f09049c46f04fd633693e5071df019d5650501a2305d636350b95af8e51bc6301732c595f099ed8434e95762d90fad01022d7a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31ffa07648eb26039e19d04cdb9b64a406f0cb71d13a3db6459bac60d327da030d92473a729414ce5fbc12f5697b7cedc00a885679ead7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eed9736b1979c53a283093c513e3d26c2cbdbaffc225f91b5f680457bd8ea5f27b38a964c9c0e199740249e6227f1789f4be2dbf54dde0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d33211a2cc92df2782719c313013fd26b7f654c77d5f1182d58550347952a6ca0a1ef77d1d6963557b66f699e439888b9a161f32e7117;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab8e6550097ea356b8edaae6090b2839e660591b71708d71f63d4a5280107168402b192aa9efb7dfc34624f283af6f1fac06692f31bf02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha002cf9e58e97478652e1fbb5afe3c16410c1634212abd86914fd556bbb5bb1c133bc9d201347a347049347c9da1e1741fe5eef43c78a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3236c07e4146c4a6407507b56338227aa3a774d705236127ba38ae710e577e95376bd91e715833ea605ecf04f94514fa3988587424bfe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3214747891c08a120b2395f55935f7cb78602bd24e36f39a53ec9124ee171586f7ef3923aedc77f483c40df4b4e54bfe56a693cbbfd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c844570c8263d359d6f0c059d28852e7bfb159e1b159e7b286c49d8c3a5da465cef2256901a96cac4005eaa74ceadc073e4b74b0755e36;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134c75f977a6488da15e5215017b92c7bbab7429bb79a89fbb589a4a023969c9ed0cf92c512e3bc362861646a9df71a02436250fd9f1e25;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf24f579b5b676b855cdeb722b48ce66c89d836829baf12bb6107c493d3db003d72e509ae935099995384b1dec7800a0f0f968cdcad9f32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eda0c1f4aaa8f35547fdfe12099507a9bb8eb357f925d9f7bd49a30d80c8cfec18b5940fb19b046a744a38a81fa65d84759eba5a0c60cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6ab08c851b5dc5c8baa318aa6415843ab6503bcdf1d029bd0d95e89e7db31d97e6ce590e5a53919565fad2de6b581c6c1b4c9e4a9a28c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf401066d15f15f5659c65ec33c393469714f152d8fdfe4847da768483439ddb7c98786e5111fc6b1a3106c3432112f358c5611e7a59ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b2e02c26bdda42bab340412633c71f75ad7ef7783dfb3608514b1b4e1fc2bebc136b73579eb5fd443b7ca88fe47996fed0ab59a7fa54a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he878009411da05b79c4e17c119ccb9ef2df3f9f7cdbb9bbba64bdf0b78e364f5509816842eca2cc580e52320eb9d829fd86a591f28e6e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7f3aa022232420c166c56a75baa8ed5621adffd63fa1bce9cf0aaa552dd3b4a69a9a2ac61aa393a32a3bf2ecb3d81ef25f6f74df8ada6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h507c7bb7377b6b2591068e53eccf4959f9c0775acc562e30bc62d1877a3071d8d3e997f7e2c106ee7081af37c3634028e25f95e8f7d40c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd02ef14c2300c9de59f6002d2cfa8f0f8db084d4f2e3f4d50c2bd706b1eb558915b45abc788f83efbc0a10cefe00b0625b32af19c866fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab9096faa604397351f0568e17d86325ff93558e26c246b0b62bac5096f414f7f53728def0da69381f55657d5bcc29542b4e032dae5571;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82866269db38db57e7b2ce3bed796b33a93fc660238fda7954e60e1d5b4bf566f7c6ab23a1d5a42b7970518515334b58ef9a7d3b306bf8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa326a7b9a693a29ef4ad0b92f9ca52d2565148114c17071d506e65e4c54282a74110b418072a8b8f920d680f51e06614cde29cc349510;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39d980edb9b26f62f8e4281432691c9378ca9edb69ac4ca318f502a23dad1b531b34f02a63953c721fe38959b61288543b312bea440c99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f19c8515cd5c544ccc29c6ea69d68badde84cfaa4cf3dd86cd756200aee04e980e0dbd77de7009a565217d7e779265d10ebc60550d33a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a8bb5aef8bcd1756d96183d3a926d7a3aa2e8d926587db95ef1a0fd865c7fdf5451ecf15a303b2251bf506eb8ae4bf7f12d1a85df3027;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7d1bc36b8cae8a8acb728deab187b7ecdd42d4bbdfc794818e0f07043e15ca3d9dfba277936d99b64971cc25a1d45f8903bc2d427b3c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a59b275f1e59decad2cd7610e0b42f3cfefeb5fe8153dc09d958d4047898728b50d3b38c270de9ca8dc3a1a555e47b9b285bf4e0451a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b6a30fa46b8fc415d183768fe67555f944753121140ad08c1652107dcc76825e77eddd7974890a3e5f3906caea352e29e954dff728965;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179b831b306b3baffc4dd080f9a151bdbd4ea76a53f56399bffac3fa998e4b8f688dad904f5f3482520b3d09434f4732dca742c30409231;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22258e3c9144cc36c5d8e4e6180c379fdbf37264c6732f59f7f59f6c505a284ca6946a8a5fea0e249510502a76f1984f96835e568ceac9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad683fa83ffd39d8a153b8f0b816a2e5307422f8b13f7daf62a43d0e93a174fd64e342c37b7862a898bb8872c8b31e646fb4de56c9cfde;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab30b8008f7808fcd9dc9404a98334149fbba7afa8255a60d1e8a2b707105eba9d8bc8bf9eb22dd834117712f3a8de8e881997a84713a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1251579b545997ed18ac74084af03b2c820597f5019054d344cf9219cfc2d9f0657d0c96d6d7cf1fa26909fac785b1776588ccdab59ffe0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cb123ebd19c53b7e8498deff61652ab3c2846f472fae491e43c3849db59ec32f82398427c8f947034bb7fbfb615aaa22b4464cbcba29e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7c47ee1d7cb468641b3c1ac54700b358894b3924bdf502cb0e4172cd97fde96a9dbdebdc70cf883ecccf6e6f59bb1bbb1fb4bd52c0a04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1565beb7c8ea0693afd85bd05637fc30eeeca81dcf1465479ebc72b4b688c37d0bbdd8763f1b51b93f51d70dcab090788940e9226e2d056;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54665d8153615e30307175065724e87a2d6e112f23d030b506e1e930627aa2ba7ef403aee63976b816c08db3eea3ac2ab1e02500b5ddd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4017534520fe04e49af2e1b25dbcd0520b9dfc7354052d6318ac74ccabb9f9bbf832b665dc0efb3626ba5d8ee4a0b53f63f06afdf82837;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d74b7b56acd49028a932662ee8dcdb85eebe9ba66baed85be7e9c31ed2e2fea62cc418b17a89d798c3a494d02784cdca3fa88cd17eb70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ad67caf44fa794eb8617f9d0be80dd94fb6df1a6d6bc95b4d96ab16497c7e0a9d3b17b2b8c10c841d913f660aea97cfd16f7b288ee13b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6e110dceb7737b47e9812fbf2255945da1243ca3ef8865ad9e71dda1b15a874236d03d3ee35d27e78e03e5bfdc099d810dcdad513cc67;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1443896df6be23bca8ee908d7d3a21d7832f34ac96772684f1741d6776ea4e0b474ac45e50df35a865035cc6f7ba6da0b7c7ab0b6df9a16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h340c1107bf52f32aaa435a29988b2b88e907774d8011891859343721182805fff60bdd82ba33d7da8ec7b0105373e77280b47ad3ee2f97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h252a6fd3c6a287b9cab9b356d32e57b0b839bc9296d04db2fe9e2b2886d7b90f654dcd91132de87a5844e91c2d290a20aea07eb33dd6f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19df0fe0986e176e5695c99fa7df932657828d0f2be9047ba544bed7c51dd19c50dbb2bdd21e24bfee8d5919ee754a4c729043aca34eb2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11eab25192f00fe16cde542dd84482f5346390c3ce99293f93a2006e4d466200053ade796b83d7de725ebce62e8ffae9519ca0f3fa812da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h400d5938e8fc60b2c8dacf27ea3e9561a15c3b99b93a337eae0b92a4f8454e2ce507e0f99867fc268df8012042e19f995911220818495f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f6ff3d248c3649d7bd21728ad48b621cede10e6b0ba3b152cffbc458ad9458c876067598a4411e97a91d5de0ab5993afc0ece9ad9f8c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bc41960e272aa9cc76d15f13b3bca607c004637bc865daf5b88b79b8cb0d68248d1068b277435a92db76cddf8d9e144b3ec5da9cac4f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e287f3de0a0a28f8200e16b1d38207fcaf06575e3a5507109ab654b03e3b1a9b0a010e2bc77bc152e8e4b24bd7ecc008613f8a1b8c26d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9bc3a39ff0fd5ea4c7577a368ff8b2b4b00cca9deb6050c8e3b1817e40cdd750e07b7db603157e27cc82e6a9a0d058afe80c352e8dc182;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4584d305cba24a1554dd8f697f49968a1e67b23bbb04feedf5b7eac6cef98e07e2e3758a21c511e1c931cf349f37bbf121bce2f29903;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf585264e07e16dd7b2dcc58b9d3b3f267b5c41b8852aa3f9fac846ae0a8298ae4246838651bb3bb038612c03045365f77862ea309df97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc91f81980f1b207dbf0ed0fbaf4d302852212b08af272150c687efccb82176db69067be620f86320da37a9986ab2bf8484c3e7e9a14494;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1392270d49d975cc908ce13c6fbd47de1f79d8659e25e3c1f3bac28225ca018d23fee7dc838bd0f127059fb7812a81d45f020bbab3fea17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b57e3940236d7374e5c7fdc1c5ef0b8baae7837db6fb21d34078de263695f61e9a2452dac3d57ac48e351f98f6b1e3e9bd9f1e549d2a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eb784da263fec68cf74f175a07ed11cd76a4763ae47d223eeff26f3af1a6d721f20e5f909aa154462c8e9cd6e0e25f7d42f64835c30bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107a3bf35757de3f96a6ebd22382c2d80b0ae5d0210cd7dc06114b65e7d20c171a1e83226cdf7c66b577231c3fbadce4ac7720d111b4b6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h869a4e0256b653f6f7e2598344572efc97453ddebc7f6e4deef5754a9bb52e0d0c0ea19e5c2b14857f94669bae7a44db217176f50ad4b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h704f98548f6ad63330b1ea159589e5e748c7764116f0f7f2d000358e2754549630f21bfa19cbfd25a515560cbcac312ff23430fe023df3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2facfe3ef063c75a3212a7ef9b1d46b2352649779b478b6e45c7edc65ec357d1e41d9d09ff9b1ec70039db048c7d29fc2e48ecc7513584;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107631e6d06db2132572c8c43d0f332409bf47b190e9dbf49230c0bf8937cf42abb9f631a7b65fb61d2f92cc238c010bee366d46f3cc1a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3c7e066958b6ecaa22694a878c8343c6bedef81a965ca792af51a21b516a6213497ac01491628816482d30f08fcf09494d3d7398fc138;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h600cdc2aeb094d22da405983e457b5ad450b93a7c87a42fc988c61773332ac895c970f88b229f25bdb6ad7d82efa5b64f42cb2e3356e6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cdd7c1eb418c22d063c93954cd888fdc3318c6bd87f50365da6f0ecfe8c0099284a3faaec9e7db578560be5863cdd140ec7179472316e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12688612b9c377b4ee4bd9be8c467d7b5415a81f48024df4b5ff6a8def9c3d560610519ffade25c4284e94608a6431c3703fea426552668;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcee84c649ac774c44f78d8c9ac01552be4e0361ca2e9536f09162467dd6fc5245194f0ebaf777fa175f1123d9b0bf2b346c79d65da7ec1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e22f8a7d11e6083db00e3b7470946128b84d0a74364dd493f8a9d4c585813618919b5c551316e71de1e7e4edcbc818f1a39e14c1fe2e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfc994a0a1756623ac491eb64caf23e326d14e691f328e3ce3f2159d246d58e61ea1e9d01fab0c5d6f2d269db5f452496c033599a192f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5bb2f01ba362f9a2c923f2424af7fad47f59e37db8c7eb9faef61766d9cfd4031edce5f4634164f04c0d9b0bd0e15c5281acb45186032;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6204074ac189244f617b0661eb54c746d2fc03fbf3c482558c33373220a68493cb2570e027a6729e4de474cc688178d3a72a5644c80b18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3da8c7f090bbc53904fa8935c2f912cfdf96becd992831a2196d50c84aed563a7509326a206ba4b10aadccb65eddb01727185e71bc888;
        #1
        $finish();
    end
endmodule
