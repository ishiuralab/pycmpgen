module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [15:0] src17;
    reg [14:0] src18;
    reg [13:0] src19;
    reg [12:0] src20;
    reg [11:0] src21;
    reg [10:0] src22;
    reg [9:0] src23;
    reg [8:0] src24;
    reg [7:0] src25;
    reg [6:0] src26;
    reg [5:0] src27;
    reg [4:0] src28;
    reg [3:0] src29;
    reg [2:0] src30;
    reg [1:0] src31;
    reg [0:0] src32;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3])<<29) + ((src30[0] + src30[1] + src30[2])<<30) + ((src31[0] + src31[1])<<31) + ((src32[0])<<32);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183219e0b87da425b7f528d0bd13577b2270de26844d9b494661073d4f7b29d85f9f5297;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h167fcb3a36a23a6a91b366b6ce1e6fa69a18558dd8f3f68034950b624d489dbc7c756bd03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20f106493c75a800edd55697d062c0d17425330b2a827a851b98e60c5e1a5172b2dd7d11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d7a0f235fe15a7536c9929ef9fbf3edb9039d09cb32ca3751d46e498ba4364f4a2333f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189fcba3a9f0a58caea36aee56c59749bfe939a52257a731cce6eb0f4cfb35f7dd5c7d853;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cd0e1512346d43353afb555846d2bfa1dd9d713267e913ceeea61331a02cf68cc1d8fab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182d2af6e1f178fd8ecef93149ef07b4c02ea3066b2059cf9e46324e8c1b4d55f33b8206c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9651c1645a14296ce13d48466cca15184f4f9508425a0046714ada18683c1c41ae5c057;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e2d34444d9ad25fa323f2def6ff79a89e0054b8c708e09942445c54ee5205d08b9ccceb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53f3ff59572ee54c8d49295596a4862f05eed1d3907db94eb37162de081d3f117a5feefc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ad2d2062092299872380ba28082719f170328723b1127ea6194da607fc1c58e63f59e7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb065316d7127254b2f16836efde34597aa2440cdf75697f7857829ecee8caf8ddb172430;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e9310ecf04f916503897cb01c6ed4c39e49af9d702fb64701a34e77d31c663dd06d44ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f91b3c46537fee7aa297de905123335f8e30970f6d7c559695ddfae6409dc236e1e3623;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea17c256b49b2bd37767a3dc13bdff4a317ab7d182a18902282b8d9479390ba627b82479;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfdfd69fd50bd073c53f6f5c82894ca9c56bbad0e58bd6b481a50e32cf056ad9303c8575;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72bf6d2ccd22ffefadde44cceb9252bd322cb868caccb0d085c16a5c3adaaeeb3513519d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haea523c4a36521a22c65a7437d5cc723664abc3e32f771fd9516c1175e42a334bcfc69b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0e57b8b89f0b7a29ec8e645ba3e93d56cadc0b2619a469554b73358a2c70c7c48a67093;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a661343513825f1deecf1230000da8462bd1b5c6cdf957a7507cbf00d31c3653a8114dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bf5dff0e51b47b78ece2b92a0a743689e785d155856cc3986cdfcec3d9f66445e5dbcf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef20d659ee6db066cb4baaccf882c647bdf0d775d8f2369a51cdb3e28d5efbacfb0d6170;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1951dcd365e083c9c5ded383767deaf0eb9820ca8099f003715c3773240225fbf6291fb0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50ca8f52dde1f957f24e446d4d1f582df36d8074c9b9874aac0ab0eb1a43e884261a8e85;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ca27970ccedd845c734abda39d0d66bb944d930418277e6b43a5a4c8445a488066d1a4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43dde6f528366969ff23ce72d60af8b0d291d21c025a5333736fc3b3ddee49d28f268576;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe26ba5a8a0efc09c5087c379847b146980f634327cb5f73378894e309760cde8c5ffe78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166b32353ecf143f32e517c8cb1d6aab7ba8bba6c4bc6f726120a5de05fa7fc5ea2950e9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158d667eeeb2e84ab1a14413d609cd6ebd7b67cb1e89d7d82a3f2dab4b62b078c919e9d4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21efcaf383da69282f1691f32371c0b6392d7144521339940af96d927bada0c1a3e27e89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173c95e15ce646b8b24184fb40a3cde6d216cfde7e43af5e61c2cbed266b6178c76cd7a78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103a1a5acdd86aa5cb336971de17dad4e36908d45328b83004d03d771edc4eb1809e15088;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ae417fc75d96a9ba18bae7396f4e2a7502c38297abe60364eea56d6bd39fde1fec3bb01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81a71998f883ad98be97aaf3e5123c01e5aa07aff46014aeb2cacabf0335adc98008a65a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118d0c7f083e9c48d6f3f74676ab1e94853d234b9ad3370085668e2d79f9d90a8b929bf9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd70664d15ea01b0db667e1fca7693a9299ee9bc19dbd2f18fc57f29c3e728a2db343f798;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fad7e1bad338acce49f6d18eee53f5216508de56cc37227cd55b993be1ad23623310162;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8470fc920b38d2d3c87d554d8b0fad395b156af499a7dccc0d9ccd68068ee425e62af4a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151b362eb2258ffdbeca54d2fd784acace87cda8006bc0d2009e1d97132b3a7330cbf7e46;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ceafa0d13569096e2a51359c1ab2d24355f4b8128ff4be691de93fb3acad20e38306863;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc13c11d0ca44776a540c53e0ee7509747ade49e5cd2fae041cb5e55486968edd24a1afc3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f64e50079d9b0814923df1accd92df39619a3a99f59321b2c7b0f84c7aa9980ff02b313;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae22c0a3e2ba1f31265cf7cf79057b48130c435f10d95ef5e071dbc2257521630de1e3e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6f4ee300b0b81f9c9c858228bdddc3fbfb965314f2a0ce23032ae0b70e64ed0674b4f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1806e332c32d119e9d17494bbd56bd8990d7b122370cd7c89ff364b5cc6ec0efcd375a2a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131cc993fac95e3761f05e9c7debb75205621734bd881bcf5bff333ca8f911a92b4159b42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9cbdac27a6e26a0f59215fc59c5a307e6951ffb5da4c6ae0f7d8976c37014c4f5879232;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbcd29817b777feba1592a00e296ed315eecd051fd428a0823b12bfa95d0f9d95bab1a2d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fcc0ec01d723ee8edd21c9474e09014799437c55b164c747d80d7960375d891f2e6dd27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199fa0e8b16d7b0be66d8e51ef184e167303945b13069f6c16f13ed58e55f9ee295518dac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc838faa3d8d3d1bae998bebca790527391071b3fa78f03cc0ae5ec745b065b20b18fdab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4a3a4fcbb8bb9a2df4783702f7e7ad9c01c7fe8fb94cbd067f2e8bd80b056968a435919;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da132fd8eb7e6135160750e307253968805d0b0b09270df4c6eda886abd63db1d9cbb46b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a9627e36a116d170a41e51aa03e29c73caca73e127b2579f98257a5dc5d8d36573a90de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c471bfb347380342a3bc5880a88fce0d1e0ffa256d05beb406a7b533f195c2cc28c7c7d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37f814c252d708ba9b7c7450f2c8536d4da8b965f1a3d01379391970f6d52a9a7baf4c4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8ce6df88e22601e5946791dbc8dd95242fa1a439d2019ff3151b884585ee52080e8592ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fde5be4d6a1c600d6d1bf51d83c1d7484df7e98c2d678f78e27b68af9d98e293df1d67e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43fb5ffbc1e541890496ed46553f041947f227f6d345dd1a61f101e5d5fcf91f3cd9d5aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1548b121df513ec87ce2aec3b11ba8de32f44d38845588668ddda23b27fa8bc3148e3fb5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h355c6e36506bf4de5d7eb5a6a45d19f017cc7641cde5a6e2123bb5d16639338f1a736599;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8aa891baa0c9e6fb1ac93dbfea648f784a543c1a3deb433169a5389c64665792bb152017;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bec02b0a6f845e9938083cac53edfc1c09eb1c2493e3dd0841280fe222a1b43a0f047e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a0d62cf9f0a799434d0b9c939f98f12a0a2d5f27667c5c401d438ce1f1625d01cf0da80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0d1027f7aaa4cf2222c3b62f8be61c79158447c43ce6f430b50b90e640ddbbf4d610d10;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14eb066a661e859b3c73ca3c4b22c1edc14db22d1549d67d5c25640d77300b762b71a9565;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3e3a3a1ed341576550267c4e697c0c644fe258997357dc563c898d60e648fdd9a4fb499;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc05f898d43ea5a9df136c66bbb7500c631623554388f6cb19c74064e4a0e413b4e82e3b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a569fc8257645ff9807c448dfc9f7c6b51c6376a3e27d3ae7dc87d841e64fc32f265dd07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199ca3ee4746a97cd84612f89004412f3705fa282e16c44a105ad37208a899e08d35c8e75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ba57df44f5d5b13728931ad334673d361a2506a772100f7d49e261ee02ee4e60a56c32f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c35a5683dc5476712f3b4d2996933873961596d4411ade946b133b592a75f299a2ac1b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4f15ddf89ee20d0c3ffcc86c07916bdea925d18915d3e66b474d8e6a4ba2d5fe7bbb9b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d7938487f70da36dd0b91aeee0878b2d356957857ff24587886e59c48ab12977febc770;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd210cd54461d2f8b58edb7b5c4b95c585fbb8fc8e0bd3044fa51f18f529dc46c15ad340a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e62b0ff8b389356fb57086cc0de7484f767f85f1309ed46e1cb4e8640a89f775b2165e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6da828a91ace2193969f2773b2c364acf7a83a38584f1b267679543f7164888bfd0444e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dae4cd45b39cc7ba03cfc468cbf0d3b02b65a949d97df39f9cfdc5d29d5e09688c64ddc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d7f967550f6e8c8cada9dd6329968a4a6bd8bedae8c63d17d30a99cac80c8bec60f1716;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e843199348745f4bbb7a9f4e9387ce4bcee2f5f2bfb59216288f952ddb2abb96c026813e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1795dad364956d3bbe5135d11a10c7530ec099670f4ffd61b9e2e61ed2e46956cc3f4e28b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89a40b9abb46f5a80ac530d98bd03c7ab74e45dcddc28196950ba229b139e7ce97b967dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hddd07be5005997fdcb1118bb7dbe1581189fe71a5697fc9af693984ebfe52fe5d66597fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6da17d364f1ce75ecc842bf566bbb32cf97237bd3fff8544e62ce30b92c30f5b4a6dad13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3bdd06824d85438c930358e439dd5e437adf7bce91341aabf62cf408161067a117a64e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155283a3415f88f2eb298983105a1e0689aa84cadd248b0bd8021d695035eeae9cab2aa38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0f74c06b46e81a5669410462c0412d09d15cda8be490b63c834e3a2e5bb1764dfd60d4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12040c0a9191ff6a76b282509f975c463b292970edd30d6c2bb7c4f1f14b6b2ae5c420a87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1722ac2243c5319b18d04dadf96045e317368a4984b95f3cfe784124a7da062b7e26cfa05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0842ec219cc3533eeddc951bc51f89178f8e30ea3c84f52fc1cdde779180d8fa72b10f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbadfcc774bb1a8d852cc300c150e7c1543195e2aff4769b6e69702fdd0a016c0f89a8d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h682e62d1c7dcf5d6cd057906fb516ee7c8c23fdbc2c082493a3316b1bdceea94cc060243;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d16a9bc0a1e7a02abb444b74df674553879c4912724cef4c973179269673cd14c8dc733a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149fa5e39509014266903836b3b34e6b1d6b05db78e47b11c3ec2919e442e9d996a4ad5e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e34c2734cded9d321312ffe1dc6f97283eb926ab48e728ffb41e7da71fb0201230eee13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faba4634638c8457755754eae333bcd8b6f46e490b28817db50ff1ec20f19521dbf05cea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c9b4fd81ea757810ac8121fe72ff8cecd3b3342ab39e764cbc365e1cd0308b66013a0bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e21468b8b61628cbf9b184232aa0017b1d10b28e709a9f11644234ac5ee44a0f178a0ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f54ee2b87017799fa007bab358aed7256308026703fff475714f59e69aebda45cf37338;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cad1306af9f00d2a1e0f3973009ae2dff5ab997597da62b5cb254d5db7fbe376c80e8c88;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cc24f324291d02305c5baf490e77f665cf0a3d20514313dd4b7d2682428bacfcc879220;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c404ce453a3b721b31a7d0820fb5a9f7ab6d1621fa9aa7309d27bb3292198bb2b0bd735;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a931cff98dfe25ab118ee55e6574b737a35f00d22b2315c04b30b0bbd6db7d94a9b5e96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h148c3c5a1359c144347993ef8580ec0edd0fcddb9e23ef14861f73c88dfdd0984d60d92e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184e4ad3efd1d42e0c730497fbfba1fe63e3d6ff6979074f2a492c1e323076925da30f4ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbc14a06e9fa1add3112f35b7873f1afd61bb358e0c5d5098a48e928397bb858fd305cea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cdea748b5b3d0f17a3dfaf5a6e63242474b9b6f1084ffe67bd89ec3e4a6cc3fd174b5e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19cbcb9e35de9e43723bef33989f70ca322ca34361a54796baf16f9c1db39e92ec6309900;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f01719b498984c480e58b633c3385a5fa1e2b612cea217a518961feb192c2a4e487c1de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af1069bd2e2e9300ea290b895a8bb4677d38efed4b076675ab8c5876ed5b27fe8cf7a01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae23338f4394e104ae25cc482ba7354f870680665f26ae5e638d29827f60265b25143fef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7e604456f991b4e95ed68bdcb5311417d135098ac36f6010bc183e3a16290fac8c133a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d32ea95382ab117937b24e06c3c2698d6399b225a3db770b5ba5f1b49e2bbf69b0919a0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1a10ef0a3adb504e06fad33861a50a6581fab9efd18415d48e8e954b9f94ab44167fdea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4ef5132583869244925eb650b4f510c849bb679c0aae30bf43283ec03ed0c69569e45a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e6df2e0cb5ec2fed5ce811a748cc74f04a654a9b3334da7a5cf25a7b2fe06b56d363f34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f2844ec3b1d75dcaf59e29d87f116b0fd3c392fb4bc76b84af36eb7ac41fb10621ee926;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170d85b014234ab3f18f335dee68bb38b1345bb082feae3a42d1e522c1ce0ccbf51c4cac3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11adce90216e1b1bf7215c740f8c177a3699d5fe36d7b3ba4c5151ec09bc5126b262fe8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c117cac76521fee9e9a90eabd77955b9e341797d9217be06cd17e38f71a3531878d83eb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8f92cba1a78e96a4caf2daf4f7c35565b5587eff927ce05d5f28240ef8b6475fa8de831;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb7499e53ae8f78b3953b2dabccd791ac5792e9dbd4c72259da9d296d22d0c6b7cda248;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111fc47b86a23259e3caba27a37f0ccbb92969437758b0f5c0136537864a24f30572a5bbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h489fb03998cd6f6224cdb1c4cbf41e478d9d4d1cdccd20fa75f6db94f79e1d96c95fa163;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa6e1ab0dbc14fbdb445cd8e5b42619ccb01e6aa1a6f4955381008840c5a89863f3074a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab67a889db7c160b0a649e8f53afc35b2d17a586c27f164b25dc2b42a6f1fd22bbc7c32c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d30fcecdbae6c2e9145b442b3bcb9c483b7551971cb7f8c3e39a150afacb75eb43337a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10028b07d9f1a31dd3f9334d08904121e52fbe3231c29edd20d3d4c67fd0855462b1d8ea7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a47e61ea4b43c843b3aec6907c8b3442213da213b166f9f33ab7efc825ce11a0b290139;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f1bba265eaf62dbfb0162477a993f5316f1ad8f191a4c32da925cb028bcd6930e858841;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa3906531ebcc37d08b7a83152f15a1de7f4ac50e0edfc3c43ce080a57cfeecb34150af6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e47e838725b622402dbc8c7ce2b582f7ccfe20972ea352712ee683256ebeebd386a7b04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51f9dba3a8449816a19a2a8e1c4dde95fa82a43e71f24a72d933c21607dfcf994e31209c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153fed1b693ada0e6669a22f4031de44eea0c111b7e5f9dda6258f688d88513fe12ae3750;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f664243596f31c9a1590e5aa8b946b0684888a99a35970e35e3160e47ec8956530b0f65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1840bfcfcd3d8fad96be08f9eb02f1922f390d48fff2509a2bada2f158c746f641f1f2c1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c0aa70e88457ccfa69165b92486aeab3665b3f58c6116f5d7f7d9d6c9c5db722af9c670;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1019ae35a43904e220ea09a2fe616308f56127c4fb6aefd158bdf6902b89bfcd45b40cc7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a7ea0a5d9408b50f2be13918847e7c17212dd2289ffc2ff2a2a2b672f60f64f880d91ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1692324ae16983f7e730ccfdc0e75a03630c5e57339d8b341fbbf064bcfc0727c3e3b48d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1014aa097fd5311d970f92d923db8f50a3896e02395f7c109684d6f8ea1ab1b27149688a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6c587196a75468d8f20330b0892c52c27f7ff8325d0be5dc048082bb24994e5a98c57c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a360758283a36ffe026f7e20ba117712aa2871716f7f939f3a8e94798facb97181889a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b7f706d0c77fbe8f36707d2c17c5cfe5fd9a50115ba3448e306cd70b44044adabe5c903;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha73edf859a2b67802971053d858b761e3726c61fdc1b18314b750fbc1516b07a5e7f3052;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd74c371eab1de11cd58031cd54fa6c4230dd08cbd43370fc8e5d50b070c73a63563b01d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63cee338a991b18dddfc64a94c5b94318e877eecd2b679c486a905dd09c404cd6b3715f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa3a3ad9025547f720964c9a5d3a5d7862fcbc389795219153ed5210f63846c41b3f5b57;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b07d602906b8a024da686599a6898be307d43b2ebecf41f8f9d7fdd78c14a536a7d491f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138fb387ae48776fc2ebf7219c81340ab605569df803d56fb2d7dcb5be3078a7357201936;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5b0196e06ca489a4dba2c395c46e24c42f5dca2a1ec286cb4928bf31eb012851308e1e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1581972ff3398e0ea09ce9829d8d3baa7ce85e076201315cd021ac1273b77101a155ab5c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165153564c0b6f9e6d9eb99e35361193491b1f3d0d02d5f2a70c5c937a9f00ea5c799801f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14019a0b016362de860ef9b5162bea2f68e9b9d1d864981eca59e1665901508c13164968;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbff1329a7e7d1c771e05edbc5d368a13a19ae0581fde1525b3de0185788fbae7b9402725;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be917b4eb60cd9bbdf5ed70caa23e125a9a0b6595feb65844ca1fd59db2171b8b7c85e40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18fa5f05c7d5e248d99c4403f5bdc8f1020c44f34ca6c6deaa30e96983373bffe7db269dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d680e8e4164263c094520752f80bbd9bba71436f817e89bc6957e533f81fa1f302fe6e79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3f5d245fab65a9c530d8e55b26a36f4da7f6630c6ba791661a0294d5906a8f0a5c20dd0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8ff1d39c15d4e00c709701c1a9ba543445f5001efd56945644d6ccb74b6de490b6e0cec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15526f2649f30b321199d16570428618647a2eed3f7e9b70238cefa77da88b28c3d66d270;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c086c4b457ca77ab15aa0ebf3dbfa34a934718b1fac85df94f6686dc1aaee91949c133f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h952c6342fdf8b5eff0dd221a3927ba8b5365bdc32d37804d5b94b90b1c4d588f3686701a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbae43a39139d3d8910d82d94997622a6e5b9d473d7dcdacfcdce3098ebbb85a2ef70408;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1540ffa29035d23b851b49b088bc38abbbf904a56d67c806d0501c4c297de844a0432cd86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h878fecee8c9cbf28b47ff85333c1bfc5eaa0d1c7818dcc147a926557fea8743a3dba2c16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db9ada40bc5fede41baf89aa6171cfaa749065de2f8e35f2f58b273f9af70016b1cb0fa2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habfd020136239c72330e770f4305211f9779b13690806b3d65b8ba8217f29db4d42bfc6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152ce7c42bd1935fbe3c0f6dbfdf50cc12db829761f6f7cf83ce9b04498e5b5c3cb2d8403;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164355680dc95117dd330702a6b16ecd5093bf35a8832b6e41cf67a1e94b033c79431b700;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bb226b217457b4044fe64e5581239134fdec4d3b6b5321b2f49e62b41873b864f44af3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8d54622b271fb3d1882545a2e6e15965395e6a09a848123ccae9ce74971b72a33c46c83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f0a6628e32607bbe9252e9bef6cdaa797602f43394e66cac0661a4297279d6f95da4cad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d554986c12c2f284767af5552e91372ef3715a8ceb83590e1f1e2a1bcecfa4619d7c2c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63c935615ed9555ea078e852079c8bed43fd3eca62ec75ab9b235fad9a0de5d741b577d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff4a87a2816e1c18c3886f6f1781a6fc4b3cacec4b715aa4c47acbb0d1b6c2b3a06dd77c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101f8bd50c8e6012abf56d6d6b738e15d5db4d614e2b5a0270959460eafcbcb99c6d8657e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha50f7c4a4d737d61007594242857beb59cb4c26b2b4d2b9b542c47842dcf8bb9bf4823a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1482b9ef2cd0bcf743bbe4a9c4d65d208b35852dde13b54fbf728dbb2f96b71a3cabae51c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf003374b323d1979e6b7eddd5483977a8d8659feb59668e845db30cf70a549f6b9d35098;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73b32d3bac2633b3ffc953ddd95ecd7584fcbee0f63d2d1e006e0d40cf4c64417e1bd38b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1320ef119b2ae78e210103df37151e393d586e8ab5e5fd5307448781becc8d21125b75f9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14afad756a22870d4c3c66a4d492ec8b71640cf46e21accbcd5c0b4b31fcecf312165ab81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c7db113341da294029ebb81518648d1acf8a6dfc8e8a6b7896350fb7f50b1abef5188db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7ff9b676b466c25a58fc8a4d33642388792e8e88bcd98b070e6d685e1b746888ae7714c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heccb204a2b51323fba1a8c8ebd4877d5e121714a223cd3b49e395520a50dc987b97be548;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he51d5ab98a47247bb1dc162f39fe192ed1fe58603c578604e84d3aac558def3f34092201;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3d356cc78ffe3e2ec7abe69468a858b424ea04cc3abf2410dc7c5a328af529895382af3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14adc23ca7fa1d79ebf25de9226a25125e506cf8172fe09966b75cc46104124a9215de8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15eb6cc3f27fddd0e9339a3cbb7298b0b778440ffb520030781a8d3bb49ac742c704b059b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf19ad3c568bea5cdc5b737b86d2fbea936ae4f39fbda182555765ab0b503ab85a58fc7f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1253950010bd2b4f4c0534d5b3776333992bd0eca8e97758deb3ede023a6c63f85dbf28f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d13d93298aa52252914dee0335f401d12f301fdd3928098831a3952eca798bae5ac2b50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b223a6567bf9a30f901f288b8ac2e4722cf10525f8ed238df3c54807cea107b24cb899a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f22f51c3beaacaa6ed434d6637ef184819ea35529b041b6b13519cf2b11b8889b8cae174;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd24f79dd0d2b4aab6bfd014bae47b62ed47e467d04c2c2cdd290fc63e79bb1bd1b3cb60a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c15c70b4aadce5a5c6da6a16cac7a582eb2d5a3db975609fcb89f2778a43e1495302317;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc29c166a563496c0038029c03d4a67c2d399563d5c8ceae0db03d0263bba38d64e6f2d5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d61d8f6d13d0445c7c8ee84d1f3417aa9c38c30a8310487f400bbe59324c57715096df0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1422823af438a8797455798e8e712e1f4b9d2fe7461c5e6ba9a0595a6a9372cde1d5cee22;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he059fde2e6d586bb71f9cc78365a3899e8c71d5df4383852e584be0f912f38ad1bb3af85;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126dd9fcc7a61dd9c85927a942652dfdead84d9c4d1591f55c6cd1744814837353eeca656;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aff9bdb1945f8028a70109c32ec1dcf0d54bc59bacdb877784b52c8f0864f96acbb7cad4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7aeeb7920b2748eb607939449467df7f2b47eec7f5f828fd937e514105b61be058ea51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf007988054a60a35bb593160305559a2ebb69fafaef0b5fc61127eb36223a91c4969c49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9b6cb8756b85aa5566738f188b831b39373f755b12354f09b35a6dda68783c0ddc66454;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183448166c92e4a457e63a65e6000f32f0ed69f60b22f346dc6461061e086453257e63ea3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9282418b8b0aac9990870a6b349a3e8f7fb237309736ef9de125c009dcd576202a271d11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a825d1963b1b9b62abb3ae567708518bfe84fed3a20dc20bfe505a5d14d64ba91b72623a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6e793ca91f3bd519238e564930c8f76f087ac4b303808c0488837365d16279c2bb29a60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132c5da354603291d506be1d209b071fda1b2cc0fdf4602d5077e570bcbbe85ef3ff7bf02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bcf04590d5e10938805d5de23eb435450e8ab44cf6abc1c77cc6b46f5fe03f88898a484;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2032a21fd0e5d18ca74d5ba670bbf2670f563824f8180cf1d7fdcbd60c8951e47cdfbe6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197120b582c41b4d8d401fe9c66305de6b45c09bfbd3bac724ba30f8870885c018e292e45;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7896d23a8fda7d3c3b0afa34b534f739edbc1a4da57281feec75c5f1e8ef18b28f20156;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec81b22bf7fe02bc634d2c908a625f6cc4fe05c13be29d929d5095684386a83812a72239;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he15029ce083919fcb1a552059cd6d21f825a4d5cdd4d0d34336e9995e665cfc6c5fc7acb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f91deadfbb5b0a218e7bbe9e515fdab4a34e1a2af8a72ba0f9f8d3805b44e5e1a5ab20a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14123b8f6a245ee0d6dc93e676b51a63c66f4da4cc6df3e120ab94fc9607a784f6e8d5f9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1d39d2c80818e6fb976616d9039eea584b307b79ee95e171109e5cb059d0a7aed187fb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfd02f49c57547302cc1e5d3e5ae72f808fc49d95032c037e2340738c0af024e879952a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haeb41971734e9c8a3b41adcea7b8d3fe5b92176ce952aff29ccac07bb41f88031e35c7e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a01cd31568e73cfb335857f80d3d2f514600ff4e2828ef12b620a8b222171d6fc0610899;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17bc29e485f7a6e049d34c976cf934d56a6e7dc4dc0319bfcc07800a90d1ff38fd348e791;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f602cb275f31799c98ede2b00643b007c85afc067eba7fa9c5e2adabbf4e1d42e869de56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19beaca228966395eb203d5b2400ada85437c5e69232071d51c876de51e81730e57834a1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1f4d4122a9c7b97714c1c29e03f425d38116c042e5616f3e19ba9a6dd1da3141f988a7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9f474cb566b5d33e77ed53eb6359662fb5a378514c8eae294be6226f8083be6b6ca26b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c01d11c05a8e034fc22541c795be6a1cf83d56f20b0257e45970e5f859a6610fe7a34cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cf3d9e393bc24a9652c6311812876ff99520823a2d66bd2018272c933dc284a275d95d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15abe388589a2169da162106b05347cea8602d0643edf3de79d1f6286b4a883398efaffd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee4eb3308dd38542af7ffdecc13be09d738e0cb6aeb80e496a9ea94bd3dc968306a8b5cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e80ec39dfb6a92572384a9999528b4e776389f229b2ebb8b5b2a9c13a5ec2ea1112245d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1075a84d83919850a7c0c6d82c5dd94fa4796f4312adfcd9dba2b04718cf4eb8341ff3902;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178d4931480542ddac3abbab5cb4505847821b0d5826cc553bc903422db63a1db0e5ee912;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1086df20f905e26efc4ac2aee4e2e67e92d4a98b26e5688ec42d162423914dc7f8b33a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb31bc0a894fb22e51d3ee14f11d788da79efc5e045933b955c3030b1ccc5285f14aa5e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff3becc2e835b5dfcadb355b960f1bd4beffa1a22123306bc5e85d08f0e97e963f4ea320;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hada1646b831b0cd0f8da903defc153765d68a9c31623d5fe455b504994aa8b97da0be742;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169997d74da389c52a868944d8b14a08f38ac625b238f7db723fa7f7e3d5788fa5bfcf721;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cf22da2cbf0890bbeb0af896d827f703e58d62908aad3c581513c91b2779a929e0a17fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ea63be4093578e7b3514e3a7df72d8c6299bbe888a804f8051c5d58a2ddb76c0b7caf77;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee2d213da904288d4b7ecb343b309f33a4c58e74df80da893ff08e0842b39f0d058acf4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19321d159b0b1ef399684cfc02106cf9becdfb330eab4c7810b2c73eda1e07d68673c7cf8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12772d180f5a70e318764d577ba62052a3ef77fc1caa97a383e973f61a64cb347a310d6ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha64c66d318e350553325c2c13818ae46c25fac372d4a0c1bc6ea230ea31f63c04d9eb0b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda922fa9fb281b22b7be2c276791399138b05ae9eb95ff44bb42212390af684e8814e66f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e8fbbb17d09ba381d3582eee600f14acd9e3da820555fd37da7e8df7137355b308fe2d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188fa881e1a59735bc94b50501182fe2cd6c3b1d2f67df11c3a935b0026fcd9d853ec590;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e2f66660cc6cb7fd16e8e34524fcb1e2967778c07e51bc66a0998685a663a07254a4f91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8009625236ffa44edcd5bd965674da88d73ad7aeb0e92c2768a5a36195492cbffc8fa331;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192e0dbc7d30f395b9562793f3132179d53f04a59558dfd4e16175da08ba7b507d91441f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae72722b386376ac2767a61301ef09d492b8c5b3a2213bb6bf447c0934da02d45adb7445;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6f88ddba886f0f2ed5c028c3a7eed734315e79e5e6793fde2dff1a1782653e249503478;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60ff10d86132d96f1d37d82ee53cd970a3b5363e7074a5372e3f91d63319d0797db5d2bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he981b13f9bd17cf1d415453f0953ee06793c34f111488b487c131393d4aad1714d787356;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4ce1a7f3c552a08760aa494173203ae9e46df03082b04c40ac001cb74a75d36d2211f11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f337ee5b8283bda2c7770936238b54407d45f91a6aa6a95825b83bc7273dea1ff3ce7b28;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf491835098e10b4eecc1eeb0fefcb881df243f9dbdaaf2ff03c051807ecebeb66bde179;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44610c0332f86df43fb4ccb9640cc0cee641c146214c77d08446144e875125cac1104395;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac2e1aa4cdf33f804812e65e56a1e9ee4d3f04bd82608c2377c5510e9e6f81f834866157;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2be846ffc6b884c3415256c46c07c03dbfdfa89172c3bcd39c6daa9277f4a9f04d88592;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71c9d107b16927286e745f8867405b9d59529c19f2c6d2f4552a4370456c3a19ac7db8bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f677ae5972999b18d8833285541e0de5a476134092d31be5c33477a56d528b0d841c1bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1368a299e7d22b0f18e1020439ee0c664afb45f754b9b6ea8e327c7d8350687ab1b79153f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d472d25ce49ec7e78a37d4119647d43298d7096fe46067870ec419188f5fc5e01000873;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9f5036dcb305df47eeb830b2b238abe63b1fa650991d32020c6a5798978da0cd117707d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8e1d864bffcc8131042bf4c471c1720f79297ac18aefba10db19a0e70c658ee8aecf571;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h426581f1ad571c7eb428a698c477408dd8c7040d355eb8a04c0f431ea7c40f1dafc8b02a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85cf172ef8cf6f0f5147fe90db4ff65d2edef3f6e36e4c336143187098665860d79164f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a17936fb8bd7261809559dbf8e455dd170bd4d31f07d857e5716dbb09b1139e5ce956e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4b9b19d86ac7faf438fd847e96d36f495c24427344cf328e9885f3b8d705e8078ae0dac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8c9f5481a8d8ee163d9625a3cf3d79d3e76b87109f6b852cbf542b576d2ea46a2f44e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1639136021e2497c193f78fb7e4a4dc5f6a3cc1d64fd5916eed61f68da8e397493cad0a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa28e1d6625bb24773a362ad416f099d5166e139a2b990b72fc2c2e44d7442a3426bf901;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c8481fb3acc3a83ec08f6e2ea5c02d789608a55638e050f13c55fc706355d8c1d7b8799;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f013dbfeeef2c4857b40790c83a4cd185fbcecc2fa2f67600816bab3d382da5a63d03216;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11f50f6b6af4e4e7f1c8f3c1269e4c803459c220eaae16a52a5facffe9d9d7e5d08d531a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ba30032f663d7e271f2a8f6fa32ee2f6051334a596f2d646ab2dedf770eafe5c47f2ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d92074054d896bd4bb743e05357667d2cb7e99859de026420753f5ce5cc86d9ed6686ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3279faf6a4c9b7ddb24783f40d134c4dfd07eeac67df072481a565c7ba17e6e449459110;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he78767703cb02ded3390c238558f7932bfd7d578e60ff4fa0f29604d8ea696cb04095191;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b18dfaef5409a2be8b659de6a67396e6a10bf94f0dc3f951c6f2387e64c77b77db1485b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162bef0ba9296bc056ce26e5ed17b00ca3ad598eb67622f9d8a51b802da42f6440c4d17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45a579029912cf438f154670cd176b5b94b5893f0c622c04af3771bb92ba0c4691885f0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3049d8ce23bdddfcd5e98c7e07485a266c2bee125de164056dbcea50a90450e770d78877;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc43de7cce806420d64e962a916fc4fde1dd38249180a2334c64f8f7c5fe2232d1862a5c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186d2e09584aa7bfab28d3be986f8c84d83bfbf367ac6e48ab50249a025d5de6c352fea8d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a85b25a4c98e30454a37d162f3cd1e14e19f72560567201ac1deb3240047a0b7020dcd01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b9f6303dcb0616d7c7da0946a1baee36f8746c744c8369e4e1bb4fde27423e516462a0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ea5242f81ff0b9d54c6a27791c64a1fd51c93c82ec011a658e51e183e1e0b95ed60e576;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd733b5c3badb65149d7d587b0be4db75d88a0f698b4300bb58ec4dfa4081ab67c0d62ab4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119ed05cad31cfb718272c9de81205c1653d2eef0f6904ef9cb1e9bb9f730d4236219c4cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h368b1f0e2f8e34c2b44fc86d832eaa67793e60170b370dde25f37de3c1e19766ccf96ff5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b4102def9231980a0527549799cae8b159c4334214ab08f19c488d72e2081147f68f5fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16bd081f138ad7abf0407f15c380567494db5307b63a1fb6114da515b5fbfa7cfe0d2baca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8a0dc34b5fbc3421fee1e84805111f66e99968d9eeb9e19f9a9c1b35f97865a2d12d7a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1a1f32c4047f1bb290fec29aebb18fbeb9fe18c2b45b33d1e18d3496ef7ca9d75ce7742;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd27d952bdb8db286e334b6152a9a4a71a9351d024039e8f09768bf83ef4c5ed37f502d7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e72a37c4b4a35f373a1f008cc49e0b5c826f254155f5ccd755a22c2666ac2abfe985d14d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfa43e4d636c8ba86ae11e9fbd2de24f012692ecdac3b0189529a1b7d073b2128b475a1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8c4d89f3100fc6fc588870b450adb4973114dbb12e33409d353164abb952ace9435fc4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc58c9a686dede331a66cc395fdd6445117af337a17d0f2d881055f762b26865626953bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h332145d398584ee20a6de1514550b634dcf63851ac693af8f1a762f9182c900c33ff531b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7af6ef73ec2613f179eb31eebf0e6198743bdc7195611f6b2ca7a2138a4e2ac6085d67ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b9deefe4c873ffe918de068f9ee887aba655a43be48166acfee4785b0ab0039e9c9306d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8ed79c3234efaf233a73f22f2921a31d330e26484a548367e115a1dcc41d3a319c4f7c71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h457fa6a365920570fef9c185eaa131e27e3f200ecb3675ce87c2d98356933c837728f3f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1910dc32bff28f163cd45e5d99c4c1854a6f4ca26297f40bc01df9562dfba0c5b0f4301ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f4fab26538daa2b6e42f416488a53bd77ac4f5dbebcf36455c4b9788f46c7f69a29d05d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2d3411301c5f4934fe1a9a53c1ad806d20e4399a06fd27fe176252acba9670878861a56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a01c3f1f93678d1741086071ce73fbe9c5dcd87646a2ca7c2605901b2fada56cf232eed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e114ed18be994b52a354ffc0ff1fb09b2ce7d7623f0ffddd17e5c4dea279c2e4fd7e7b90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h604a8a691adfca9e83d0585eb69e7ecc3756d3230dfed846eeae95d4ff4decba2b247a9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163f8a6e85049ef5a02c137f5cb06ab9abe15fdafa0151ec7de7d000494deba836ca990ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f405261d1d44cb408a34e0969b636d7eda1ff6b4ac5035bea8e2537a067093533743686;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4a35de94de38f7ee9a03a31b9bb365d9f4b365213fcfd198d1b2665dbcef29fd984ab76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195af8f878a92d344d56d5735a823a1a452b5417499697ead8a5fd13a0c5db39aa4025183;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e0852ff1bbef3bec3a9e8faf8d49e07052b4fec24719d52cdb7637aa61befa18237f1ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1957ae9a241398e3f33d8763f33eb0b2215eeace8dae622af90c1574fc87e952a1d404642;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c803d33428a4f2e656fcc82016141a85ba0672ba318ecfe6a0862ae71d4c99cda976583;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc041cf67d8299d80b452175f4fe2b1bd0e52d20cc6d91b81b0156ee0fd2c1c3bf3afe93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8fc3a65a60091e1adb45b60bc4f647c431164adc907e739758ebee19f822c8ad7cbc914;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93a880c30437a3c4b928aa8d8d6fb00d73fe69592daa96ba4a98892f8406cd9b9a078883;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e57563a2ead05db06edb5effbede98687c261b79a03dbb160bf7ad4120c0ff4f52527610;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16dd08c7ab878666d551db01873d3d121f873e7d83f8d7497e0b190fa03176dd4e8425373;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd956c6e7da090b36885f389d5c2940fe9c35208d9531fb7b19d0e891a8a46107a2271e7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28440e9fe17ad9021dcd09a70159db6c9da024cffab02f2b6778406ff61b6141abe6ffbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1736e0937ea292dd0e84376d8950f5b94fbb2b74ad0633d68b2bf648465faac7cad3e96c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12da97d80b55014fc01ec9a8d96188625c61893593a1b74891294ff517600f2409b5ce2aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51f9c0cf290c362cb07a8ee6695919de762ff2d65029399c564c86b64681edca3081d794;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfe800df014e7e7196667ee1da477fa3e1c2185ef961effe85a570fc146224d22cd35b3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf566a74f2b2d893e5d59129ac78b019528c1e98c12fc20a3cfe78947b9b7cec552e542a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf440ff83bbc5bb17c170712e2f32bcc06a522f6a938504b173584d89ae00c6eb609521c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1005ed72d09939cbbf2099a611258b6dc0d241b65545f7f009da70ea18e7de7944ca75b97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff767829e06710b823045ef504a77235a01dd368e729171867e3a5c655a2b95109d7621c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c52683058eb91e2d7aee88c71127300c7a42dea5ed4ab65e54bbb3cd661ff911965b5a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ec4ba5e213c66cb63da4ec4fcf227f1333b444a7eb6541256bc3f1af533745092ed2376;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he0c337a5a753f1981be18ac354e08f9a3a93c4cef693623a379c84fac41c6f2a7e0c5f64;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3498ad590826b257722221e467090c32d504185074513cb942662218a6c762e10f226d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117e9b175e8b3369b46b98c4f8f0c87d4af7e7aecf06ae0342095d80299eaae991f8b8e17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ddae7ac38c22bafb7c0f6fe3162a1bf374fc8b6851bc90177870fae1329d81231614422;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7e2f060dd0d13c4e13fd3fcd8e909bc233d9d4e4b85f4fe2d62de7b261a53280446f628;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1429468861ffccc62939fdcac9fa4edd276454864423af1b0502ea697f24d366cb15421c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159a8a1f772ec6d90c477509fe62caaad95b05d66a32e0ab505cbc7276257758e0c2dfa06;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad56cc954e4377951620b4f44fc2da1b9d895d3a35e289fb0a927cc1e7fdda731f1aec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef44446222c70e99d1ec16e3c86cbe6a20bc41d1c6a6d3fd929f5115e7cd38dc6d7e21e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca331765caa9dc10346a6abe158eb4ccaecadaf96446da05cf80d34fb02cd8b590245fc1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13afbefed73451cdfa7a2fc1a837f9784876198da01c56c56afaaee515101093295789e17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bf43830e76f464b04de80127bf59e998407d1d3b2aafb837521d13234dc2be32df1a4b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d80c70f6b11a1aad79452e8ef903c74138e073d6985ed10e666bea9546761c6f5c1bc8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109185f9959cfbaf96cd03847b5e5418b4d5439ebe749c2423b808af5a31983853a8f90f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fad42661803ffab8a76ce066a322451c8054a00e6b29f3afcd7f3ac6f2c5c300bdb350f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ec5209ee4fb97c0ae31225d2e3defffdbda5b29d7d6ac382eb1a018e4d06256fc6b5e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c83a8ccea4c02258d87404b09e96ce5622249723c4218d7f5bbe7b02137af7cd7b03a488;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h46da0773008818318dc38303cb53eade01e9772e35f77cbd8be8e3817a53465d221d8b2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5b39be9d4534703fb9bf357a2aa9fe66a43ae7cf86aa2d3fe6a7f8bb65012915ddb5cb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4568d21be8d57bf8b588f342e7ff39d829457d660ebeb181857be8794932984daddee0f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193aea849d62585f4a1560c30a1c488a1e14b081bdcad0457aae5a296ffb2e4becf05c2cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0fe619c289539feaa41d15f6e2c8cd87a8186ec1bdce5584a799bf4b75a6683c9d50740;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1889250242e95dab58d9d344c5dc338a0c607e7ce28eda8bec876b89abe91fd288bd11107;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7aff9a88b3d04fddb4eab82f3072e48e6313933b75714b0331444658c9a6900614436c18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb51da9310f52e7d7fde3eeb2c88fd94e98939156bb9bff149576a33dd301b7e4acfa233a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae0a3b293904dcbe55633d77a7d65690bca1b67673b682192ba3767e9890675e21414406;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffa6410150d2378a13f568028b48add13360d9d01bf199652dc10806d48a011de97c6c63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3fee333729f98c05652342b9f826c91fba71075fd60f0f3752006732e30155eb2a12b25a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c5eaefc96e76bb4c54cec44487d350519323e9ff270bc4304a32019e659091cc8290826;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189c6b6b1cbcc2d41b6941326fa858937ef197bec295793175737ac197c07bd887efe2d0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1680fd260701c07e79dea2bd8b6dd7466f4d5f0e94faf8c7ba324e343166d154e78c79173;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f2469dd76fd06b06c6856d9ae0f5fee5d9822eb9c3ee57393b9a7d0ebc4cfaf6f67e993;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a1a8280fde345fc3a51a603b01935924001334346542fca5631e57255c101b5f5ff62dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h649ab1fa87dfb09c31af4d6686b75cbfbdc2d4cd13b2a0e9c7b81187642d809389f87962;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1b5cbe2909bf4969fde9ea4054b91ff36ef3223ba3ff7690d54760be5bff433081767b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194b3767bd795065b3c000ee7be90c67c4cc02d5fa90543361e618bb7c0e763ea5b5eb1f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a5e8a62e8e986d7183f326a3ebe3f5fe527c548ec896559061e3bb03c8774ea6cd2694b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f1204f189e2fec4275b779ad85324eea8e2fc103de4308a6cc61bd521267da0a5d9bd43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17dbd3b9910929e091fb500c9c1c73b2c5ea1b5a7c6b068485424610739929e2c377b1b7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecd6c6b945b9bf14facd6112f1a6d6cf0d8b821dde16f1b2627fff0d43792dccecee2101;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9eca555b6b9bcdfc2fc2d8b15f949e8f4973813fa72d1f113ab67ee1786b1d6f4b97ef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d0766cdd988e6a0be76eb008262aa63d150930e44d329349961ede31a9d9ce7cbd95d72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5798d4144c250f23759d32904f65f3a068ceaa36cf6611d6613afd7974fc2cd43ae6f4fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1e939a8276c1bcf841b07a2bd3bb5126d74ffe5cd0752659ae770c617adb3f8548ff4d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fe52bd45cbeb5e21ca7b36057b01e37193c886e9bf3d9b2e822d6528548b586afe9774f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f2e2ecefb40024ef521912ad711dc440e6851be35a858f176275911adff5b12282774bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fbf1f050a689ac2644711fb647d92c231e276b6eab0f0d52cc1aa87548666c4a775d128;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1c49c1568406a99ca9ba190b8833c935416f3b6314148761704e999b9dd4fd0309bebb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a0073328e546719106db34788e28cbf33e3637b1cc521f44eb27ec2284f74b9ce001f1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169e7dad190e523bb0e94a601be3d781d22aaccd977fa02e2a796a9bfc15df699f2c50396;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11685168635500c2988115ba56681970821b92b898e1e0ec34efe7276431a7d5d3133cdda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1563659c60dba160079701bec7f71d69f38e72b1a1da974b8aa84aea494d2720c4823928d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd273f4fe88ae1f446b42467ccb4eacda37cb8a969e0938cb5ac431fb701c204797bc08a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd104a607425022379c6506e309ba484f8525cc714f7fa1bf1ae505add08481a223fac44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e9654cc142c3e2994fece30e4057281378c44793b0092f8bcd30e585079da9ae0821a63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha64aa0e2f31c5002303ca84771c889a1909b0b4caab6322809e03fee6409bc7765f181c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ab593a638d1048287120daecb7410b6df522f78fea6be8c6d564aaefd573fa2bb3a4e9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ada16bc9765af5283aaac8446aef1d332f54469c74cb18acc4edfc4366cf1da8594402bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3b8fc649125c68e1019cc5af3f4b1c0e88e6cd9b13761e5cbab3487cc214126d97e191e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b86fc48517becb5c20339ca127effe127306a50f350c5a783302ac5c54fe915839d6cf4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ea5206aeeaff12afbbc49725898998afd7d3e58d4415a874b73a36de8160359502d22feb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h995430e20d8ede47a9baa36b66abdc8d722269846fc3d07ddf1a57ceb2f44eed39f36413;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129ac0f283205489d0f9193aa97dbe1787fc06646b315161261f1879d8ecfed1ce3306e81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c50aba17b47fbd3121fb1affce31287abc567bfa08b4ded4d1f93814829cb27b2a7de817;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba6a330fe65b1d16ca29139c883408ce5e316be5d964909dfab4cd9677ed7757e13e03cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195ca8b75c2f6183026b814f96694c2883ae04d37d8100861729ee0d1bab4c7bbfbcff3f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afc2f12bead43673126b20dc9cb236648fd38428066d7af3935f82a087191899da721f6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f717ad1112689800b3cd82e8c69e738ecc573628f16c593b244042ead0fdade495e9f7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3a66b56709bf17bac2d9338699aa3cdb03278a50590a1d3aaa995835c90316c419629f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a82a3aa5064c2110ccd92eb1f5ae24564a56cbd0d1934ef67e880e57cfc40b1a71bce6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e855f45fdcb38e68ef1023890f2f01d0cfbc395faf48d07cc9bf3b5ecf4c49a5d64f22a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87240075c5f2001f86656da345c064cf432aa0bf652b3aab66b96095291e34674e8b4cbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d253fe506f0e1e6610a7ac632bbe041cc464e731a8abccedd49ba8013b7e4a862602a22;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88b8a3d5e2c6a6c6a42beb529b5e4b40eed6d11b3441c6c73d9b2896eb1b6a2bb8c8022b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1edb52dd5a2d1a56c3b63b611b5dc9fd03ebc34d9895a110248cd5cd9cd14d11006662e05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c4cd2d4dd52f68a6ff2b1cf3fda7f6b12586f67ff497489d7528d1065093de6d59c8e3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb206e7772fb5591f7d5ed36222ae7fd5372c78ed9f901bf170ff39d1fb983c6071b756;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h784a1043d2d9d61801e6219fa51ef164f73078736e6391d4c97428f57b300c85433c8e8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdec6f554f00f91617e5f4a7ba890ce89c0c443fd5a3f0da5f2b7cdf3b446ca1b124ccb6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb55eabe1c2288d76a83d6db10fa59f91f7186c84e46d416869e946db8f829df4bcf59c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1178b36ebc9f87942ea61a6b3d46cea68a074e7480ccc1f14fed238854dc4a9a7ddf8dda6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be116a0ad2355896691baff7aa8929b00e7c3c25d38bafcb699afe5927e3f34ebc850000;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa1ebfa576f2c2bda17b4568b5da2d91278078accc0ef2d98dac0c0ac6d68c75a41bfdee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6eab04ca5ea07490b20fac66091aff4c769dbd09167fa09b0033dc5b1f38aec8c3753db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b875e6a39018a7b92812afdeee1a01b84c301a223f4080047e8bed8d3bb2fb39e3cc3e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1359241a73c3a7ffaa818f74da35979579a12e952b6c5c95b8d115640813d930a12734e99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186c58296969f435015fc9d2d5ad6a48abdd5c251d1d12d4cdd7118858d419a5c0aab7a5a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h219868008e6936017df7e24d6f7576ec0ec65c1a31561dea93e6c9fc7a7bd7712f1045fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17729fcae2f3cf0df54f7fd89cdc64bc9e854e933a990c55694ef8a8218fb007e389ed40a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1080ba8febfbf8eeaa285321a954291a22e1f64e252293c9f36c48b8b970cda8f218ac361;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130fddea9524a1707f80059bdcaa9c23dd81e54195044958ed3f309806f7d68807cb3121;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1468706102641a4667af69806e3d533269ce5b750feb1b7cd55f229389fbb7ae92f4973f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17efaad77ae975fc7a6bd40453f1d7112e7d81bf650653f28dc58d4473379081e3db769d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da036f925dc77e04c35c755f16156352ff9116f6b49727218d430273c9b9cd2f7d52cdf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9379d6e126d287500fd9af04d6dd07fac9e28fdb64f5258a7e8d7496f49c5a6213b1945d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b9014f7eb9f23b873b1ec1041c641d491e3dc2d70b7b8e0959019336ef0819814fac3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a16977a66314ce34575b3e97f9b7f2cf861afa03c9b385e0e7b3ba0867f89a91e487c18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1c14390ee05cd74d05cdb66db31aa8668a0e001db405e8bde0c2cada0363101f67174db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f5ea883f2b81290b0f5b8c2665879da800ea82190530e8b7e2fd4bf0df0c241ce42aee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfdcd8d1e6793b07f278658d6ee441d21c7423de0be0534b25e6807f20b3ca79a0ace773;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be71a59afa1f0bf0d91edd704fac4131be3c7c8b3fd2dbcc844a650703c9861748bc4bf8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha20d2aeb0218e58a3404552d268db54cb4b2d21a6e01163302a7bcc86d0eebddb28ba2dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181f06936a656baa4d6fcfe3141201e951aed00e1ab8891eba2962d4d9287faefbc658eda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c12d23db98ed513b5fc6943d777ff5da589aa7aa1a50d263a85daa68ccf10cfb1baad37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd2271ac5cea6bf9dead2e6b7fca916fefbac71a7520a84119f04ea2214ff472d98632d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abdfea63e731b76f5c270868276cf120572e5355ff752cf43d5388cae7639353ae16261d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb2ba69132e0568bcdc73666286164e53e6c888619329177a653398f233199286ff983e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffb94b5ffd84bb4bbc2fedb4a195aa0f7c04e40064f749188461e9f37ea99e2f26be63da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abb3a45d15e3fabab87cc4b3dd17b459e7c4f37adab3effc1d6b7f7ec771bc59ed98abac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89f1950c197f135524cab351b310443073f5fb8dd16b57c7dc3169b778e3cf78d97b2137;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b83556f21225262d16657050166a1d0301313c49d14d98d8e38bc8400501c5b858fcd0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e890b650bdb309470b9649416a98818eb0c6dd99608a1a9ec2e857fb020d5655ca010496;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dce43dfba07dcbc280e2d728a9866060043077d8f22f8230f786e126f316b580f98eb876;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f403f8ccc66773c87b36281713eaa9f5e47ce60050379d7f038d68953d70d081fcb63942;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e1698b20bcd4eac9fa7a1dbf1bc5c7935c2104c794394d99b3884200a4defb8228c2bb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0694a8919252a12ed7def866022b744ff1b0cc7984aad5612d869a78971677eb13cf800;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76c32ecfa68c843800ed6972fe9c296a40494fb33997f4a2f1b47ebd1907f847b4f7310f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1406aeb3e8b78bd2e8f2a535c481396b1748888ff1011acc5b79e9c42243e40b0a0ca88b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h213971c440a54170ebbee253e9fa8e4ce23f178b6cc5088c1b3f465b923931bd974b9b67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124051fbd65f5088b37b9ef218ddb9ae913fb3a074f8daba6a9cd1e7ed47404406d4aad0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ba33387f00b32938b2ab5beed533226224d5295c31fafffa34830d782c3de2c363eb56c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63e0f471ffb53aef8af847d2a4e66e0e2f7b1d65b16d1945d0cfefec6aea11d1118b3be4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13505b4659f32ef51c78dc76e8481e9a95daac01de90817aa5871b573dd9f15c2aacab6b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10106e3c8db2de7c474a31100ea9c175eb8eafc81f389722825ea609bd2435ac721c9ae90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185e7b54cd3d9880c03cb15cf6e1bc88786e465207fea7f76e054bd5a72a28198429ad62d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0c2f7c08dd813663135fa8734585d7e62347cb1e48c6dea8e666c9f04f5db414838df72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a84c36db9ff011006aa1c6bfe880d6c2c5bcede04fa11c14ffe06fc9b27da3104b58144e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hddadc3489120ffc90b77c298d62f3e91229dc1a2aec1550bb5131241297768cc49be8925;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h148fd9ca38395ce062b8608cda0f7a58956f7b7d7e1d6e8a3f3fb2ea5f067cee037485368;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193d0c77bdc2e117e37368e2a3c42980100b96e086961329a1ad198e56f538a68c32b5af0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfc732985abaf02bc8fcb3ed7a355cffef8dd9fa5f158ca12c1ce7cb802162635d7cc4f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f7f55c77f2f504e4d1125dc2d96c1a3ac614f22d50a6cf295bdbc589b25950fb481b0c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a7f06861d4cc40e689970a9e12769b504c38e64eabebb26f785c58765ff884b1250987b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h729a66bb9420a17e9d204b06ed5a10642d7402f7bcba00b33d8b9a2fa8027f1df351fa4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a345c4695c5d7441d3d962e055ba194238678e5f103f929bf05f5b89d152aadce0b69d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1619856df4decfca767efc9e967fdfb0966a21755d5486389edce151e29bf4404e21d79fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdf584dd56ea7968e71bbd279e52989d09fda5c5b2bf3f60c10b3f75bc2475c1bc4e15b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fff66b125de09a4162c036fbfa2a291efdfa030279fade2f67801c532450583530fb9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116511a256b83287c5b584f95f3b75bb64ce7c77a7f270e22b34dfd3dab5d95b6454b9589;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he951dc602ecda5ebf26455e4b7b6a5fdbd2454fb98704e5dd2f55b8d66049fbade589383;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a957c83ba5ba0fbdecdb9857c7e0e54b7f35f6d7f8de6fc9fdb8d7e7aa414c2fc6242de5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3e5ed2b9ac73d086d765b60c582f4f923507809f37984e815394cb09113c2aa5cca14ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec3d891b2c776bd125ed821771d556c3fc34708473661bc131c60726d8d872115aa78501;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h325114aa9b3ba403cc9882d8e61bd53fd72fdc397b2f43c29b97b10a383fbc0d9fadee6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cfcd5d5021830a1b6a315d1d6dc5e385f5f2ff743950c6af0ece1cf43ac64e3c62886f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b938cdc2b08535dba13b907715c9ba0fb4687f6348e71be0c74503a9dfe4360274eeb30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1928d3b6b40cd61c8ed06ef34dba92666ead101ce657693faa59d599542c24c3896aaa43e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140197e56a5e9a9e028a2ed4d7fd9fa7260860fa8b58598843a5e6e33b8e9d604a093ffe1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h513897e6c033e4cd746aa9cb73d5535eb1934fb15459000f1e2de024bf10b9e310a24675;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e49233ee19fea27d5401a4281d24a0335ca916aec934f295a25b8f53041926b1e90bf64b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48fe18aca0605f63bfcdc6cfce6b6b176cbd7469294cb0510d28743468730943fdcf6a93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138a6f5b9a1255eb640a09297e63680f1e5e9992066ccc54fb1dce7038791e744a3b08bf7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164673dfc91f4daff9d7c50c7761e579ed6dc8b76d2d32c5d990048556dfac4602a924e45;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbdb5e910f076354ba07643e85deb95fb6c973c99b47729b2a62f7f60b16160d157259227;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1292a47eeb5f3f72827f830310d768433d5a4ccb800f724f4fb0f0cfd69268215958b0e78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7497f33ceef9a96e3f3e0d12f00bafe55636cc80163d65e038a87d18f4362895019f03e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44cc0948fdc0d696a7bdb2e4773b9436533926bf37c5db7c92d468f9af3a86079913e0e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f05cb5b2ccc7ed3523d8ce93d0da8566a678e1bfbb0ecb3e22a1ea82ab9cd7483ff55b43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65e1ede789439fab63298c055f0ce71cbe43d1da20558d7052b5810ad2f41c4cd334381f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1841de44e81f9a2f1aa72e5585d6619cbe3831ae570998a42dc21b0fbd1be7c6147ea8848;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h728b8d6084dc52218f7c145ef740c3bee66f09fbf1ced0d94e68bb5f7fc6b69d1d5cc110;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a852f782cbcd823969ed7d1b635b1954e0dc95f45416419308cbcfc0368ce5e3160277a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164ce06f13ab4bb11d1bf92fa2f06f516bb9a6f70e178aef3b97bde9dc771bb02fb597867;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h92fe277894873d560b9353a7f4dd6f7fa06d3ea3a9e4852a17f2aae675523ac275b61f5c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d87385f304769ca3f0145c1563e58f647f57480ca1f69d33055fb30ace96dccff6500349;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110078dd0434cce5ae712d34f3ea84bd971eb00b5b092be4eae38665d2cbdb05d415e0e1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f74f6c531a74778dc1d484f46c5e3b3d4d752053f26ceaad2ebb618f52d7f03810cc329c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee36e417bf183d0b3bcdae7e9ad5b51a44f8dfc54b5376e47cc263269ac795c3039c07d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132436e1ab3f53e423675b2eae805786cb644298f982a405642ce4467b108ccaef1c3c916;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h788e37ec58ab5d00efe38f54d6fbe96028a79d7750d215f00c4d85957bf4c73d1ca5d6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc582bf407026be28e0af66c5967db3f3b850704ecb0a2b991a331fdf38446d5e26ff5618;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8dfd7d3991f292b00a9573eb116938b55fec436bf92a306d83fde8808cf30bbfd99e76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c2c4bb31d3953a0177d1eb8fd5b7076668f2cb141faf82b4b0849e64f460c2a72a88d67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145dab2a2215c5057422b414595c08b5f77cb41b1fe9d290fac36aaba0e42a33695742f98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c884afe1ec478bd8cefa4800856b694ed4295d0e154f758bcccb7dedaee31a1b20becf38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1efd8b2a6c6ba6b22be7a076c651450c10f35d2d2103cf593cccdb8c51b0f55811950923f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10635e985cf62e09dbcf0fab7930176423ebe3f244a0b2ec332976d77b03b69671e1a6ffe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bd3d50d13fc9d90a9fa38ddc1716bdcd0251ce00c865e0fee47c235c54372740b3fd6d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1249eaaa6ef25839773b281d8f88d34ffbdb24f5d0e90afc26b46ea85d56f69fc0600f7d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25475ac044938705b090c217ec620546d878e6b02c827a63387fab8be18ff92f1f0128e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10229b5205db1ce35c115a8577d2938c0a667070e39edec44ccabd5ad40af59a76892132c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194adbda9d7e2c26a1438ab9ef932e62d4e181602a64d339b6a4087fa93ca5e47efd4c5f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187cf6473fa678df33a14a93133c144228a7fa2107b0c10e0c8a291ab7d01d3aa5ce9f078;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bcaecbb98654ad44d50f7c9304988b188665ac44fb9fa54b147be5d7435018a6b06a546;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf32cc4c3d604501276b2d752572d267a87adae84b5e50cf1b438d4b4989701bb58bf3a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad8449616f444b43fa8792c35a9a0b694519c7ada6ee050d1f3c881fdb654115838924c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4566ebf0604b8d53e658dd25b9b04fee74f3e7a4fc83865c544370bfb9d8368a3c12d75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a29cb8acb514a6affd87d4e8a176756544b8e52caf1194cf8e1da4bd30dc1d08446b036;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aac7e753625905cad16b78e072ad75c57e9e00e40b6d184fffd86050d939202efee95ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda23ee2afa786c205d2170f1457e2d0674b4df6eb79b5d85a0f6b6b9eef57940a8037e4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d58e2e70f3938363d593f7fe1365cfa1b1b430a7b881ac77c9e1840fe467ed9b46ab320;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160f188510413911595843383a9c2f7fd8d9d1ffedef85adfebacb6ecd312dec884471490;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172677377b04263f57f358e06336fd805786642aea3428b7af985c4afdbafb2d5c6c9d47f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbc06411aabcbcc02f6991443d841f5819f4c19e0f9437516d4828f3bc680035563adb92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha98b8e0bf4d57a794bd57e4c816b800e711560c5d67c1dda7ee408b5c7f652abfd5c4570;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9ec8e4ba48d6ff81d1ddc72ceb3d844479c29b0716a89533a1c779a2987badc7b00e16c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129b8bcdd182a9f47029347e1c2d31e0bcc74bfd4c71cc2571ca887e88af7f064438661b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20f4acb8da53e64505585aeed90f728461123bbc90ecb98ad07629630683d6b7064948b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3774dc3f37c3af298e4e9dca83f47734953c5090da733a80777e636378fe85a816ac3409;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ab45c67444cb3d49cca8599bedc5dd703fe2c313c3aa71a8954ecdde724f7f7d582e886;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b789c7b1fc0d0bc1d586d1da7f370417783a9825c58024ad2eac05fb78afd359424ae2ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd7c789c150bd5e3de74ae5a27d5cdf655501a1463ef09fa0ea609fde765038c837e0e12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd36059e80dfff094c6218b668aacab8e79dce6b62d8265f421c641fd053fc84e9ba28ce4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9291ab0a7cb6c8bd2893f339d4af657f875687fe1119c4120078a8ae4cbc211e300045;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7f04f6c2e3c972cbabbe30344e0f1962ea5ce499cf1a61a8b80ba31115b68fdd1d5cbb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7fa4e873a8b8e94dff645c127409118317133b3b766fad44410e816d78b35f22739e547;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c5fcf2588566d78496c1eff50e1486fbe3a518a547682b68a1b09a55cc8975ff7e99e75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda5f0e22557b9876e98fc3eed7fe5900d41ea7da215bd47e2177d91c872d6a192ecc3b4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121ff70eb236e747d935c3db5c57a7ce5794063bcb65d8abe4113d6c2a9b10d997bb92db6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12577e69ccff47cd3d4be22f89a973b3f20520a62a914ebd40545c2927f833b54a353a594;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd78db56d47ada9434e2b9775682b14a5c0a9a8755560a8cc4aaf9ebee7b35390ffbb39bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h688af19cb32263e8bfb802d04978edf3bce6d2b73cde731c5fe14595d7fd0633e28b185b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9714c1c9a609e14c153c3b32a4fedde25c67a7f2e874fa831a3f7e9f6941769bf367894;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50eef27dd85ee1a17fa71bc762d70dc9abafc22c5566df5fdd5f2396659929bdb56b95c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b1aef61b845cf085ea7d7724feb43d1306ef202b27e86ed4567fd7c7e53c5903c944daf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9efc1d218e845ca810419a080be4ae90c241e7338961cea69e9efe440ffb560245434c95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65f2e365ad98c8bcce807bb07a054d6332de13317fde5a66aa587d738d63aefcf6da63f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h436bdd87852b24b58705bfd4cb85ee93af53c295eea1073a62788984f6d5d2fceeeca255;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1906be4652686bd3c72dadcf7d8cf88fb0be63d5644edb6c1fad121d953739bae2c54a5bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9faeb19f17b7d4cd49d65654a94243e5009c427207303b7bfe2d1a4ec90f549111cfdde8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146421f3be4312c85f9a8b756752935ca5b3685f41933a51da25f78117982cfea2c4204d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb16a1cbb9c5116c04341c71f759e1930db5525638f1e107f24f090bd435f2c2607621c18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca0faf8dc84e1a744e3e4bb7b27a96dce8438c91f5efaadbe8f9c2a7f7c856051ecdc3df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51b5b7775446ce15b858cf25914f4b51c87a9f10410ab89507edc2020bfb164bcc78aba5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18eddf9712f39e3edacc522cc8a25aa9ea903eac38f603549a62504dcc76f7f43747230ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1997a73284db4c3d12aa8cdf513e2d3107d108fadef8a50a693aa1e97f722ca447e6ba55a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfb2793c7dc06dccda30c6b6c31a85bf556d99efe75725e1bd2aaa9c0eb4a6b62644c7e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb0e4a2a107f29bae35dc9fe1769293e27a46bdfd5dcead68aae789eee9d1129ab659d7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a2b2f2c76b0cb54563be56a8689b27aa29688740509caf772ff0d5a14ca81dd633901be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18395b2ded7ac30ad94f97145d995a841540c844ac24538e2c1e489038ffac7e6d12e770a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80fbda20bf82c845cc8c468bb182ac0242281298f28399b10780ce2c3fb5585715865885;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34edbc18bb00e8a5809ac1c1752600ff728c89379e2e8ede50f79d72bf0821b0e51cabf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37f1cca42c4b657a7b500285d9cfd612efbd58ed588d24ed1643de0ab5284f63cc3fee16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33fe2f2b4911d00634a76170f24a81b13a3b98fdc6b88e1e722dfe976b551a1e5e7a6c27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a5619dab2b74ea6cc5a8e6ebccd295b4ad606e383ebdec7ba8266fe9545bc2602b4e341;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c96ba711f52b2cfc056f91533a75e3d0870d4ed29d4fa9c4261c19b2cdfdefc70ab9963;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4603de26e5a43675dece45317ce670c4d282324544d4821cf251e8dcbc5465852022b90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ee77550e8a995bd30eb362d9f09261ff5391f87231518dd4055dcb3a514ea0d7cf7ce92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acb8987a8c704c549e71828f0b7481e4bfedb4188e446efade547083ab884c4861354296;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80ee19e710ac887ec5750c705099f51be5b144ec09bfcebae6e4288e122f3ccdc27c324b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1035aea147422b94c9faf477e459738d11d6436c358d27e2d7feb8c478599748446950230;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h213954e4119d1f8738c859ca580a6b373b35afc1976f466ef0385a095dd59eaa9652d53b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5d7a5d48e5e867b7640e61dd41b1ca14fa2e4ac21c6ad120992fcead5cd7c4c159500cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b4e7a8abf1499400ddc9131c24612eca7974e7112f6372da0550bcb34e7f2bc10c8c84d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1f9f7a847cc4d5c6d56567346dc86fbe6f3c744445c70925f6831c50f16b8eac5d2d446;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153537d05bd412780c7cf61b5a60243e8b4452252ae6dd20f458d4567b9a12cab03838d05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c7e1d1ec8fc565ab58eea8fd7d772674c9be2fd742f992ae15a5973c648a655e8bd6727;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1efb624556558f6fdaf54865786fc82342cdc18e5e3c430ea447786a9771f94f7805e7e8d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a2c24b773e957a939de2d22ae69a5ab4debf1bfab2bee1628a7b5e51190a6fbcb638ba4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41dd3c15f34be8c5c4e95ac8ed2e487d1b0f92078d409e191167504706b465c39e65e8be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1081b84d6b91ace857c7f94e0778655b5967e778d0da689de5af92f7d632a6e627ae16506;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c11ed06d55b5f111c7b19060e594a604c3b81b67e533e4b9a003911a26188e746798245;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d76138a87175cd14f054a5bc8f650ab9afdedd13249ec1bfd081ba0520fbc129879b0417;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc38378219c8adcd5926a282230b1dc70e106513da057db8eb4f56977894df426f8e9675f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8409d8d5b42f7221030d5cfa745209fa6edb6c7a52f543f2fc3462fa05bffcab6a32c13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3838bc2ad4fef709985b951d5fe752c7a7a9b3ca14f8bba1ba0a738fcaa76942385c1621;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d6b47741b04f4f4ed47e9893c3313a044d3f5e26fa6c932ea4171d559ec2ba19c9dec0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198507ce15ea50ea45ff77ea8b621fda4e718d0ca48f80168990295dfe44552e40ccc4e34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18525574578e4a3b0c619f312e25eb2acf1c762a46e9fe4f1d68bb292183d2c88eaf8d3c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1836eba1fe3d6365b7521994d91340e326673b27675b6e2a83c8be709ed21c339fad16644;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12701a69f436a8688462e156d0b1a65a11c67db30679593ab60f9f4e0cdfd35654c66fb13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35a3559a9c8da36a7397f3205f124e6f4951c5c007537a07781d8240cb9d7bd94d9ce26d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143cdfb0d5ead186011a3775b14cf27c6e1bb1b3f0100f69785da37a067d4d60ff2bd501d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c927350dbec1a9938813d4c13cdea79c50a6a1c21f28e612da98f09c0b0a71a50d45cfcf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbab3405369acbce3d1a6071adf128461b22070a7cbe2d32dd7ac4428e30ea207d3a7ade8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14454eeeb4a3b94020b21457b245a8b3dc0295e375e729992f756662ee08d7fcee14d4359;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2223e262ecc4edd90982e1ef22ee328b8d8517dd1a85118e9f6f1850117cd95a8d9b55cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc06edfe8fbde537d082416152db13e51e6c2f457e71417aa579acdb8aa0d6536c16d497;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3bc3e00448b5dade9164a93c3ff1e587b8ad51bd1c9f51cfaca9bc577556dafebe100c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29ea9b233df49c51770f276051fdefe105f1bd3d0be58a26d13fb8784b326edd195489f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123e89b61b0d2c503fb1dcfc3c6d7900615c518863410a5eb0aa2d49228604d035b65515d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a137a66f8205a33f5f9f60215e91967e551619ac55d5955403ca9c3b1339418d419f80a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42b9fafa0eb5a04cfbf73228a73fd3af7c029121051f393c92b90a93f928e574a171342b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166f4224dd0bf267162094b9d03e28e5d29e65d583da04831f7670ae297f6d93dc77efd86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9725d42b569c8164f0d6854adc07de3ecfaba259a7c1cd0662accbccdf93a321b419462;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c479148856c5da5aee68c6b859246696c07b146331beafa9ad468a095ad8da313552afa3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1350f197490f6ceb1e020ab5b18e52d7e875cfb5a585bb2fee04ba6ac7ae5c52456a9842e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17311cb8c3c3d1056d39ed201376003c8dd1c481f6ab90a66e0268ce2507137f93d3b3397;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfacd0c06695f6f149c69d0507af38a87bbd293e2396aef3caded4c1d9cb0ace8a1f5eeca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab816221f7d48d6b33c2a1605f59208a5b40a30b9b3e506fcb0c63637e6768a76d606291;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7aa2090d8190611ed162ca51aa6cc5eb5d7564838f13d3020e8740ade3f366ade59388;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1301b01f689664ef749bbef58d269390110482e1543e3a5788422312c3e3b5a7580ddec7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2802155240cd138de42e57e5b698eabec4b4a774823ab980350088cbf090aee6678beba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2d06b5565fb7305df5e3bee04d9d2290fadb9f54e60e422fa0856f331ce213e97d92ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a3d06e005e48d543165a26605c6e24904686cab69a38e4ff280c37792c5da74272c32e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1599ff19ae51587f06e35468c937105a01a64dc0f42a895b86f8dd44611b8bf8a8d5672cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef9af783fd6a6543138394d26901d5275ae5a3a1d817a19f566a44cfa63844552b84fdac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9239010bcd331eb391b34e7c04776fcf49508150a0315a24b33b2492b9680612ff037de5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ea6567e33b790ff87616715c8bbb826f9b5605a8af7c6cbc49a1b2d7c5e301f862318c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e064736c1e6cbe8bf3997ad119263e9b973cdaa344a9ca76f929c9c29be883db6216eb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8aa789abba3d5c9ab421004cf033076958fb55d0015d8eaebf8b55bfeccd8962313625c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1b4c469d8665ccd84c4c12664693d09257a2ed937a88e257e3c2b0a4525cc49d3ccea69;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ab697c0c333b89c8e57309761e654fb1ecd20aee4f03384659d4cfee5a0ededf66d829f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed9e3209dc46f96d42ce37802142c31a0452072fb1ab5f9221cbc22a4363025d292c3b17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28013fbeeb2b9a3907efcbaafebd5a7e247a19d246d240424916315e9952def14af34ced;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbacd21fa1a880be5f95db8dad9592f1c6f405df33f50d731ce843bb3f9b039a633d2088;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d1c3a1a551ebd0bc9bdfa3e2b676cd0f721dddb82664d03f4d5a50c595a12c00fcd64d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1037c097397f2ea78e8aadc5c21425eac73309af4d2cab37e5fbf2f746dbf67d4100ee258;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8ba7787d32da00efbe49780b79c75630b174eab484f36745b45233734be1421d8eea039;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba4446ef3dc22792cd1bfa81c6513f304a9beb21fe819f4969fdfb35381b0976cc35d6de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h863da252d599156730d61f4c9c69c185e194d2fc88054d6e27234150c62cd6ead4ee1e54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1773c84b2a3c1ceb31d3a4f03c93aa069bce10715f158d7e7060c39f02bf09e6ed24f83ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c29d0423df62db42fe5117900daf9b5280c33b2ef480375d7dae9a7b260160e42e5fc0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6c07822081147f985aee9a2c799f9c6cc1dee5906deeefdd562e7d4737111095edbb4c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a1af27a8bd6f2a126987353c319f7e3ed164fcec2dc879c031b23635eacc4db36b753ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e39d1bdbefda8b15a75964943299e8fd511cd337e71c6a645455d7a9c98183eac1c8176b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2753b21fde907010addc8e9ebac4e02e9ae402b654fd83f597e30821bfb8f61b982c890;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a62fad14f04470ebb92d3698e036522b760dd9d08746562199068ee92b87a3de7f88c924;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aa4673270cc724bcb3deac03eb1d1f6cf1fe7335e360e2091f303349beb8da971275867;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d6437bd0e77611e4e242cedb27c49c147f251b35a8ed3b0fcb7ad150f45bca4b2c74701;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54716e6399e7c59af1fcd94f2ff29e4c306d5f06cb408581224ac17f126b4fb666035130;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4932576a0def0f0b62f5ae1391dc11ac5d601936b77c7b3582a11b63b71e9663038c988;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b431de691408fe7559372b435590cc7a5a39e9bbd8260c5a1bfb5e5fa96aeebfd14bfb62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc29377100fc678395986ce7502ff62a44a82ba18d0eeb5471326d4bf2f2aeda2086523b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147feb44a72ceac512e20606ebdd3a8618e70b39f8383fd44bdce10d504a79cc0b7d68595;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c24ba88966065a9bd3611652f6d072ad51e94d562c2802da64e571304ef77143a66ba75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h941cdfd6e46dedf97b01aad6bc9dc638625c7bd2057e94c42db65801e98968f8e474cbef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127b0979a22d263478096d6b7f28a17c65cba4dc9d41b8072b3fdb18ac8bad15ddd66ba4d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151274d94a94b7884955ea74e0e6cda0425f612179955b07b5e8c60332a84562bfda25cfb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h335a1984cbfa196d95ddf799f3ada1ed0761fa27c5efd90c68a9a1c73ee3d90ef44d284;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e32196f02195f6aabccc974ca492044fd314f16658ef0de3f552dacf8070fff0de1746b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d274b1818727c3a124c3d09ea0b8f53f25a86fdf3a3f86b7a241492a048500ded6420fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbf5c228682377b5042732517e97a10495b6b9cefb43917a851bcfa94615725c9f3530ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec42f17ea374434b7454a1cbeb8ffd5675c1a48febc9e07ed23c1027aab1ccf260ff06ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4e959e2bf019d100ff6577f82017e315a493f1954ad2e573dd1fb7014756bf64b9826d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11808e48528066ea68a5d9c824f19ac0cedac550f1abee08072ce1c94aff25c0feeea00a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h793d6ca488cc0d06a93c656fc6bd8557a305304fc55baa41fc5cad887bbbb0cb1745a8cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ae76f632b9d77d2fd5fe8e8a4575d2d3b2689c0b0541ff76cefad83916145b8ec5fc178;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36152753063703aeb46403bafb0ac75d5594dc1b4286f4034271eeebe1c9ac8fc2dc6d18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf995539790842befe7aa5309f514ec8204ff92a4e0efabeb8dba50005db0058e97f324cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7b39e55a78cb31d5882c28d4d1ac11c50dd53483a617a61467586d6e5de1d5280990d14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60a769d4ea650c8b9d8fd06bef08ae4148442dcb08aef7feb1dd13cd8b4b81ca917b8a7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f09fc22c6fd34f187174399aad52664adc04c4ba582bdeef236bf0d4df8fc4a2a806df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10661323792516916fd38f49876f35c5f572216ba8d452a3d924b4f640ef5f8e16dbe023d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he779353ef28133db8fe6967d120a698ae3c65283d18904577c92a5cbefba7ea8ea2f9190;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7a46ed0b9c97192277ac17842eae67f884fca4e922bafc4f9ad51ad42c03e41bb5bc5bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c1c72c0b430ee7c469beccf0dfe165a1544d62081cbd0525f92f6a227c8200d09c34e0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ec70334ea051a7b9c9434158f19bd159432f8f4834f116c20945b5074ab9d90ce83a03b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1267a42607767a19a2d1cc13d643feb164e479ad40c4ed839d06c28145a6e827b1ce300e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c78bd0752494b0e32362a0a9d014877ad092257131d78ef2986248ac67c4bb21a680ae7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c088fc11c9127e0b4ee51f573d03697854e5f04021cf7191f8b4e0833ff39742aabbaf81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1432ecf61cd84c25790ceadc42f053b7631a9288bde8db4d7ffb1325217f151ce96f8c013;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea771ba3e3874b956bae0f0f1a148a12be88f72749d480baeeb7cd986cde6d7cb1e13e5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a31e4da97d002b1719c64ce8b2ee06762dc7cedfa84019948a5b47478ee42ad3c9fc21f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45dde632ad1ffad94835fce8eb3f2dfb77604076237b863f11617ec5aaa1b57f7d31b6b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdafcd428fc10707493873fd08f72cf00bdd6acb3ffd49461aa2cea640f578fbb3167b77;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c43e7aab7e59940ded1bc9442b8842b083ffab840d3add8b5d6a9ca3aaa2c24a89cc198;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb48baad1905eed2f081f8c95086c7c7407f700b5d85af7a98075b3272af561630cac997;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bbb2f12775ca382d40df21f2fd5d57926bbbb83853e5109f0ff817f0f8946f48ad19c35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0f5ee7828519bafb0590f3382dde028e4100d087a780b70ccbe86f7b365010d0517f0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfea7120d724887b9cd7dc2d5d12e32880350437e5ffe132a7690df63454da45789caf58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1304c8224e39d810116b393533a3b9988c377f09a8c16b2aec7a7679ed588002fc0defeaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be94a6e81f6813c0db93d15e3ed6c0ec17e4ebf9ffb637273f79f442ff1454772389ef1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d741c91f62cf550cb259482abf95137c508cae0648a0ba1005fe1b1e979cba22535f971;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b30f93fa4cd1f701d150108965ae05b257d2857d6b9b52759de07162c3acf9637d425d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c92069bbf1e7c60ceaef9d8647217f4b9d790892f8f843d4302a50ca7b6da6ecee65aade;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1db05c292f72733388deca1cb9da8d740a9cb4496f77e16e2260245313bc5c7bb13c7ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d25c05bfe5544076de6a23ebab138b8fcbadd70b472ba9627d4bd0d76c90d2c265353508;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16644b0c1a7f37b0b2575ee9da780aa2d9a73cc78669cba5918a21ae2a67d54afb04c47d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbdfd10b5c04ae94ca636c6370b6cb6b2654ea7cea61a85bd0b5b124dce6607aaef01d61;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5fd926526561d766845c9411fc495a11bc5eb63577605116e17d9e996a82df20f7474574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13650fede75a9d6046a0dcd9db96776ea6e2fcd5e66d86f09b834d3334ca34f80ba068fd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5426e261ebd075274d9483740497b33d451ef7ac5c7ca0f71d5e7860634cd48ec821851;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6098cf439b9c3e51f8ab1aad84691a3cf0b02e9d40843c9ddae470f6e6c42ca5a96f95d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heecdb038346b7a2c53b4267065b1d548bde288b777b5687fbd5b373fa0357ea161f13eba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0797a2f1008dd873391cba16e890311126463a0c372662bc2bd82f08322cb96796b0598;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c19db6c8775826d2210364b23c9dd5dd66af679ccb4ccd9e023641c051191df3594e49b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h46dc0b8e01e9162d3afe87b77ae86cfab7db22214b9099a4d3bd296602025aabf0958114;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e44a32572de4cdad854c68968022c49af7926352bb896066b633d863d2a646c81cda964f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c24c75b05adab5ce1039d7681bb0bd79c677bae8cffc37a08655bf11c644d5e20da12738;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a8cb7dcc8620b175c3ab6d63047f60c7940e5b00762056d46c0c4adf5d20fb0c9c5759c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1ba930547df9bfc04e96c022d31f858e5d4cb4227eebf8766e2317da4a4294e28488c6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1beb297f25aaf6e4c9d1d347348990e934032f06ff1559bf159b80aaf9b540d7a9b78b0f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a14c830a1e022ac1cbf56a5c2a482d45d0bb50efbe31836c9495d86fb333bee90673f48;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd5a17be0f126aaab63e25b5f727f2fa38436d96664fea5dea453d0d37cf36e953a2cbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd24c2d6ad472cf4282dd8166853d2e206423ffca6d87adb8a993d447156884f90417af62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbbcfd5cae54feb70e9fc0c6b8e144158e805adca64efebbb6a125c8787d3a1c14aa43ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5f9b1f0be383c0b0510582778a84896bf4e69ed2796da7c9418797a625eb3a9f2bbbec5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b917b15463a8c598eb8555b9ef994ef51225440abd6292b5164a15901547729c3bbf87c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85bdb7f64bbc3d20868b81a47689a02a1025ee590e352df539f89053432605c422065148;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1610337a40a38621b70270f4e9847d5e145979094632bce737a11522cca18919338110f7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d73fab70734cf24c7894d02aa7282adc78de5cd9a47a4d23a8bd6ccc8a1096be49b384c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb7ee33da11482117178522abf4fcf4610b487b0d12e3e151f94164527340fda775dcf8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7af165ec7fa9e65da6d55fe5acffbed7c421672555f5f99dc586edc1ea820f31609da583;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172b236b99cfc3b9eaa92866723fa4f182459863c90188092fd3dde502f7a9c745984eb6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b25eee7b828b63aac5c68cbd053b684739746706863c9d48ef11be5c0814d6f4d5e5863e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171f363099ed84acdb2dc07e4e45a7808730acfd3c21bc878c3126a6bdf2b79d1c780a8ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacb0f53e0cf2deeeea0b82764693d9895b0cb0c49560c984f1953c0a618ec72ebe1221d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1516484b7b298bae82ae10752f44074b8eff12c1e509a003e805d8d8fcbbe468cfb24a183;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f2d134b87c98f524184404e6da34f3ecf30e3e0511fb1fb77407b4d3061066ac3906cbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ebfaf831372aa3e7cd0b092103ddd2e9748630f13b20bf8152ee2c87d2da07c14350769;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d718e620fd8b2cb1506e492860d182a74b740f1bc7cd2b8bbb7a39209d7bd6edafe94e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1556b9682a69bdd4f253974197c0ddcc30d40c3a847baddf97ce87270acc66e3bd8a80968;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h932f386928516bb706ba8f21838d8e6418ebe0f31b961b19808c6d61c0a07619351d4995;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h417d00a2b94143bb5cff5de6bc27eadc6700277080880255327f7317c50370f706513d63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1723925a6efb4b7ebcc6e4b74c8ef4b526eaa42689ad35a43e5197a9fef3aea180b1b38b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bb8937160b4243b80690de787a77ca40b441b57d8ddb62af692a8175c08c372d47bc46d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1411407342affe5f4c4f9068d7b1806ccfa3991ad10cab2df936bb4bcbd3b41e09d8b0a0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174fd57e7a059320522b5d01ab37dd1d59587c7219e47b397d7287c16690cec48ca6bb3b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dab8a935f6f0c98ff722beefaeb4ce1ca21c077486a535c34088d722a1c02a048cbbb03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c47a66c7be21f46f352f1affbc453d827a62f4fa548cd9604fddb0804d9724bb5fffdd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afa6222e766d289b811b323d4dbe72a41c427cab6096c0506f1256c513bb7313538c146d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f125927997860c6755aa888142523b4b204231d3038ded0f3cd56456ef98510e32cdcd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179df6f6058604ca9bc832eebf9b43b3eacf66482303081a3e2c58a47ab75c7c8e58fd107;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6ec39dbef7fd04858ea1fa689a430ee64137ed44c9c43e7729aa1b6e48009cb65412744;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ec4b7ec9f4f94358090e4c4c78599ba7a63072c2780060abae85ea3f679942a1606e06a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1509d4009d05c92dba68faa0b7a57803c4eef9fd35335762256f84a12f3d2cd48eca28a31;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2706c4add30715a87ef21cf11e4b350539aa351e9ab89694d5cfec198a12520891c9ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde39abc774a4e41b47f4dfd9ac02b6f5f5316c8b014b99c52e466e82b68c627e2adbc1ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e9f5f8312ff6f22265a5aae6a70020b7a18beb82bd25c5a38a98f5524f0fc4a4760c09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129c5237f53b14b5753fb11d3fdfe134cd04a4488cab3653965c98709da9c59c56d5b7446;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a8f294841a4b38577dbfbba05524e11ae1f799f57349893b9822a2ad56023b4291ce893;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a554bda28b78778d386e5210f2acd5f57c95002f7f1a3f803fae824fcb6730e85624b5cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190d267f96a3031222483e3495bb107ff5235a4b7dfd36ab06519cafdce173bf3eb933c3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc11ffd13d06231e751c4aeba31be80074d7427ef3630f27cf657f4c266f06aa49905d9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100e43010098614fba76455e098896b61d9b8b9d3b07b656a5896d42acc9cf21f51635f78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec5fe1264632f2bdb96c7d10e3d0772ccc53bef17744da8903c514c79a884ee1f7ad68a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h319b813415c324649d94f2b9697574fb57f3a562bde3ff713dbd64680b473a1287c00937;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113dff9609f6ea018d89400bc6ca27b7c6f7db3dcbad0f3be7f96a6e4dcd1ee775d094dff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h721537d083481aade96eddce38197940ecd77371605730b779da75a40d3ff535c19164fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a940032f88e4719cc1bd9b621ebd8e6841c2367717f55e887048165297a0df07c76b138;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0a79c52507b7ba95d926d95896b5c8f709eabb7377af8c5ee789c6903a14cd770a973e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb7cc685837cd0a15564a5235ffa7e281ba200410aae09e4f5800443347471073f574381;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebb502bb3c8f7a6bc03af92250154d0f97361e694d88cf9164d01079abdbb7ae54da8b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11843696b2e189084da233d2e6c9bfe07a9ffcc61478e99b5a030fc0282f095f1e044683b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5150682313298ce2f18c60ed1701bd408fa39693e63c271dbab5b13ef63fdc40be69807;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h218e44bcb03776abbfb5ab9d7556e61b145972959c7da2da54ab4cd125c16e28d3a99499;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1503acb3fb204aff79c951cf55d95b02af5e3850b0bd11d4d4e2a3908fb1ab1a088cb1a22;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b05084d532f0751938dba2b6c99fb2c7c7e502cad0a162b5c132e34b457713564c5c9a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1081ee30897a6b27f2e197aa9c194eeae944458f72db443db9db9c0105bf7c0922fb128c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h983cf4a41ba80fcfef6331e53620d13447babe764d506fdf43cc145362f20a93f5e1bf5d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73866776a3dc98d2b6e08eb343f7b1528a3b889eb9d0757cb7ae8de1fd22e34bd531a4be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23dbe09c488fb91292f5053ddc81fb2c1c8b40356f283a7bb013cce8898ef49b8dad23e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6c42c9e0a85abff15929d8312a4ea123813870ddcbab9510949de712d95c242ef7ea39b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7ce6981efe73e07cdef92b0298f0e85516d0f101b27eedb7a298af82518ec4c8fcbf450;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc95af3a83de876545677cbe1cd8b91f895eef23fee0a295b0845c25dc59f8c254940bcd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h867a44a2ec62cbf940c6acd1c76c53c17f281a6ac77879b97ed302460f82520f2875be81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c85067063857a2740da265c0ae6f4126cdc3377260cfff45dac9fd014669fd3e83357fc2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5933801ace83afecc1989a49e39d950970e3a1425763555ba3d44db3c8d7191a8aff3ac4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd53630fb8ed7b08ff2cf99d817547380d1498c2138fcc53ebf133ff4cdf05144c1b5d4d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha71976520d565e340e548d3f64d39dd65346ba1356b1af3ffb6249e639196c925d44ebcf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13be8d1cf20922e26472673fe1629d69fcab3afaba1c109b89a3a8b20a2884b1bd205991e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc107ada3ca75ddea9c0bdb209db3d85fc117fa9a95e7cdb1c1798e35f629acfff4e64ef9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15daecab65c22ea7028c9d9eed27a033712a7f0ce1ddba1479e3c9ae4d7d1b21c98f194d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e0bfd34ee53dd4918c9aa9837f7cbcbf35cf2a736ef1f2fc237b0ee2e5e382d700f26e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bff80993b60cc5fc5828269a000996f8887f3d01db5a45c79ae7f628840f481edde34355;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habceef7f922aacb39d96cf479dccdda332a2649cf23bb20988f700b22c4075d0764007ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc89593d60cd89fe59d5aea158a292640bf3d6e68bffa3b4aee00e4c9908420d52b282a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fac89103dfdb6364277d9a3dd215e9a83cac5bb1986159e5ffdc87d669ff04e301e3b94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e808cd6cebbce2415040c59bf3715803bc7f8eadf8f36d70944a88c2ffe566ff8078b34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc8981fbe1ef94f0b1627b19b08307e59e3240605b682b5ab15bada844bfdba648aaa98b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7e2483e66233faa327707833881ba92d6db3852cdc3a49bf19d1cce2d5f7ed2d71a2ca4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1389866c8651c32bc04109fb81f63a006fb64a633201352dd5b538d3279741120c53f3b0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb856cc9ec12b35b543d5915719842c620dd1ca8d7bcab174475f9422fa15cf3192446b60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126133992e360d030977c7997b0c6484a86514e0f02ba68aaadcaa2b04b1cc1fd1a253e82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb218e3ff4001e3330d678992c725783ca0ee80a2875b08003b0e768c26341701a91b75d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc7e70bdbb7e937944e71d7cde93cdda508ee3abec2493077902d4eefe6160c5ae5d112c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24650a6af609297cd4d1102fed8b2b7576d0a023154165c9043af4e32ed0111a117ebcb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e00babb7e9a7dca7ba16bb299564734f400837053494f1d07e92ed6996f35ef86d31792;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fda3fd4117c6b1a6e83f21442b08556986e24432c7d92fc37128b2c79034b150466c3e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107b813873836e1c7a043f16f2ce9a62dbd009c1a07d9cf7a89f1c3a5cdb323f77d6cfda7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82a1852b66efe94607114e8812e16433064e1e9cd279802c735816de4f79d90b5fe2829b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h660b5f99c7a1f280e550bb60d256f12e6f136f0c1ff279105cccdcd1d8bd3edc28a57dd5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e590d225d86077e96dd5cb0dc17df3fed8ba5b39d0ae3a14ed77e6a36bf6974942fa72ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f27822dfe27b433ed9e8f2991ff729bd80c20942489a0f1aac33022986c2ca1964ea436;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a6f49cd9c0272affbb8142c8a30134c8a6192e18be5dd9e3363837533afef832eb1f01b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1364cc77e1edb61b15ba5a322a79f4461afadaf0343d7244ec25cc32adcf429aa69a29775;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5e5a98ed931d17afaa8dd986d9de9819bd816a9080d45418a6258cc4f62fd9ae4c7af0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5fcba9b0a7f33d02966772052599b11972c2714b27a1024d6b3a5224a37a8bb8eac6789;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17779cc12de425df5b49e44c84eaaac59081a3f6cae2dc6d87dbb03148722b392d50a2bc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a96f627243e5bdf776d5230171417092675551908b688d01b7070be44cc41b26f9e43f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha16ccc83eacaa33d875d8692f27f573cfc728929cfa4152e55256169f15fc5408a1ae9bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1934fb6cf965213afe649f67b4637f1cc65528539cb50e12bf7f8d06ed3984f052071022e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f65ad7e929645d316406b054c9472e8be08c9e1f2ea1d094b66b96d20e6b485dd066a84;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d54b9d643d8401ed6b7d76505d6cca751fc594af2fce263f42ceb8e5182cc379894cbdfa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b99d6c114c993b8bddca0db3644e9b33b3ef285edc056c7d3026deaf113c52f13774e44f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2e8a423e642e8da8d8e082550667eedcd7bbfe202f924ab83e7884d320ee301ffa34b80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17cda6d359059f5b83b40d7374fc82f0c5b1d47e8de0b14ac797d874458a9c5d39a5f4c2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187648e809ada75aa988ba7a678e3436187807bbe8086a9576433de15167fbadc5ce8bdd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94180410b2906ef0dbb8a00f47aecae9d3e9c9bca9b67b1ac01c061a63a704fab2362aab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cc6168242b49d495b1f4f23a12ce8a804d1961957c68f6a2847855aa302e1758ac0770c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b2691ff61667b04a5050e657ba1b2819df6d620976e33d64a5e723e3e2eb5e160cdd10f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc819712f43732a0eec98aa58409749582cbd67d5c0d5c56da115eb80312b679e27dbbc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8e8568bb851dd50417457860db0cc03860f5f4e7a3a627279d57263422f9f9f9e510f2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78e9098586b08dd4ffddc5ccf8096ccd6994ad0e0c6c4dff383e6d8b95372db30ab3121f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12731f9c1eff20d0076cf8f134648aceedfb5f73be5e647b50cbc4d80aa79550b23865449;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h608226a47069f6e4ab37545a90a13d2bcecdf82c40c774405f9a46e156b0ded9063511f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103a3f9d89dd43de57dd8dbb16f86d14a089364e093779bc52c689338fe9e2b982f1f58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19525ac8c9db58baa0ffb5aaa0793ea20036bbe468cfd02bd3bcb8f839d1e798cd899977a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5af993ed10b1bd6dbd7edf6caf191f3f6f23670c3e675d106f2e5ac47f5bafa681e3d2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc8fda943d448cc4e48aeb18d105e91fa274ab97d348bedc04635adb47338301bd5d1c3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91f234e49719c7900a1233a1490a6e249ea4d6b2783604daa2f9c1c59b3aa1a5871bc312;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfd9a90febaa3de03db578e77ceab9cb2300e7376c0a67c532cedae8adca1a90caffbeeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1946d36f0acb276c303b39f3a9e8d1f7a651f6f6fa70671a5b2461b3a9e2adf3ab02cb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a7d0e35377781db1be92bd2849530ff81ef1c0ca0a99944db38b3ffdc5d0dea0e161e5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdca30ee387335cc2bf20c720754683f3d7a161e01a51632d763f440515eee1b48e9a0380;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183bc38ed8ad2061cbb0dff8a73de592f6a7b80162168c9146b994f3dd408372cd758a7e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20398dd3a1436c8c7cce27310d221cdab654a452aa1f4535a8fe0039c3a3b10f22ee09f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee6eaf17d8b465a740ab4a637db51ba331b7f40bf42ef063d1f70d2239564f6fb978b90c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df39d4394a9057fcf5753326bdc270a4a522b6a49ea97530e1d488593240413016404dbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc1dd46f235a9cf571e5f52e8cd5c995e30bb65fdb49794619913dfd6288f7e45f8707eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11941e09d72e060d4ee0b08e98b342ae95c3f328dda254e5812b6ee866e86231ff3e509ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9139ee95c5e51689df7f563e40cb3c65b1ec179a6f15d48fadecd8686fad72555cf33b08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e270ac92442d766a5eee0b1849625bf9b4ba9ff4a132be013da536c04399c831c72240a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cae9045a3bd6595fb99fc1aded5373587987cf4d5c311b616f836622a1914d3a17f67a58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b7ed8b413cd10be9b7b1e1ed5e3c3d74b2a7cb92fbbeeb340fe44d626563c73e13280ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176fd0e2d554dff15204109a6ae0821eb603ad48a9a1d9fded568dd6f84d17cf7a2c8c65d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1249ef1fedd5b7744a652a530968e1064888a6dc88b559eb9e8f835ea6a3301c89354518a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h465447b936865271cbb8677678b59f1c360f30664decab3223717c15e64ebb491c10198c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e420ae5793633bcb7794135df13e09ca01916f228368b30427954dc3274c8e26dbde3b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c81c4000d8655f9086e107104caf43b0f69da6130ed63196049983922cf752ff23d3dcd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42f910f3b1ac038fe35c6b8054b19a8c109c17617c7fa4887aafa978e8c1708ec89f2453;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfb5b62251151cbd78c75fce4131440d5f39d536955a2416de35f3b617c0183773d3f520;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f45b3356dbfcef108094de32ac2ee26f4be48483ca25be970ff64665ca633e5e6b25dee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1653b82804ac123558d050e7701881fd62a3beed50c29a62751bcda139b0d345fedce5569;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18eaeed1d292108ca1c1f987ece242debb0ad08f0d0b4817797a37bcc01598224369a68af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3137aed7491f492f4c4c432874e39438febdaa01cd0135d38ea72ef6f3c17bc030cd335;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e92b4705050a03972944a93e72ce8234a688a5ac71baccc7050dc879a0d078053b5ff63c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c871adba22e152e06f9e3ce111a4ab03e8af3a81ad20af50988e1767d93f6757ea27765d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1f72ff77afc8b9347343876b05efc4118828dc5c7fbf53fe30cdcaf848c2e222b53a452;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dcecd6a0aba495ce38a0e0bb57e6f27086e344cf18d0fb2283f4b91e879fd80bd045cb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162985c731089e056c00c51790c8e4cd8fab3018910e18478b5cf3858808febda39b4c432;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b17d3e3390fb03d93007c32a9584f8938374e60cbb4c256e959d1e8401010103635dd2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c39adaa6f0d41e1f269692a031d6d3c4c3f2d9fb219609f963f55a003ba0c8d61c5a206;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f41ea67382dec4d255a78707076d25e52f2cea1c7b6047a60fc447aa42dafe413d8eefe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb281a039824e726da1aaba7f2402a674dac4cf35d77e12816918ff04ac9592bedb966356;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c92b279b6450009e60d93f612abcd58e26321d698dcdce08b7baff421d0dec30ef2b6d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0e2ca051a17e7164606cbb0175cd89da02fe27d6f95c6fe04d7b71f097ce23a85c4c0bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181bf10850e5acc9bfee4ac627bce49786c789c1502893407febb8fb92f829f04d8df4da8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa7f70008c3cc8f40c41ac3a941e159c826c2a8e984928bda87b21c4d281091753698bce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2aec516ed82c823bb2768046b9af7cc1af895b67e5ad448712042697f0e01caad2091abf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e68304e3266b6e2724254a560e5e91e0d31e9831f68d40c8e0ded890f6cbf065e962707;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h450b26f458906a0ae5edab714a9053cd07eaba7b310b654d1884368bb9225fbe599025e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34647125f859b81d3cda00bf162057466f9c791de9be0b0318f63d88f7cc1c1b0faf297b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1a87457530651c08548659c3029ec4dd075f6f4053886f61f038f74aa250d0c9a20223d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63fda60498adbfc2d04bacc59b1c68e8054ce58282bdd5036060e7015073e81034b5af2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a247e4f1c8947558b3d9c4f924dc6978f073261eaf794a5ee8756e5b8a411844efe31af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d61f166e5baa5d741b228d909c1a57c30c98be2b8121036af472eba4113139356fcf2551;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c9a0b1de12c951c7748f0ed04673f10255dc798efcc80e76688657971be65022ebd7d6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c67ea70b8a190bae744973b76d17650f0940da8fe263ce5f84cbef11d6a337512db7a6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1552cca8cf47019f6c641cb21073654537e12f7fcebe9afa470e20e58782539368748186a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h357849788052adfb87628aa579a051ef75a9a78a22deb428e4c5dfc507363ba3566f50fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110a99c67e6a1f96c2b82c2535f5e7e2512cf0e4aebf18cf4a81a9c6d45104738adc26757;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8090d2efc4db59e6b0bf3b7c7f3fa6dd5171b8fd4d3f57a3a34521b92b84eee346fcef6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd14d799e38cf5b743c819197968f62ee856416eb1330ac88f5f44debc71353f1546ee38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eac33050fc593a659f2b63a7c4970161861b3e81f7d54342a3a2fae0e82cb2044881405f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd70b6d8732ad092f2b1c2ffcb138c0d5ed63323342bdd00431c306694f3ed4c37bf36e9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cacbc31f3f77da74fef77e44415eee69942fce9d69d93d23a8faa762e2095f7e1ac96f0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hddb6dedd99d7aee80919a41a227b9a937bc351696188ec9ef073be07f403c8cb8b92aaaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5070f6544f24512315a5727caaed688e0ecfc6e3bd9e7611f1db0c7731cb9ca07cc33d7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e90079c2293dbdb86a6b5bea308a4ffeecd8179a9396011a80db4b226651d073d5cb9cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d02e6039d706378213e1532bbacba58e8517017dd3fbf75d902ce35cb012e1e3912deac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ba4a4e03e206d448e298e9d533c07b85edc03201334796e592ab4d28ecaab38f602dd05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197c430e13cc5d52f1eff71ecdec02e764a25670ba6ea9ff55709a6d0451187b8c14adf23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af15be9b7b2b834742be66b45a721a52b693cca25ee7f7a9ad77348e4fc96cf06782a4fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3de7cde887c696d397600f09d3cfe4069900bb974ef337e5e4ec359152a0bb41bc538f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3318f541e699b3b262f3ad2ec99438ce8db2262817083e7ef29e695b4ef028636f33072;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9db0d4c00a73d3969e8a54403be0225b995d7c0747a71b06091d620ae18d737a5032d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19351dcac035acbff9aad3bae89e55c46f30300478dead410e7e80f2b7b32642db5b480e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf3893c1b73f8cfc6755a33269b5c0fb0c47b1626b7b18e60fe1f33af016b1cf9194fbd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10317d487516fa73fcf72208d7f9c605f875d47ac487e71930c20325021fef4acb0131fae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h426b15016e7be027fa27d45f9289e5902c1025a21e8959f1a67ce491441f0ac0075f4122;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1163c016233e93829dea555fcc77a3fa7db2f54a6f9248eec72f28fde0a2e1c056a1a3b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebd6ab961765c8b17c251cdec03dd9aba2706bd1aec0122cd10c53ddcbc4e4d15963e8b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb244c924c42d329397cb53b33d01f13596dbad64536c55e536aa470988be4b3e17b36f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe28a3aa7ab7d2558f4581403e8ab79da7cdf69839463ede2d54d6f3b1cd6a4b58b5af13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ed0ba6fc6d1a6897583bb40a4e2d326abcf494054c467d890d86854f40720c831a8e640;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc9ef325236e880db31f39206899c79bc9da145e311cca368d7c32913fd413b7c04cd7906;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h516b2f4aee186292a8fc9e6023d1a986f8936273627dec844c32ea771928d42af92c51f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ea3a9bf27c99eee5c4dacab77dbaea86d16fde7f49f34fd2a812e70f8dbd29bce1e716d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5320f30fd8691f0ba8f1d50fc13a3dd4d8db15a68a66fbbed92f01b5235d1e5025f8190e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9f6b7bcd677c81db1d8a55388b12dbb953dabe5f00efddfc448fac272aded8b48c627b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cff7b80f248c0f0eb1b7a0e17d0fc1a9f72ab50cd8c569af8464d126b3f5a487dd235e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155921bc02ecea0fae4a72edb0d90a8a83573d6592581e6b2babaf9e02731e34c482dc3de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h681a51161baa613d3e734373561c26f67895af6e7313ae7d5b1cae959b25d2f5b6d8971e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7acad9c0b7815545640aca6e472956afaa950358789a9e6e864231f2261fb7ac2f0e3674;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4911724e86465a1dc0944732b31e4b2a0fcdbce4bf20942cf901e4aa0585e37fca2dfea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3678282dcd91d44d2180d64346342d7addee91bc56ec3f0a142e5a23c74eaa8b5287561;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c5bf52f7a598c5fcce368e965e0d239286e400145595dc44bc9db5e6caa4973eb2ee58a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16166ef67e8e0cff73a1b29aacef29e57f3b78c87e371acedf7b82c797ab2962cf0d5ab94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d67af38c936490fb254e860a0b53175d6e126582a2815ff72263295f3584d58ba2bea17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1433ec9ce6d186f5badedae8bbb616d2b42757fe56e6020072374260493224728a22b2889;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138570afe0149a1345c19030ff98c6b23d245658ff1322b6028fce5f98ba01a1ccc725b72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e321c922cde4a92233dfede9da8f63413cf3100be6555353ea421165af43d5aabffbe72a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9eaf315f6fde5945fc3aa5a8f75d62500e50d66c83417f0490f5a78e52e26c1e18f17ce5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e37b834c73354c0c119021d1e63290614ea0e7a6da232341b32ae3c77545c791964b8a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe832c54db872b527b7e229417b620b54862faa990c6f2e4b1833b06d45eb5dc46302e0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h40230cc13ff50cdd7287000c51251008200b887c76c08296d53eec174f6a243386e132;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1989330259beb14457908aeebadfafd6798a062c883e7b2a725d2956a467ddf90d7b5527b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18781c91238c50bb406d4dda7677e613a380e6b44cbe1de89ac24e50c5f137b1af8737f6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a226fd04932a02f585da914d1e99270d544c35867809a6a18a1edd53eb9cf96ef06b053;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h746e81de6fe7385d494e537bf853505fffdba9ded7983dcc45cb51802eaaa1826b90c80e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a5ed50f8a4b80f886547bfe13140c9dfced5d8b51a58d77bb627d807d2c0936af8b1f7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151b0991251d155c59dba0d99c142322a09e048e56dcb65af4678a8ab30a897840a15ee37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43cda9b66ffc3a9bf2c0f038b4de12e8e939f9e4509e3150777a8fa9020554549d6b19d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81c2104ca3c1a70e3c2f17744a7bea53cb17232ea932caa55a717562cd0e5d64a0dc5e52;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5073467fb688dba53b2277df881a01eaa53281407e9463df168b41839a7e3ebf04d1a9c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef68dc54413b787a035bf624f5b5214dc52a5c430085e5a82bd39c9846bd1ddcedf6e027;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9f974cffe1425a28c3c2377de0778e03fea3a3e4d6bad73317edcdd18f93d0f4d2a84a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5111b252dcbf828eff9faf4dc3ec609e15a8740a4d8dd3c4cbe362fb3b5494034d4cd09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118fbb0be03394f0875bae20ae44752ae1f7a6c597d7b7a2d0e8a087c534f9d4fe7e28574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf643f9c140f2313280151371df259cef4c937e727c599833f204e721bb86702c57ba216e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25aa90224e8003d945000c69137eec506e696f2fd56cb295d1b23279c869ff0913300304;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14964c1e1f033ffac7821c03e63dc2ca055cbae28a2008aa2ff487e789a9ca76358c278f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee29a3ed543d16eb4fe9f0d6e7a12eef3e78988bbfd99a6f85458d7731e7965cf564c70a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bbb4df5285fb016b4afc169c98ddd87cb19ee74983eab9b598263fd276993bd6b3403ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1f1b94098dc8b2f7142c2c3336bb3197608501f35e29015dcc6ad679a43beeb4ff3d125;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166633011db2cc2603c69632774da39b3b81109b2dd5e0f33c6088d605ec042b5d9f3669;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac78b452613e705e6968e6cf0fad48628b600ae83f33bf981b5897a073362792be11f37b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113d60b979f1560e25d7b6f12b2ebc0b2daf1a41b4da1c4339e34e0bca42355eb6904b29b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84bac5a480ffdf8683d71a798d0d445e0320e529d4afdfefd8fc0e589ede4a5211b2339f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c63d795d1165c92dcfa242d7c8ba1edf35df560f65cdaec34259ab17a1e8df9dc172dea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c754e625b8e81483610708c9a72b6fb15dd611367dd588c73a62e9c2db5bc0beed4b0530;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7df32bf693d8afe92da027975e3f0e09b9a037a4c78f04cd80238731249aab571bdf9c62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69b227f8a7863f40477738cd44422cf66030117bcc32a6dc9c46a84252eccb0fa10ff631;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1600be4000c26eafc6a6699d2bf074664b71d3923ef111db6d6ff828e41d3d24c2ecc9bc2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ede6d6fec70903e1551a8956c81a05e1e637beb3da59498c6ca98716638d0dcb0600eec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95a5bf96c3893927b994455c2331589f1459ecef09684d141144731a9317e223dfd724bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d2c06f186d107f1e76673e1214c9076ec9d03f6b73be249949fb0a44a58f20ac426e64d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c135dd06a87d4c1fa6aacb264009a381ba59716800d5414c7dfd5172a5e09891dfd7bc56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12eb4b9f8b1403dbf4c10541a5bf0c6686595467c95738ee20a254b8b32c85598cad628ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6b7d96a9cd406049ed34bf8728357ed06d2232a2f0bc559da850b712f45900428c775af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f198d59531c4f0b4e507e4b2728c49857c4d3cabb0bea51995b09e11c471fb0f0f90df7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7a1cbb9cfbda44b3d1d034b47fda2b28bd2be82295b68fc088fddfc0588a8e42c9bd9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d93306dad55184945727169865701a8eab48416297577ba5b6b9fb191a4bcac0f11dc1d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139716b05d29a954f99765ab9157eb7ea201c024f26035595190190c309ee65bebd085bba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d5288df6b9280e2530da39255af6e269f46e36b18b3abaee5875eb3be058c80b5efbfb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9be32c414f4feb26dedc7db7628c2fe94c80d107189f815a27d4d667eb23319f1fa1dc83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199fb52f2fe8d29583d5facaca3968dba4ecdd6c16f07cff53b1cb1351a21617b6b792d8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8fbee4b8ce3e5abf530952b25a900b2427252cbebe602ac79ddd5176a6799e2ae8f7626;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe3819356c368982a2eafaa908fa4947d01681e3349c7077d582894d390017dc83563826;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc36684d5d7b5ff9256e19655410a501c61c6999210bf97e0b3c1c6010d9cfff0e3eac1c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha656f75b83cfb8c1615a1227e66e686ce3cb37b1aaf3c39021d81d3ac066af57d653f11c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c085cfaa8e64d343f11475054a48d1531ca4340401e4f4d5696f7421df9cf33f1f85b95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119acfb1144214e30636fe27eb8d30a6ea7900fac41cfe4a000177cbcb18cd1f82937a072;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eeefe17028ed450485ebbcf2960576255706cc2a504b0e6fea2367119f62f5a0018eb84c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abb5c69cb76526fff4486d0bbcb38147232b8bd9a8b00f94ca46a043013abad440c6c7e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f8aad65137fce4e9a6af66b763afe2d2f8aaad6844bdfffe891cdbdab98be527d9801bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1bdfe009e6ea8a481f5a9e75388787e1e16a601e60bb190175b60f8d591e944c124e812;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11614bf3ff949038f82bf43c8c8f7497b34c0afaa432df2b1ca24ab83b12120925caa27b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd70999cdf1884fde5b455fe4e8949c7523db144369bc28dacb9bb96d32831366eca8d930;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h345406acdbd48fb671fda2ca2ebd81f646f75ea0bd22c165fccf5cbe5aaca4dd229a1471;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1041c3e00c8aa40769d25e44d112746a587873dbf1d809f49db8481c83959cca1f37829de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d43305f8af3fbad5aed8ba37de1ea85a639682b8739f71af7a69e407e50032e661a6519;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d61039de8b2bc98815d7697beb7716fa57c526befbadbd759a429c20ffde39c81d05fb7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f940d6de711991822a45182810e0a519dfcd40b1dd1d8de65b6e8e5117918f4e3c209234;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de1d98044eedcf2bc6d104630c3877700bf9a0ee7d21ba53acb832b83d88e36dcc7cc61b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d714fd4b07a4b33a3211a97c26f70de26ab3f166428e7a3f13a548cdc9dc239202e2f9dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdde5fcb3967068c7cd4dd828ecd4e57e4d152d56e4b7837015499d1834487702652657af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb20fd5a75671c821570e26f0a913bc9790c6d71b66624f31db24006c6c8f90c3dffe3a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf8f100052c75e066cca12381e25627038367dd5d556606c1ab5143ffa97835c4cc0f1b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1008e3f18e76dfc122d04c45c8a96b54a6a4ffd9aec0709ae0e716a4da21c9a512e196b8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c701dfca7ffc2d9ecde3b134f25a96f238a27134667ed123bc150d7b8e2a4c45850140a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8401f0dc089b09a58b4434ea933e83f86b4e4945b29489d3b44824c54ece9d0fddcb62f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h925b9f3172ed1bbb15c2599d4f220a569a154c1ee0ebbb33461def96a0d5930068956c37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149d81089d6d1ef5f30da01817d9239020820f9b4b842112b1bb191d8b22bb65a4c0547fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4afb97b30c2d8c5c74e5f0acc4c2c6947127b64000155d39b557ee15aedc1beb0905580a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d75bd32c2429a4f4a772ba6103fcde8f5567cee49f68063e5d4a52e0ac1fa36c86760b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he168f5f5a3aa9509923a31ada740ba31dce38fda03c41a12786672efd22e358bece37cc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ad80c1f3120694c89f3641c3552db1541aa7f38f61c4c64af64fef6059558021c8f7bd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d047366acb66a84d42859496165cabcbc940b45d6efa37a25b0dc37fd21af4f38523f30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131ce1c253a357cbf12f48d785b55755aa3520f59e331ed9b890b822a1f0ddd13b21c47ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ba2c49532dc23a150851c04da46c22baeb4598f483b0e261b7bd6ae4092b9ba862985ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78672eab6e51f3522f1a4b689538e71e86f0526a6384291286071fa3f0b7626d2fc0b83c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3a338b3137eba6d2df58796db5a8b13d8c603369efb2864ff9233d84ca7461695176380;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bc8d36b937decc25d00488ea14bf4b23db114215f6c828a2538f40981e90a8e4ad277f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118813cc122d123dc9c377001e0f3a784af31a90606711e75f0752c95eb71b5b5d10983b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he79164ad8070e478385416b7eead95d9a713e7429750b6b8be68e5edb541a1c32b6e3701;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfed6fecc9412e53eb20215dc13f1fba5acb940f7f6d380942c79de1d5357615ff635812f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cc0f0f14b74646e29dea2d5704e3e91259c8353d18cb63bb71da92687990b55e228bbfa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bda549c5fcdfc598af1537b8b6261ee5380537e6ec4bb5ab2afe6f63cbb4b5ba181ad9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1446055b0010c6bd2dab99df24a6425c56e55d63f94f97190dbb0657b80d5e6045d250482;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h515c595923cd5fb4d2bd08a34749ddf137b911a12d795b966d523ffbb10c99a758c45a9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1531176091b8e4edfc06540050e33439b71cc5ca246d5e8d318f59536489a56fc8478e56a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f81cc78b0b15eea0fd679251dff64aaef0433b964eca76481d95823eee2d01637c9181d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdeb4a018b53f27e517ce4d70a0ad0b2faf13ca2bee23fb8f3e59636806b5537c3e6b63e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h270958bdec03f465cc54c6be62f6b70b86f8b68f2d971f54588dceab34378041b530d644;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123178581d4e61eea2cdd85e728420f75f3d27d50863254dbc8984fad8933037ceb9033ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24d3da6c0f3455f1d3323c9c2376bed8ec00b07d8e707a580c53ceb534cdf0d33ec023cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d51e58df914e2e71e777df281200581f422ae990334492be91ebd067c1aaec1a93b4a45;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfc14527b45cf5819602942ddc4248c13b1ddf0d3d2f6345d39e142a36dee6d850c16a90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e640c9a06e7c571ad6ae80297c7addbdac9a232b5296c382819b88da1f0e6d1db718222f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c0a4f96e6ec93159ed4d8296af4aae6a505f2c52c2c726ffb6e4227b670405f73769af5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56e2f4a5d9de334697f389b7b8ecca6c590da71756d5279ee77f8ac3b5f56a464fc50448;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1985d6614cf42aaed9c4b3e985605aaf00f4da9721016e330d45035f8fa1aff0897de6e1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6125fd56ab74f6da6ff545976d7bee92873379cd1c5b2c7c2b55dd6b9df6c5e844a537e;
        #1
        $finish();
    end
endmodule
