module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8c2e3452aa89669;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ff9ce2094abfd38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ef0ce03063e0c15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90a570adab253740;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h248ce68e028613f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ce8ddd63c0bbb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9b2f4ad71ab45b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f5f4ce11e1c320d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8daf4ce93354620f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32d74b5f238f43ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1e21fd89d87a5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc1e5e9a353c7220;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had6a20dbfaed13f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c0542b0e092958a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf187615f695e5a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h669eaf3e43a1dcb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d5db2b8cb8edc53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b685d01d1916085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae6dbaa2f224e13a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2365824cfd7bf85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40629333d98887a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h309504905d3fdab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7ee7eb43d80d36c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bd2e19f77a777b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab815d56c7fb6279;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h470c382cce9b35f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf07f23a068a77111;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfafa3e04c67d1117;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec344fbe82eadac4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23da32a7f7d2e15f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bbc428230417c73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4f12b4a54a6f584;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6eb84cfc70b246cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab2653e7155cb0b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80a474c361ad8ccd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37df4144548c7f47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e9fe3000c2ba96f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53134532b7b5ff4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h891b386e0d65ebd9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0b8fb5dc4c490ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h258f72aecde11e26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81586c715869aef6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h570f2c9aa4b6bd98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f4d027b963947ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e1a5697021357c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba3c549a34807376;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha98793e9c2217e73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20b9817bbd4a903b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf74f770e5fee0938;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb307b0bf4dbb104f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d85c4d14837ec0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4de0eb5b9d8cda13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee4715e80c06a34e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92bbf69dca103d39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e1cee254f031a7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49f4a698e471546f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2aa2477aa0191afc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8d3d237a99b0af2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf29adf0d5ca00024;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8e30b3d120a1990;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h174a001bb2ad08e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72090ea09d04b97f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dec92b8870bb7e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e3647fe002a0bdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h757bdb4b8bec849c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d846702da3d8eac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7438d1571424d78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59f40a0289146a4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc135281592985646;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb795f85dc2fe7a87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ec76445606ce69d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28cf1dff6612c154;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha04394dadcf8c4d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9795f52a099d4997;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f94aa66d3a3e6f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab247bd08c35aaf7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1074b8cd7335dc4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ed51d99a9947ac7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h547b60e00b2598bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h685f2a2004048c50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bf9e6baa0432a20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ea3dd59795a6af0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h361b47a8cee89f0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72d1a5b4a972b6dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38fb4fcbb675794d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd570dff98bebe59f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h632bd37d721c7fe0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6841c9fc080ece0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b16c3d37a77e8b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha44f1c324622e3b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fdb09a259913f41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52d8036e49385f2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h483634f2ea799ac3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a4e592da10de3d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaf85b9830f2aafd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96d2931a024c2dee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h360a01842af155a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c8edb98d8281b3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36350b47b286dd81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha86a6bf0a0a7209c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb477bee349e8e538;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h850d053654b09261;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc13227ec725cb5cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h467da381c64d30ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f7d3dd1001825d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40eef1e374371561;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8787fce34bd55ce3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c056a42d1268570;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb432e11d90910121;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha595c3c02bd9c23b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e3862df4fe38730;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h430d5a8c0eb272d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb12c4c6d7a5e9154;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77d7b13e64cb9dd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7da1fb46b8aec6e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf27020791fd12ae5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6779323991f7373a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a2332c7d297ede5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h662bc8565116b64b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8730f4f52a47dea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb085ac4e1ead6bcf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8db6bf0535609d4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h438d447f83cc9b3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a61e9346458d426;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb077986f81ea615;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf710573fcfa19b39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cfd9c29de45cabf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6d89540df38c45b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5613a2e15631d15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6a0e0519b9d7d25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1a2362d87f037f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac66d3e1a9cc10eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65d9a7d1a573d564;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbaf1e19940799879;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fb24fd30b77564d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38278e30695c1df6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf6aea3ad4e0a7ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha90a2acad9807282;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h957bb6df608b9192;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e276acbadc5f90e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7c7420ce04bbaa9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc85588dd0ac9c772;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8fbba01be3a7b177;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86de7cc3540ab7c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc1046a7478cf77c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc97498f29f13dc0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d02dead4f1c72ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3662da7cfc89e2cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd71b14f6e515c324;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e48f22af7f77e5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc52f0bb15377fdb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h208758f32946fa4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dcf74213c043672;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a4d88757b5749b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h427a091e127c6c83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15a5eb8790f19867;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90ee5edd246fc39c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a187735b81d939b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd925f016fc5e30c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67af415946cd151c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha588b302d2a93c8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57b64b81937238a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30e121ba7ff92f2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h240052d329a13691;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd45f3f752618d248;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e096b8249dc88c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha88df5218b4b618f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h807cb81f9f14f8e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41721403a595e9cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56704c645be02271;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3be211c0061f9b05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebd3f4c9599c2b00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee0994c55248c28c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2ca73c542e1e383;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5914438c67850564;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a29e17a9a59dfcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb58677dda7dcfaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha37b9a08f0d32433;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96f7225a30eefa66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1865331f4e16ec1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42c38d47070c7650;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf00720f8537c7a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbab89f5cf0c144d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bb8c063746a96c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34cfc94563d7a0ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0680fd40ef0ec60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a3f7b19de60ba8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1415aa410b30bbc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43af15afebf0f83d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cfe786bceabf528;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ddfdc951d9572da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2907e8dc2036972;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e35b6e11c216c78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49f4a6442bb781ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h155494ed99022c66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72cb7a2f578b035;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5df55dc5aee6c97e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25b00b8033410003;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d404d7d1903d159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9e7acb925e83749;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2e8bebdc511af73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc45ddf0c52966752;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3a517fd56c50150;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15dd4cb6aa86e2e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5388f9b2849eb378;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15c41066268bb60a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22cabd73f7c6e3cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d790a5e4edc1e7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfab4bb6e53723308;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60b6deb3a93135f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f1a8bed50dfa039;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadd66b2893d1cab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90ec5faf5b610f1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd402222b9ed07bbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h575ff830a7e4edb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5420d2dd0ba357af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb58e550e6663ccb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21d4275b3f26cd14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52771b87ba06346e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd6bbc0c8e3a72f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h385179938060711;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38ef8fcbbfdb282;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9de6b32e34d5c87b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1139701c722368b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b93d9587a77a915;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fbf1ed752e038e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1faa13b971b448be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c1249f0f7b42f9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51d1955aa0b0d81f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dd52038f89fe11b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb49d9dd99babe47d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0b6046c9bfb0c79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc5404936906894a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha27f586170fefe13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29c6022a6bb557b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5aa4546f54ffbcb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8864634ee166ea63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec6fc5db9c0fe7f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28ca9681d3894211;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39edbcde6f2f3ff0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h839c8c5134445541;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2872983813825745;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25a188891f290e84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f558d2fd7de8aa8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9d23e52a35cef72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h230b1e429a14198a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105a93b7fe78e1c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f484d48763d0b87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc42830c1cf305e20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7f7055a321aeff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha22920744b8aba01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78ff839604d4514;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f97147edf589f39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h246f4f2f52e2a29c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62d953c7af159ce0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcd22a9201376bf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he01b535670a9933b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4134f7c4309c9865;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc57e7d00116f29cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc56a3bde153777e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e3742c7e69669b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2805b86b7a3b1904;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5d6046456c9cf20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47fdd6079d687640;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e79ddbc2671ed9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58930a2fb05c91b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he579decd736a366c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha12f0b3866f79368;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4059dcbe85b51186;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd1f2091990ddb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f040c43e9fb07ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77d81416a23caab2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa1fea25121f2d90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he623a7620dbd9889;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h792d41503fc2d838;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0565b4a15dc8974;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb175bc35b1b0d6aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f4b5ecb7a868ce4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc33038cff21abc1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d26ed79f87b8cde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9febdfab19e11ffc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d505c4b34e769a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfda990561c33e2e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h889aa126ebc46f7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe721660c45b0b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f54a61b9a10d8ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd85a9b65249b0c45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he94aa67335054636;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h241cc80f9efc625;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7d3b6731be83ad2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69a1b80fc254f4f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd475890e59a485e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h762035f20348a30e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc39259fc33a4b84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fc20b5d88cf5d9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41b506fc28bff4f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0fcffee94137f1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4f80f4bb9356e6f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6fda21cd47249ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4b79f464432730;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d28487e6545b9c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4b792713d11eb34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda18b322859b8577;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2d1afffd262012d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63dcf330ecf84c50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23270981286381a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he79c262b2830ce1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb256663d3a777046;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa1f63ab2920ef4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb7f2b1e2d3c2590;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbbcfc5534957821;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f017fec180221f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddfeb988d0925e7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87784d11113f007d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h878ab1e99d3730f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7896bdbbf4f818c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca2afe8a65d17b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a5cf937343af820;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a9647e181e5c4d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he03a0624a05330ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a043d81de74fcc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86b28bed425f547a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb502c516d34ff5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1016dc245ac119f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28f1bd320ae5b243;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5396dadd6a905cee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9b54825933ab46e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4aade53f70f47cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea03d6b2aa4873f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0e19b9c56b1db8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd350b49a338da5b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75c94f7e629dcf15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e4d9f46e770a68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d24a8a43a54cef1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8eb28f70872ed7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b360214e48c1b52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1de0c0d27767eaf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66563a0ba30dc352;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a3815daeaa5e74b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a2ffb24e74c0abc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9453bb95aa58e97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68ae28f38e16149b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13b6ef6cb1ad9ded;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46639d7584d2684f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d972525174c34c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h104cdb3971700a46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51fa63f68ce1b52e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ec34052c296ea99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h554d964648c6388f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9523919f54974be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb3efb2849b01914;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h649e785b424ed567;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf52fc5869cbbd4f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c3c65446a319f65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a041fba5bfa8dc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc97e6d0b0125ed19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80c92217431d3502;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5133259a20bf07bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c83092b830989fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h221035f1fa89bd3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h620b14f245fbe8ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7517ba8e1b051ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6c8cc12e8f5d890;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc0886cddc1c1998;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a429ced33016a28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h673caade74b7e12f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2071ed2df21219a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dab654561ab8bd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccecc006ff8a5b34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b542b7674d62124;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2563cab686967fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa73cbc84870f7a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24cbbe93fff255db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b41f2769c9c47aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4050d8b2170af612;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h805825d12a54c27f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9b4fe215392e159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d0fbdfa0c41ea7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f19243f6e601354;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ab438a8f1ce772c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36120177097ae499;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d9b00d1adb3c590;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9983afe37a545cd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb799ae7b8ff94bb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb17b9a8fd9823d7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe5c80c20942eb77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42f1b3c1f6fdc656;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68ebf9551955a1c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc86a384052a12082;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h920075ce62f8a356;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35f7f7d322b67e53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ab9d6f8d2539b9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd34c84b1e30d460d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d2c320812df220c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91ec5814c6c05d3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a17f4c6d8c7f0d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc0bfd5fc281d163;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd797ee9bab43424;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaff47414c9f2dd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b62ce4f7bea0594;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2a25235b0db9cd1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71b22e083852ce6f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad0d9649729039e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65cdfe63d96d7c67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c3d1c8f9ad4a23e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf32aa70c66cec94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7378b6d73fb06e45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e485b92d6e8f65c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c5c7ed1d7225ec4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb486420d7a72c372;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha071bfbcd6717ca0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc56543f31e68f065;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5a02b9708c7522e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9bd1a785a86e1a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0fb545f4d5fdf80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18cc93df9cffc4dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h358f0fc542eef9bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb11bd5065fd9be70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78b9a3854d3ec62d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec787b7da50d1b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda90150a27baddaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98daa78aeaa099d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56bf7d17a18c74c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1c34c8d9cfd7069;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cdc4f54d0162012;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h789af71ac8893214;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5e4d804aa391e0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he749ab3ed875203f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff960b59e8317138;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ee22b4344d35bac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd889cfe7a2e5638;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8620d4e43dea2c22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h949503f305513d4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b5e25f466227d1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7df6da1ebbf9fedf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb614fde0a834d15c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h343f9c81aab70504;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcdd3b5a039608aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0709e9ff6f54988;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed5505ba1f69c04b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9536074a6702492;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5922f319a92f58d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5efc471ce57f44d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h957cedddc20bd0fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7e0b09e9a5c24f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0c0c8bb716b6224;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f27ff8bc869838d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he52db6c9846a5adf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9dc329fc7a56cc4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cc77f328eb69380;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha93c28dca4d4537e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8a7368ac44a6eb9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba950a64a0055566;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61fa984190072427;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0a0ad2f28c9902d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h402f40c114be1886;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h634c8a3e42dbe8ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedf73fabefe67a84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a15f1ec719fae2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fbb27bc8a6c1a7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20ae24fc55a04051;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h178d60f113b08817;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb672b14e94a445e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha339925235648aa2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4cd955548d7da4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cdbe9366438db97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc19be5a03a346539;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9cf2f72150d12be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84f6b7f144b478ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2cca3b1f1a37653;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e6da35f591174ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfed00d24abc06729;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18e1d6efe7f5284b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6d05721312ee265;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7978e1beb4a0c13e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1db8977b0f56273d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c320f1911911e19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2983582736de4e27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h725b83bdb7676683;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39d7e02b73f38360;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3ed447c7137d0d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had820d0ce51e7f6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda5a7fa3d2e0ad72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3946e5d5c2bca006;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bbb18b14b1eac5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf643d29981c677bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16e8f1585a9e1b83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb8e22959f7c1545;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had5d3fd7c017b63a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha07215202ba9dd9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaf9b68e6a4e5cb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0011132bec49e88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb69a6b308cb7b3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50238962da99a941;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7eb1f88450141d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha896470dc9e2367;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77d611b7db3b36a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2770dfa96be24377;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc146864511e646fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb78e46cb905dcaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6c3f0ea97e3ca3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6cb3c4ce74b43dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf54d3075fc35d7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96638d8a84ebd3f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he37e57ea097ca753;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4aefdfd41171f135;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a2a44e7e507bddd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9b6e463b966e95f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a314abe198ae767;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4271f63ff381b6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73d23069e8ceefa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f64152d2e49750e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86ecd59efa2c3992;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h741dbc87f55de1e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4cc024c83b80f42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbb71f2a0262a09d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h471209d5770f96e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19889d25029ffe24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a5f734ce3a40fc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47bcd8bb4227ae67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff4fde1fdab09ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b1e322c7d8328c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb67bafd65ae554ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3be255c776117d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8826bf76f6da482f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbbe28b18da4afb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcccb5ffb4fc938b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha230bebda6254f6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heea286d084e8073b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7388d892974f8b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4df4214ba77e9ac4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h663d3836facd3230;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha68cb4d4f71e0fe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h156ff0b110a508dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha642d43a6d4c74b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd449522614e2efd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa719400efb4c1de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48e426b1f3d83379;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6aa2a566edf379e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb383e5532b618eaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb380767840f21ad9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64eb90d079d099cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5acc851d3ed5367f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd42c76a67d4fb139;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h955f008c84fb3bb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe090b3b8a55f78e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c1b7fae19f0c0f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b0ee88cbdcddff6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2af5bad7dd13a028;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habfda0b53df5e051;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67d0f255efeaceeb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8bd865492761495;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8442543220698ab4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd27040e9ea7ba02f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd92b4e77788b07a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2456b8bf2e2ae1fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec0c1facd38db629;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h642a864c27b0c7ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0e9b41955672f0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8968025122a8b335;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10b6f4a31344584;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9109023111e21d1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1902e032334c155;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3242bcd68ee214f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89abd804e5791f72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d6a04b75b838de0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5bfb426f22549911;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7de654e0995cd279;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c40a89b0c111ca0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d2760aa5f1e705c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e0b1d978ce8ac85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9107445f0a0aafe8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff17df87631d0b2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h765c62aa19441c92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9efe50901e4f79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4837821ac08647bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8ee65c26dafea07;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5855a97d21094430;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3d643317d228bce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5bd61c93e6da10a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8c78412503f2db6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6bfa6fe347a5990;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ee32d84d649223d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e43af173693dd5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42f5c17476569e29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6782e7672fd020cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f5415aaec180818;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9225dbc6c6a1b989;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a789d778bfa0a6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf90bd9a30d5311e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2565da04203f9eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fecda129f154740;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ef0681ab67f1d5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aceee425ca3b430;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h877207abaa9b0abc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7af5a6667e983cca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h556e19629e121edd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c2364dfe149e344;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9c3a9c138c03feb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb20107836e3a9378;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a2cfb9cc512315d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafbb087f76d83695;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h510133048b0ae73f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h240a58e90bf443e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7320a479e6e9001d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e3119000311186d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3543872a439192d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9a3bc59abdd0f37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he13fdfdeb5acb8f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c4bf569bf79612d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c357b2b78cff13a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b589cafde636c38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd13da170b0e576c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89104383b2a5b4f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a65e18f884a3ab6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5602a9f26d9af9b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h884bca130ae5037e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc46b3c6cf2565cc2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9cfd4b4996d6bbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15b31527d7ce995e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3b6e7d7aa8be3a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8dce4d437eadd48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51ce4ea86781e93f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7408bfc7ba4acdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc26159b5d9615fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4f7b28878c82128;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d89cf62b6e475ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cdc82e8053c67db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79465caf01c58371;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10bd0f3f5310adca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc384ee4df8116029;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab578dc59fb033fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcee7fd596c0bb7d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83823941ea213fb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61baf647173369a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e143380d822b7ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9e67208b0297be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0be5f9585c0e318;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5bda2a900fbfff8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2fa80a2ae2db822;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae14ae573e69ff2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49732d930087561;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27d592b0e5b1964;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73fe0c9d5f6fc244;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8171ba9a9b23a41a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf64f1f7f1bbd4776;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h632bf9417c137235;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab125b7816f21485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c95e2ec5cedad7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cd80ddb8e22a407;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h390914a5a8721eaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1484c64b6dcbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c2d20e4dc35e9e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8352f30b123167cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdfe11bb85fce60c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1400b98022688e8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf9a9acc50949123;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80443ee865bda824;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea055630a047cf60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94bbd1ae1e313b28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h524ad524d0e1b0fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e33a43554d08d29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6b3d4321eacfb7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h528f6c5527a314d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78a4e5fccbce9cec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he208c31c77e94ad1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heca26471c37710bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc10cd6f7c01835e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77e113ff72bd9992;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3098fa03e7b3e309;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d0a0e40aeef0f9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d825640fe4fab53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13388c900ff5c0e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h120a040cbc4a1f4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f1f3a55a7cbf544;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39afff66b60bc12d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8d04201ec8f13c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce1ad31549af22c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94454179b2c9097;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17796d5ce7f4d94a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cb48c5d2cd0dd00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbff52e1dca4138e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd900d661a378c50d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he54254679e0bd634;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5233762e6a1bd22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0813f52ad7152b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34e342f0aaab21b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23d5358eefcf7637;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a4ac86e87abe012;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c73828744a1a9dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa511b40a1d5bc2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf2234d474629966;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cb33efeba9d66f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h970f5fb436482a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45e30d64288440d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20d412a09913bbaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1a9073abc5f3fbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc387b1186166adf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99ec6ded45919b0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24faa8aa56053207;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9556efe5ae8a51b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h380ff28bf9c20a66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd50116501a06bcd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf992686e3119634c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5941e063b7c95c3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaa76e21e9bb620d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f17c3a8915ee18f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h271dc2ee49707f6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe3b2f379c351e06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3242bee849e3a0be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc35d13c4322e1d7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33f6199e744b5066;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1f62b8203ec4c20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d9e900e32d2375e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4232d4a308564f8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h572f52cdaec5ae1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91876e9f64ccc618;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5ea3d60ee78e975;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3e0ce2d55b8eb50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1726a68c3def6e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc033b303ac0b41d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7be14958dd41a233;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7514360e3529b8ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9265e263ac015de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf306c741c9de38ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h125ce07861be4284;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha65049e1a1604f1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had78f479898713;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb750570c78c579d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0c8cdbf6d9c582f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62684d600c42ab11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf8f77a1de4846b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3965af601bc8cf70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a17ec8dd50af3ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae101bc07950d7b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he40ab8d23c487bdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf367a869c00af191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d671b72208d160b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h511ea9aba7d41f4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b65add364d01f1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6de1ec038219041;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97bf80f36553745d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1eafc5a7be87ba1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8415d47e521e08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3424e33f906ca5b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b3698b79a20ba3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75876b79556e93ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h938537fab89d4225;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h485cd046c4de0bc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62d95c3780aca076;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he47cbd8268528bf4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2004a4e9095c2a60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9256e5643070bcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc03833ec48a2cee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52071bf351bfcc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec54bdc75921e637;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9d965c2ed7b0914;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h799696f3ac759220;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h804feed558764fde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4424bf567f4abdf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1890a1bafc82a431;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4fa889ef4fcbb38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7f8547457b0d95e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdefb95b9e2457e37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e42fd9995fccac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a39e3ce3b2f24e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac8f3466a164ea10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb846135b6d8b3823;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf04a718246e7412;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d818d8a1b6603ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30805d514898268a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31ce15da98395d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7b04bf5c31dc129;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45073ba8c457e5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb99d42c2f26faad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffa87938f4629303;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bf8305027c5367f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0ba892b66f983f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h311f32b3d9706bc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc54b35ff16f8e803;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf60f67f8a4458fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb94e2a83c7e2890;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb994606a2255e5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e6ddc5343027cbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed5e34b1c23a426c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6b840e986c48bbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ee94df9ee827239;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f865d9e1491d7c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83783d7490877aff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he53a0db875b318a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5090528833428a36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3cc6deb85b9bebf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7732edafa1f53127;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1217957275cc6998;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a6c8b6ced36fc11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9954ee1f083636e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96df69992a61afd9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21dcfd6df36b3d10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc638421b113362a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89577dfb52cfce4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56adb4c67d12425a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4b152a4947dc1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha86e438b906fbe84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h735c49b7f375af92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he28f466ee1ab4263;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20eed556504d73a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd871b5aa73488ba6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcad9031e29f3ae03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd32becd46058b016;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he468028e2f27ed61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8ce62efb10e3a25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b0e04f39e9cbd19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fd460c70ed9fa6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27a7c5085d05b4b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca456a1379c5c2b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e3ce19978d525ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfe79e20cf9ee844;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85f36616eb141e39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h641e2cd2ee160455;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f4c471a30f273db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h292d7360cb22b57b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe7d9757620a56e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41db9428e48ef515;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c65ab0eed682378;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff8e758bf93d2f37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he379b5c6c6dabbbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c0d39b9c5b312d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8107e1baffe67ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9823ac59076093f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0697ebc6a782a3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6535803e9605629;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde46a9b111c341cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9773fad6a76cd798;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd999e836a84a0cb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95da711c9c567199;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heda5b3f5c3eb8611;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b07dd641ebb9b1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40735824d6e1d13d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b3857edccbc51e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab2b1d783fa26c24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f9765a655ee2660;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b97dfe9f757d40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8de5d79bc1fdd93c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35059b3c72281b85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71e5e31c5addd188;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6dfaf549cfa559b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82a1fc67a07f40a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f9f628fe82d3017;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6921ae29540d8491;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h372bd190451995ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff8c05abd21618e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7d80928e218473d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22dec28169ddf8a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e0599d015d4cec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5807da2013ed8819;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3beffc345ed886ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cd4d8412e0056f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba8b56d44d385d2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb508bbc68406f7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a6bb4e62c81462c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ca3b01818eab848;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34f0388ce414656e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58475abbd321d5f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h424d215fecba9cbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14037bcf772aa659;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he78b397668e25969;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd39e7a430df0e914;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb81c24313241dc6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h960427a17ca21836;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2133d9c2af73c73c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fcfee384b8dd86c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7daffdd2519f6e7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4db869411a62ec7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24757e61cb95d2b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f644d51bca2098c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf71a6c8b44127dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e20b2c0a00b4cea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h680046cf6103d54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc98264e215a96c3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9283ccbe24fb1c73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6773214bbe2019de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7c53765451dc19f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ea9c51465c2bd93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dae6a42f670ade9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h834c5452ee5431d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dee29e9735e0b82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19c464eba036c735;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20c0eb89c4198ea0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99315ff4dc7533c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h280efd9e546251aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ecb80aa618910de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c24411c814b66d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1878e876c60c2ab4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb21a06a82ff20e72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4b50f0c551b3ab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b1e1970364bc371;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6631161ed6dca2e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c25d01874640f90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he960ad2d7ba52609;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5bb8397bd7a3919c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he73bf4de59790343;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3c88b1aab67efeb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7a94dcf1af591c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h159ba40e2b8774f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1c09838d6f7d40f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5504639f87beee6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e563f06cbb587ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb322fa4b76074;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84497efb2baa6e88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h787cf985c5ad8e5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2566aa31ff9ec8da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9029c511086846c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f34c2f83c814de2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92c3d42961abe911;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha277ce04ea30405c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0573f5bc5e9f646;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8fccf08596e505c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad7f9251ee643fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha28506e094ba0fee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdeb99547dde540f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bbd6554f6380bdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9ab365ae0d8e134;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12429779564916d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41a9f907bf4d60cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h547744268dc4ed55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ed449048aeac731;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h747392f777f91d06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h717a8e7f795c29d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde060d9bc373cc7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4f8c517d4b51bf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbd01a848de91de2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2b86b6fcbc6f2e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha554988ef3afbd00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d55bd9d2181e7fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaf4ba7807f7a593;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a204c4840437949;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f47c20b8ea8866a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac271060e38273bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9aef4c7eb99141a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6f9cbcb445d289a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf35976a41d091c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h683070a67a94e89a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5f781692a6ef0e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3769557913d2824b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7831ecdb5c455f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a06f04c070d98a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf687f67494e130ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52ac208c242531a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22634bc75b59cfea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h763a358463e0ac8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4feb26d34a41e1c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h939e5c45adf15141;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c108b797624df2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8ecd1296512f8cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73bfc686bac1c5b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd96bcedcd8db79b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he68d0001b645e018;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf21c756b93f5ad7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dfacedc4ca28ad0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h712af64e6fb17eda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e19061698a9aaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h196fff1b5c264b43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda13a7b891fe5396;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf83e0a792571741;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a2763b242a4978;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd6b5592666f6bf9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc381c8eb8e5e111;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd04b60b8e47599fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb103529c4de52ce6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h110698c1a90c1ce9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef97e9d55f22ce0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha20f4a676da202c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57413865ddbd7464;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2aaad2bd891dd0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45cd9f8d52e967e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haeaad94d534cb03e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf614814e88f9c485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h363bb2d9aa38d95c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12d4167bc8ec29fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbce6fe1f490ee7d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h393fabba5873d6bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8879329ed4af4b56;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae479612b4f9130;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha43ef42bb8fb77d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13516fd478ef5d32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ec6e79b479072cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7364b36937eeb53d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23b748cef1b590cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b10597385f70eb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80edae3fac0bf393;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h852f94e65c0ac717;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h397931a7d8e1308;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10295d99215da5e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6e5ea5d6623d272;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f55b10075289b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfba6f89cd18afdb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16c2e9eb2b7b9149;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc75222a1b979e819;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b220e94485c4b8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb988dc4c615b9d90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16fe1a8f2e86d87f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9be25b4dbaee5c6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6416925fcd8d63a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf692bd68e71eeaec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38b6cf6806db9e59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6709b56f191f0e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5569e283208e3960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ff2c94fef9b9e57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aea1114256221c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc865f64e4d4ad7a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h175d8c88a156d285;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc127120d4fa8242;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h385d7088bea5b73a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heede9dcda08bcd73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12a6f845baaec00f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h743a8677f3be677;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33bb85a5f8d28ded;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c4deebecbc24e85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8795d9015ad66092;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha28c06ff1e486d83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h893eb8149dacb027;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebe08311e38bdafe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28f69937ca02168e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedab691fb5b1d590;
        #1
        $finish();
    end
endmodule
