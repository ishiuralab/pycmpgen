module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    compressor_CLA162_32 compressor_CLA162_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA162_32(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [49:0] stage1_0;
   wire [55:0] stage1_1;
   wire [55:0] stage1_2;
   wire [75:0] stage1_3;
   wire [94:0] stage1_4;
   wire [53:0] stage1_5;
   wire [105:0] stage1_6;
   wire [65:0] stage1_7;
   wire [53:0] stage1_8;
   wire [76:0] stage1_9;
   wire [92:0] stage1_10;
   wire [66:0] stage1_11;
   wire [55:0] stage1_12;
   wire [85:0] stage1_13;
   wire [68:0] stage1_14;
   wire [59:0] stage1_15;
   wire [106:0] stage1_16;
   wire [63:0] stage1_17;
   wire [81:0] stage1_18;
   wire [66:0] stage1_19;
   wire [60:0] stage1_20;
   wire [79:0] stage1_21;
   wire [81:0] stage1_22;
   wire [90:0] stage1_23;
   wire [66:0] stage1_24;
   wire [77:0] stage1_25;
   wire [54:0] stage1_26;
   wire [66:0] stage1_27;
   wire [77:0] stage1_28;
   wire [74:0] stage1_29;
   wire [62:0] stage1_30;
   wire [97:0] stage1_31;
   wire [44:0] stage1_32;
   wire [18:0] stage1_33;
   wire [10:0] stage2_0;
   wire [16:0] stage2_1;
   wire [16:0] stage2_2;
   wire [34:0] stage2_3;
   wire [40:0] stage2_4;
   wire [27:0] stage2_5;
   wire [30:0] stage2_6;
   wire [33:0] stage2_7;
   wire [32:0] stage2_8;
   wire [31:0] stage2_9;
   wire [45:0] stage2_10;
   wire [38:0] stage2_11;
   wire [23:0] stage2_12;
   wire [44:0] stage2_13;
   wire [36:0] stage2_14;
   wire [33:0] stage2_15;
   wire [43:0] stage2_16;
   wire [36:0] stage2_17;
   wire [28:0] stage2_18;
   wire [27:0] stage2_19;
   wire [37:0] stage2_20;
   wire [27:0] stage2_21;
   wire [33:0] stage2_22;
   wire [43:0] stage2_23;
   wire [34:0] stage2_24;
   wire [30:0] stage2_25;
   wire [30:0] stage2_26;
   wire [32:0] stage2_27;
   wire [29:0] stage2_28;
   wire [32:0] stage2_29;
   wire [36:0] stage2_30;
   wire [35:0] stage2_31;
   wire [40:0] stage2_32;
   wire [23:0] stage2_33;
   wire [6:0] stage2_34;
   wire [1:0] stage2_35;
   wire [6:0] stage3_0;
   wire [9:0] stage3_1;
   wire [9:0] stage3_2;
   wire [22:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [16:0] stage3_6;
   wire [18:0] stage3_7;
   wire [17:0] stage3_8;
   wire [18:0] stage3_9;
   wire [14:0] stage3_10;
   wire [14:0] stage3_11;
   wire [14:0] stage3_12;
   wire [17:0] stage3_13;
   wire [16:0] stage3_14;
   wire [15:0] stage3_15;
   wire [12:0] stage3_16;
   wire [16:0] stage3_17;
   wire [16:0] stage3_18;
   wire [11:0] stage3_19;
   wire [17:0] stage3_20;
   wire [14:0] stage3_21;
   wire [22:0] stage3_22;
   wire [12:0] stage3_23;
   wire [16:0] stage3_24;
   wire [16:0] stage3_25;
   wire [11:0] stage3_26;
   wire [12:0] stage3_27;
   wire [22:0] stage3_28;
   wire [10:0] stage3_29;
   wire [13:0] stage3_30;
   wire [16:0] stage3_31;
   wire [15:0] stage3_32;
   wire [16:0] stage3_33;
   wire [15:0] stage3_34;
   wire [4:0] stage3_35;
   wire [1:0] stage4_0;
   wire [5:0] stage4_1;
   wire [5:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [7:0] stage4_9;
   wire [7:0] stage4_10;
   wire [9:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [5:0] stage4_14;
   wire [9:0] stage4_15;
   wire [6:0] stage4_16;
   wire [12:0] stage4_17;
   wire [8:0] stage4_18;
   wire [11:0] stage4_19;
   wire [5:0] stage4_20;
   wire [5:0] stage4_21;
   wire [8:0] stage4_22;
   wire [6:0] stage4_23;
   wire [7:0] stage4_24;
   wire [8:0] stage4_25;
   wire [8:0] stage4_26;
   wire [4:0] stage4_27;
   wire [8:0] stage4_28;
   wire [5:0] stage4_29;
   wire [5:0] stage4_30;
   wire [5:0] stage4_31;
   wire [10:0] stage4_32;
   wire [7:0] stage4_33;
   wire [8:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [3:0] stage5_3;
   wire [1:0] stage5_4;
   wire [4:0] stage5_5;
   wire [1:0] stage5_6;
   wire [6:0] stage5_7;
   wire [2:0] stage5_8;
   wire [2:0] stage5_9;
   wire [3:0] stage5_10;
   wire [5:0] stage5_11;
   wire [2:0] stage5_12;
   wire [2:0] stage5_13;
   wire [5:0] stage5_14;
   wire [5:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [4:0] stage5_18;
   wire [2:0] stage5_19;
   wire [3:0] stage5_20;
   wire [4:0] stage5_21;
   wire [1:0] stage5_22;
   wire [3:0] stage5_23;
   wire [5:0] stage5_24;
   wire [1:0] stage5_25;
   wire [3:0] stage5_26;
   wire [3:0] stage5_27;
   wire [3:0] stage5_28;
   wire [5:0] stage5_29;
   wire [2:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [4:0] stage5_33;
   wire [3:0] stage5_34;
   wire [5:0] stage5_35;
   wire [3:0] stage5_36;
   wire [0:0] stage5_37;
   wire [0:0] stage5_38;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [1:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[0],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[1],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[2],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59]},
      {stage1_5[3],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65]},
      {stage1_5[4],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage1_5[5],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc615_5 gpc38 (
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76]},
      {stage0_3[72]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[6],stage1_4[38],stage1_3[38],stage1_2[38]}
   );
   gpc615_5 gpc39 (
      {stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage0_3[73]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[7],stage1_4[39],stage1_3[39],stage1_2[39]}
   );
   gpc615_5 gpc40 (
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage0_3[74]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[8],stage1_4[40],stage1_3[40],stage1_2[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage0_3[75]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[9],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc615_5 gpc42 (
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage0_3[76]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[10],stage1_4[42],stage1_3[42],stage1_2[42]}
   );
   gpc615_5 gpc43 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage0_3[77]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[11],stage1_4[43],stage1_3[43],stage1_2[43]}
   );
   gpc615_5 gpc44 (
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106]},
      {stage0_3[78]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[12],stage1_4[44],stage1_3[44],stage1_2[44]}
   );
   gpc615_5 gpc45 (
      {stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage0_3[79]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[13],stage1_4[45],stage1_3[45],stage1_2[45]}
   );
   gpc615_5 gpc46 (
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage0_3[80]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[14],stage1_4[46],stage1_3[46],stage1_2[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_3[81]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[15],stage1_4[47],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage0_3[82]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[16],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage0_3[83]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[17],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136]},
      {stage0_3[84]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[18],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage0_3[85]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[19],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage0_3[86]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[20],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_3[87]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[21],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc615_5 gpc54 (
      {stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage0_3[88]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[22],stage1_4[54],stage1_3[54],stage1_2[54]}
   );
   gpc615_5 gpc55 (
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage0_3[89]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[23],stage1_4[55],stage1_3[55],stage1_2[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage0_4[108]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[18],stage1_5[24],stage1_4[56],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage0_4[109]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[19],stage1_5[25],stage1_4[57],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage0_4[110]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[20],stage1_5[26],stage1_4[58],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage0_4[111]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[21],stage1_5[27],stage1_4[59],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage0_4[112]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[22],stage1_5[28],stage1_4[60],stage1_3[60]}
   );
   gpc615_5 gpc61 (
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119]},
      {stage0_4[113]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[23],stage1_5[29],stage1_4[61],stage1_3[61]}
   );
   gpc615_5 gpc62 (
      {stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage0_4[114]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[24],stage1_5[30],stage1_4[62],stage1_3[62]}
   );
   gpc615_5 gpc63 (
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage0_4[115]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[25],stage1_5[31],stage1_4[63],stage1_3[63]}
   );
   gpc615_5 gpc64 (
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage0_4[116]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[26],stage1_5[32],stage1_4[64],stage1_3[64]}
   );
   gpc615_5 gpc65 (
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage0_4[117]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[27],stage1_5[33],stage1_4[65],stage1_3[65]}
   );
   gpc615_5 gpc66 (
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage0_4[118]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[28],stage1_5[34],stage1_4[66],stage1_3[66]}
   );
   gpc615_5 gpc67 (
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage0_4[119]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[29],stage1_5[35],stage1_4[67],stage1_3[67]}
   );
   gpc615_5 gpc68 (
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage0_4[120]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[30],stage1_5[36],stage1_4[68],stage1_3[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[13],stage1_6[31],stage1_5[37],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[14],stage1_6[32],stage1_5[38],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[15],stage1_6[33],stage1_5[39],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[16],stage1_6[34],stage1_5[40]}
   );
   gpc606_5 gpc73 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[17],stage1_6[35],stage1_5[41]}
   );
   gpc606_5 gpc74 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[18],stage1_6[36],stage1_5[42]}
   );
   gpc606_5 gpc75 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[19],stage1_6[37],stage1_5[43]}
   );
   gpc606_5 gpc76 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[7],stage1_7[20],stage1_6[38],stage1_5[44]}
   );
   gpc606_5 gpc77 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[8],stage1_7[21],stage1_6[39],stage1_5[45]}
   );
   gpc606_5 gpc78 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[9],stage1_7[22],stage1_6[40],stage1_5[46]}
   );
   gpc606_5 gpc79 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[10],stage1_7[23],stage1_6[41],stage1_5[47]}
   );
   gpc606_5 gpc80 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[11],stage1_7[24],stage1_6[42],stage1_5[48]}
   );
   gpc606_5 gpc81 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[12],stage1_7[25],stage1_6[43],stage1_5[49]}
   );
   gpc606_5 gpc82 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[13],stage1_7[26],stage1_6[44],stage1_5[50]}
   );
   gpc606_5 gpc83 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[14],stage1_7[27],stage1_6[45],stage1_5[51]}
   );
   gpc606_5 gpc84 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[15],stage1_7[28],stage1_6[46],stage1_5[52]}
   );
   gpc606_5 gpc85 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[16],stage1_7[29],stage1_6[47],stage1_5[53]}
   );
   gpc606_5 gpc86 (
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[14],stage1_8[17],stage1_7[30],stage1_6[48]}
   );
   gpc606_5 gpc87 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[15],stage1_8[18],stage1_7[31],stage1_6[49]}
   );
   gpc606_5 gpc88 (
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[16],stage1_8[19],stage1_7[32],stage1_6[50]}
   );
   gpc606_5 gpc89 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[17],stage1_8[20],stage1_7[33],stage1_6[51]}
   );
   gpc606_5 gpc90 (
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[18],stage1_8[21],stage1_7[34],stage1_6[52]}
   );
   gpc606_5 gpc91 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[19],stage1_8[22],stage1_7[35],stage1_6[53]}
   );
   gpc615_5 gpc92 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[84]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[20],stage1_8[23],stage1_7[36],stage1_6[54]}
   );
   gpc615_5 gpc93 (
      {stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_7[85]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[21],stage1_8[24],stage1_7[37],stage1_6[55]}
   );
   gpc615_5 gpc94 (
      {stage0_6[64], stage0_6[65], stage0_6[66], stage0_6[67], stage0_6[68]},
      {stage0_7[86]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[22],stage1_8[25],stage1_7[38],stage1_6[56]}
   );
   gpc615_5 gpc95 (
      {stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72], stage0_6[73]},
      {stage0_7[87]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[23],stage1_8[26],stage1_7[39],stage1_6[57]}
   );
   gpc615_5 gpc96 (
      {stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage0_7[88]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[24],stage1_8[27],stage1_7[40],stage1_6[58]}
   );
   gpc615_5 gpc97 (
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage0_7[89]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[25],stage1_8[28],stage1_7[41],stage1_6[59]}
   );
   gpc615_5 gpc98 (
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88]},
      {stage0_7[90]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[26],stage1_8[29],stage1_7[42],stage1_6[60]}
   );
   gpc615_5 gpc99 (
      {stage0_6[89], stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93]},
      {stage0_7[91]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[27],stage1_8[30],stage1_7[43],stage1_6[61]}
   );
   gpc615_5 gpc100 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98]},
      {stage0_7[92]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[28],stage1_8[31],stage1_7[44],stage1_6[62]}
   );
   gpc615_5 gpc101 (
      {stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103]},
      {stage0_7[93]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[29],stage1_8[32],stage1_7[45],stage1_6[63]}
   );
   gpc615_5 gpc102 (
      {stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage0_7[94]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[30],stage1_8[33],stage1_7[46],stage1_6[64]}
   );
   gpc615_5 gpc103 (
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage0_7[95]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[31],stage1_8[34],stage1_7[47],stage1_6[65]}
   );
   gpc615_5 gpc104 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[96]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[32],stage1_8[35],stage1_7[48],stage1_6[66]}
   );
   gpc615_5 gpc105 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[97]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[33],stage1_8[36],stage1_7[49],stage1_6[67]}
   );
   gpc615_5 gpc106 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[120]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[20],stage1_9[34],stage1_8[37],stage1_7[50]}
   );
   gpc615_5 gpc107 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[121]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[21],stage1_9[35],stage1_8[38],stage1_7[51]}
   );
   gpc615_5 gpc108 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[122]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[22],stage1_9[36],stage1_8[39],stage1_7[52]}
   );
   gpc615_5 gpc109 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[123]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[23],stage1_9[37],stage1_8[40],stage1_7[53]}
   );
   gpc615_5 gpc110 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[124]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[24],stage1_9[38],stage1_8[41],stage1_7[54]}
   );
   gpc615_5 gpc111 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[125]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[25],stage1_9[39],stage1_8[42],stage1_7[55]}
   );
   gpc615_5 gpc112 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[126]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[26],stage1_9[40],stage1_8[43],stage1_7[56]}
   );
   gpc615_5 gpc113 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[127]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[27],stage1_9[41],stage1_8[44],stage1_7[57]}
   );
   gpc615_5 gpc114 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[128]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[28],stage1_9[42],stage1_8[45],stage1_7[58]}
   );
   gpc615_5 gpc115 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[129]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[29],stage1_9[43],stage1_8[46],stage1_7[59]}
   );
   gpc615_5 gpc116 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[130]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[30],stage1_9[44],stage1_8[47],stage1_7[60]}
   );
   gpc615_5 gpc117 (
      {stage0_7[153], stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157]},
      {stage0_8[131]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[31],stage1_9[45],stage1_8[48],stage1_7[61]}
   );
   gpc606_5 gpc118 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[12],stage1_10[32],stage1_9[46],stage1_8[49]}
   );
   gpc606_5 gpc119 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[13],stage1_10[33],stage1_9[47],stage1_8[50]}
   );
   gpc606_5 gpc120 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[14],stage1_10[34],stage1_9[48],stage1_8[51]}
   );
   gpc606_5 gpc121 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[15],stage1_10[35],stage1_9[49],stage1_8[52]}
   );
   gpc606_5 gpc122 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[16],stage1_10[36],stage1_9[50],stage1_8[53]}
   );
   gpc615_5 gpc123 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76]},
      {stage0_10[30]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[5],stage1_11[17],stage1_10[37],stage1_9[51]}
   );
   gpc615_5 gpc124 (
      {stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_10[31]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[6],stage1_11[18],stage1_10[38],stage1_9[52]}
   );
   gpc615_5 gpc125 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_10[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[7],stage1_11[19],stage1_10[39],stage1_9[53]}
   );
   gpc615_5 gpc126 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_10[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[8],stage1_11[20],stage1_10[40],stage1_9[54]}
   );
   gpc615_5 gpc127 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96]},
      {stage0_10[34]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[9],stage1_11[21],stage1_10[41],stage1_9[55]}
   );
   gpc615_5 gpc128 (
      {stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_10[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[10],stage1_11[22],stage1_10[42],stage1_9[56]}
   );
   gpc615_5 gpc129 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106]},
      {stage0_10[36]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[11],stage1_11[23],stage1_10[43],stage1_9[57]}
   );
   gpc615_5 gpc130 (
      {stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_10[37]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[12],stage1_11[24],stage1_10[44],stage1_9[58]}
   );
   gpc615_5 gpc131 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_10[38]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[13],stage1_11[25],stage1_10[45],stage1_9[59]}
   );
   gpc615_5 gpc132 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_10[39]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[14],stage1_11[26],stage1_10[46],stage1_9[60]}
   );
   gpc615_5 gpc133 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_10[40]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[15],stage1_11[27],stage1_10[47],stage1_9[61]}
   );
   gpc615_5 gpc134 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_10[41]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[16],stage1_11[28],stage1_10[48],stage1_9[62]}
   );
   gpc615_5 gpc135 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136]},
      {stage0_10[42]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[17],stage1_11[29],stage1_10[49],stage1_9[63]}
   );
   gpc615_5 gpc136 (
      {stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141]},
      {stage0_10[43]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[18],stage1_11[30],stage1_10[50],stage1_9[64]}
   );
   gpc615_5 gpc137 (
      {stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_10[44]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[19],stage1_11[31],stage1_10[51],stage1_9[65]}
   );
   gpc615_5 gpc138 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[45]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[20],stage1_11[32],stage1_10[52],stage1_9[66]}
   );
   gpc615_5 gpc139 (
      {stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50]},
      {stage0_11[96]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[16],stage1_12[21],stage1_11[33],stage1_10[53]}
   );
   gpc615_5 gpc140 (
      {stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54], stage0_10[55]},
      {stage0_11[97]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[17],stage1_12[22],stage1_11[34],stage1_10[54]}
   );
   gpc615_5 gpc141 (
      {stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60]},
      {stage0_11[98]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[18],stage1_12[23],stage1_11[35],stage1_10[55]}
   );
   gpc615_5 gpc142 (
      {stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage0_11[99]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[19],stage1_12[24],stage1_11[36],stage1_10[56]}
   );
   gpc615_5 gpc143 (
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70]},
      {stage0_11[100]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[20],stage1_12[25],stage1_11[37],stage1_10[57]}
   );
   gpc615_5 gpc144 (
      {stage0_10[71], stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75]},
      {stage0_11[101]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[21],stage1_12[26],stage1_11[38],stage1_10[58]}
   );
   gpc615_5 gpc145 (
      {stage0_10[76], stage0_10[77], stage0_10[78], stage0_10[79], stage0_10[80]},
      {stage0_11[102]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[22],stage1_12[27],stage1_11[39],stage1_10[59]}
   );
   gpc615_5 gpc146 (
      {stage0_10[81], stage0_10[82], stage0_10[83], stage0_10[84], stage0_10[85]},
      {stage0_11[103]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[23],stage1_12[28],stage1_11[40],stage1_10[60]}
   );
   gpc615_5 gpc147 (
      {stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89], stage0_10[90]},
      {stage0_11[104]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[24],stage1_12[29],stage1_11[41],stage1_10[61]}
   );
   gpc615_5 gpc148 (
      {stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_11[105]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[25],stage1_12[30],stage1_11[42],stage1_10[62]}
   );
   gpc615_5 gpc149 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100]},
      {stage0_11[106]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[26],stage1_12[31],stage1_11[43],stage1_10[63]}
   );
   gpc615_5 gpc150 (
      {stage0_10[101], stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105]},
      {stage0_11[107]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[27],stage1_12[32],stage1_11[44],stage1_10[64]}
   );
   gpc615_5 gpc151 (
      {stage0_10[106], stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110]},
      {stage0_11[108]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[28],stage1_12[33],stage1_11[45],stage1_10[65]}
   );
   gpc615_5 gpc152 (
      {stage0_10[111], stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115]},
      {stage0_11[109]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[29],stage1_12[34],stage1_11[46],stage1_10[66]}
   );
   gpc615_5 gpc153 (
      {stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120]},
      {stage0_11[110]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[30],stage1_12[35],stage1_11[47],stage1_10[67]}
   );
   gpc615_5 gpc154 (
      {stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage0_11[111]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[31],stage1_12[36],stage1_11[48],stage1_10[68]}
   );
   gpc615_5 gpc155 (
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130]},
      {stage0_11[112]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[32],stage1_12[37],stage1_11[49],stage1_10[69]}
   );
   gpc615_5 gpc156 (
      {stage0_10[131], stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135]},
      {stage0_11[113]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[33],stage1_12[38],stage1_11[50],stage1_10[70]}
   );
   gpc615_5 gpc157 (
      {stage0_10[136], stage0_10[137], stage0_10[138], stage0_10[139], stage0_10[140]},
      {stage0_11[114]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[34],stage1_12[39],stage1_11[51],stage1_10[71]}
   );
   gpc615_5 gpc158 (
      {stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage0_12[114]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[19],stage1_13[35],stage1_12[40],stage1_11[52]}
   );
   gpc615_5 gpc159 (
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124]},
      {stage0_12[115]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[20],stage1_13[36],stage1_12[41],stage1_11[53]}
   );
   gpc615_5 gpc160 (
      {stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage0_12[116]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[21],stage1_13[37],stage1_12[42],stage1_11[54]}
   );
   gpc615_5 gpc161 (
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134]},
      {stage0_12[117]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[22],stage1_13[38],stage1_12[43],stage1_11[55]}
   );
   gpc615_5 gpc162 (
      {stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139]},
      {stage0_12[118]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[23],stage1_13[39],stage1_12[44],stage1_11[56]}
   );
   gpc615_5 gpc163 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[119]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[24],stage1_13[40],stage1_12[45],stage1_11[57]}
   );
   gpc615_5 gpc164 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[120]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[25],stage1_13[41],stage1_12[46],stage1_11[58]}
   );
   gpc615_5 gpc165 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[121]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[26],stage1_13[42],stage1_12[47],stage1_11[59]}
   );
   gpc615_5 gpc166 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126]},
      {stage0_13[48]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[8],stage1_14[27],stage1_13[43],stage1_12[48]}
   );
   gpc615_5 gpc167 (
      {stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_13[49]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[9],stage1_14[28],stage1_13[44],stage1_12[49]}
   );
   gpc615_5 gpc168 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136]},
      {stage0_13[50]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[10],stage1_14[29],stage1_13[45],stage1_12[50]}
   );
   gpc615_5 gpc169 (
      {stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage0_13[51]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[11],stage1_14[30],stage1_13[46],stage1_12[51]}
   );
   gpc615_5 gpc170 (
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_13[52]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[12],stage1_14[31],stage1_13[47],stage1_12[52]}
   );
   gpc615_5 gpc171 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_13[53]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[13],stage1_14[32],stage1_13[48],stage1_12[53]}
   );
   gpc615_5 gpc172 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156]},
      {stage0_13[54]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[14],stage1_14[33],stage1_13[49],stage1_12[54]}
   );
   gpc615_5 gpc173 (
      {stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_13[55]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[15],stage1_14[34],stage1_13[50],stage1_12[55]}
   );
   gpc606_5 gpc174 (
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[8],stage1_15[16],stage1_14[35],stage1_13[51]}
   );
   gpc606_5 gpc175 (
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[9],stage1_15[17],stage1_14[36],stage1_13[52]}
   );
   gpc606_5 gpc176 (
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[10],stage1_15[18],stage1_14[37],stage1_13[53]}
   );
   gpc615_5 gpc177 (
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78]},
      {stage0_14[48]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[11],stage1_15[19],stage1_14[38],stage1_13[54]}
   );
   gpc615_5 gpc178 (
      {stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_14[49]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[12],stage1_15[20],stage1_14[39],stage1_13[55]}
   );
   gpc615_5 gpc179 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88]},
      {stage0_14[50]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[13],stage1_15[21],stage1_14[40],stage1_13[56]}
   );
   gpc615_5 gpc180 (
      {stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_14[51]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[14],stage1_15[22],stage1_14[41],stage1_13[57]}
   );
   gpc615_5 gpc181 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98]},
      {stage0_14[52]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[15],stage1_15[23],stage1_14[42],stage1_13[58]}
   );
   gpc615_5 gpc182 (
      {stage0_13[99], stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103]},
      {stage0_14[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[16],stage1_15[24],stage1_14[43],stage1_13[59]}
   );
   gpc615_5 gpc183 (
      {stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108]},
      {stage0_14[54]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[17],stage1_15[25],stage1_14[44],stage1_13[60]}
   );
   gpc615_5 gpc184 (
      {stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_14[55]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[18],stage1_15[26],stage1_14[45],stage1_13[61]}
   );
   gpc615_5 gpc185 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118]},
      {stage0_14[56]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[19],stage1_15[27],stage1_14[46],stage1_13[62]}
   );
   gpc615_5 gpc186 (
      {stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_14[57]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[20],stage1_15[28],stage1_14[47],stage1_13[63]}
   );
   gpc615_5 gpc187 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128]},
      {stage0_14[58]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[21],stage1_15[29],stage1_14[48],stage1_13[64]}
   );
   gpc615_5 gpc188 (
      {stage0_13[129], stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133]},
      {stage0_14[59]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[22],stage1_15[30],stage1_14[49],stage1_13[65]}
   );
   gpc615_5 gpc189 (
      {stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138]},
      {stage0_14[60]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[23],stage1_15[31],stage1_14[50],stage1_13[66]}
   );
   gpc615_5 gpc190 (
      {stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_14[61]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[24],stage1_15[32],stage1_14[51],stage1_13[67]}
   );
   gpc117_4 gpc191 (
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67], stage0_14[68]},
      {stage0_15[102]},
      {stage0_16[0]},
      {stage1_17[17],stage1_16[25],stage1_15[33],stage1_14[52]}
   );
   gpc117_4 gpc192 (
      {stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75]},
      {stage0_15[103]},
      {stage0_16[1]},
      {stage1_17[18],stage1_16[26],stage1_15[34],stage1_14[53]}
   );
   gpc117_4 gpc193 (
      {stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82]},
      {stage0_15[104]},
      {stage0_16[2]},
      {stage1_17[19],stage1_16[27],stage1_15[35],stage1_14[54]}
   );
   gpc117_4 gpc194 (
      {stage0_14[83], stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage0_15[105]},
      {stage0_16[3]},
      {stage1_17[20],stage1_16[28],stage1_15[36],stage1_14[55]}
   );
   gpc606_5 gpc195 (
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9]},
      {stage1_18[0],stage1_17[21],stage1_16[29],stage1_15[37],stage1_14[56]}
   );
   gpc606_5 gpc196 (
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15]},
      {stage1_18[1],stage1_17[22],stage1_16[30],stage1_15[38],stage1_14[57]}
   );
   gpc606_5 gpc197 (
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21]},
      {stage1_18[2],stage1_17[23],stage1_16[31],stage1_15[39],stage1_14[58]}
   );
   gpc606_5 gpc198 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27]},
      {stage1_18[3],stage1_17[24],stage1_16[32],stage1_15[40],stage1_14[59]}
   );
   gpc606_5 gpc199 (
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33]},
      {stage1_18[4],stage1_17[25],stage1_16[33],stage1_15[41],stage1_14[60]}
   );
   gpc606_5 gpc200 (
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39]},
      {stage1_18[5],stage1_17[26],stage1_16[34],stage1_15[42],stage1_14[61]}
   );
   gpc606_5 gpc201 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45]},
      {stage1_18[6],stage1_17[27],stage1_16[35],stage1_15[43],stage1_14[62]}
   );
   gpc606_5 gpc202 (
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51]},
      {stage1_18[7],stage1_17[28],stage1_16[36],stage1_15[44],stage1_14[63]}
   );
   gpc606_5 gpc203 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage1_18[8],stage1_17[29],stage1_16[37],stage1_15[45],stage1_14[64]}
   );
   gpc606_5 gpc204 (
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63]},
      {stage1_18[9],stage1_17[30],stage1_16[38],stage1_15[46],stage1_14[65]}
   );
   gpc606_5 gpc205 (
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69]},
      {stage1_18[10],stage1_17[31],stage1_16[39],stage1_15[47],stage1_14[66]}
   );
   gpc615_5 gpc206 (
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160]},
      {stage0_15[106]},
      {stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75]},
      {stage1_18[11],stage1_17[32],stage1_16[40],stage1_15[48],stage1_14[67]}
   );
   gpc615_5 gpc207 (
      {stage0_15[107], stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111]},
      {stage0_16[76]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[12],stage1_17[33],stage1_16[41],stage1_15[49]}
   );
   gpc615_5 gpc208 (
      {stage0_15[112], stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116]},
      {stage0_16[77]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[13],stage1_17[34],stage1_16[42],stage1_15[50]}
   );
   gpc615_5 gpc209 (
      {stage0_15[117], stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121]},
      {stage0_16[78]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[14],stage1_17[35],stage1_16[43],stage1_15[51]}
   );
   gpc615_5 gpc210 (
      {stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126]},
      {stage0_16[79]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[15],stage1_17[36],stage1_16[44],stage1_15[52]}
   );
   gpc615_5 gpc211 (
      {stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage0_16[80]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[16],stage1_17[37],stage1_16[45],stage1_15[53]}
   );
   gpc615_5 gpc212 (
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136]},
      {stage0_16[81]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[17],stage1_17[38],stage1_16[46],stage1_15[54]}
   );
   gpc615_5 gpc213 (
      {stage0_15[137], stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141]},
      {stage0_16[82]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[18],stage1_17[39],stage1_16[47],stage1_15[55]}
   );
   gpc615_5 gpc214 (
      {stage0_15[142], stage0_15[143], stage0_15[144], stage0_15[145], stage0_15[146]},
      {stage0_16[83]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[19],stage1_17[40],stage1_16[48],stage1_15[56]}
   );
   gpc615_5 gpc215 (
      {stage0_15[147], stage0_15[148], stage0_15[149], stage0_15[150], stage0_15[151]},
      {stage0_16[84]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[20],stage1_17[41],stage1_16[49],stage1_15[57]}
   );
   gpc615_5 gpc216 (
      {stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155], stage0_15[156]},
      {stage0_16[85]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[21],stage1_17[42],stage1_16[50],stage1_15[58]}
   );
   gpc615_5 gpc217 (
      {stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage0_16[86]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[22],stage1_17[43],stage1_16[51],stage1_15[59]}
   );
   gpc606_5 gpc218 (
      {stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91], stage0_16[92]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[11],stage1_18[23],stage1_17[44],stage1_16[52]}
   );
   gpc606_5 gpc219 (
      {stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97], stage0_16[98]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[12],stage1_18[24],stage1_17[45],stage1_16[53]}
   );
   gpc606_5 gpc220 (
      {stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103], stage0_16[104]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[13],stage1_18[25],stage1_17[46],stage1_16[54]}
   );
   gpc606_5 gpc221 (
      {stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109], stage0_16[110]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[14],stage1_18[26],stage1_17[47],stage1_16[55]}
   );
   gpc606_5 gpc222 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[4],stage1_19[15],stage1_18[27],stage1_17[48]}
   );
   gpc606_5 gpc223 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[5],stage1_19[16],stage1_18[28],stage1_17[49]}
   );
   gpc606_5 gpc224 (
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[6],stage1_19[17],stage1_18[29],stage1_17[50]}
   );
   gpc606_5 gpc225 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[7],stage1_19[18],stage1_18[30],stage1_17[51]}
   );
   gpc606_5 gpc226 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[8],stage1_19[19],stage1_18[31],stage1_17[52]}
   );
   gpc606_5 gpc227 (
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[9],stage1_19[20],stage1_18[32],stage1_17[53]}
   );
   gpc606_5 gpc228 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[10],stage1_19[21],stage1_18[33],stage1_17[54]}
   );
   gpc606_5 gpc229 (
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[11],stage1_19[22],stage1_18[34],stage1_17[55]}
   );
   gpc606_5 gpc230 (
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[12],stage1_19[23],stage1_18[35],stage1_17[56]}
   );
   gpc606_5 gpc231 (
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[13],stage1_19[24],stage1_18[36],stage1_17[57]}
   );
   gpc606_5 gpc232 (
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[14],stage1_19[25],stage1_18[37],stage1_17[58]}
   );
   gpc606_5 gpc233 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[15],stage1_19[26],stage1_18[38],stage1_17[59]}
   );
   gpc606_5 gpc234 (
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[16],stage1_19[27],stage1_18[39],stage1_17[60]}
   );
   gpc606_5 gpc235 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[17],stage1_19[28],stage1_18[40],stage1_17[61]}
   );
   gpc606_5 gpc236 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[18],stage1_19[29],stage1_18[41],stage1_17[62]}
   );
   gpc606_5 gpc237 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[19],stage1_19[30],stage1_18[42],stage1_17[63]}
   );
   gpc117_4 gpc238 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29], stage0_18[30]},
      {stage0_19[96]},
      {stage0_20[0]},
      {stage1_21[16],stage1_20[20],stage1_19[31],stage1_18[43]}
   );
   gpc117_4 gpc239 (
      {stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35], stage0_18[36], stage0_18[37]},
      {stage0_19[97]},
      {stage0_20[1]},
      {stage1_21[17],stage1_20[21],stage1_19[32],stage1_18[44]}
   );
   gpc117_4 gpc240 (
      {stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41], stage0_18[42], stage0_18[43], stage0_18[44]},
      {stage0_19[98]},
      {stage0_20[2]},
      {stage1_21[18],stage1_20[22],stage1_19[33],stage1_18[45]}
   );
   gpc117_4 gpc241 (
      {stage0_18[45], stage0_18[46], stage0_18[47], stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51]},
      {stage0_19[99]},
      {stage0_20[3]},
      {stage1_21[19],stage1_20[23],stage1_19[34],stage1_18[46]}
   );
   gpc606_5 gpc242 (
      {stage0_18[52], stage0_18[53], stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57]},
      {stage0_20[4], stage0_20[5], stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9]},
      {stage1_22[0],stage1_21[20],stage1_20[24],stage1_19[35],stage1_18[47]}
   );
   gpc606_5 gpc243 (
      {stage0_18[58], stage0_18[59], stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63]},
      {stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15]},
      {stage1_22[1],stage1_21[21],stage1_20[25],stage1_19[36],stage1_18[48]}
   );
   gpc606_5 gpc244 (
      {stage0_18[64], stage0_18[65], stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69]},
      {stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21]},
      {stage1_22[2],stage1_21[22],stage1_20[26],stage1_19[37],stage1_18[49]}
   );
   gpc606_5 gpc245 (
      {stage0_18[70], stage0_18[71], stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75]},
      {stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage1_22[3],stage1_21[23],stage1_20[27],stage1_19[38],stage1_18[50]}
   );
   gpc606_5 gpc246 (
      {stage0_18[76], stage0_18[77], stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81]},
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage1_22[4],stage1_21[24],stage1_20[28],stage1_19[39],stage1_18[51]}
   );
   gpc606_5 gpc247 (
      {stage0_18[82], stage0_18[83], stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87]},
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39]},
      {stage1_22[5],stage1_21[25],stage1_20[29],stage1_19[40],stage1_18[52]}
   );
   gpc606_5 gpc248 (
      {stage0_18[88], stage0_18[89], stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93]},
      {stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45]},
      {stage1_22[6],stage1_21[26],stage1_20[30],stage1_19[41],stage1_18[53]}
   );
   gpc606_5 gpc249 (
      {stage0_18[94], stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99]},
      {stage0_20[46], stage0_20[47], stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51]},
      {stage1_22[7],stage1_21[27],stage1_20[31],stage1_19[42],stage1_18[54]}
   );
   gpc606_5 gpc250 (
      {stage0_18[100], stage0_18[101], stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105]},
      {stage0_20[52], stage0_20[53], stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57]},
      {stage1_22[8],stage1_21[28],stage1_20[32],stage1_19[43],stage1_18[55]}
   );
   gpc606_5 gpc251 (
      {stage0_18[106], stage0_18[107], stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111]},
      {stage0_20[58], stage0_20[59], stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63]},
      {stage1_22[9],stage1_21[29],stage1_20[33],stage1_19[44],stage1_18[56]}
   );
   gpc606_5 gpc252 (
      {stage0_18[112], stage0_18[113], stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117]},
      {stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage1_22[10],stage1_21[30],stage1_20[34],stage1_19[45],stage1_18[57]}
   );
   gpc606_5 gpc253 (
      {stage0_18[118], stage0_18[119], stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123]},
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75]},
      {stage1_22[11],stage1_21[31],stage1_20[35],stage1_19[46],stage1_18[58]}
   );
   gpc606_5 gpc254 (
      {stage0_18[124], stage0_18[125], stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129]},
      {stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81]},
      {stage1_22[12],stage1_21[32],stage1_20[36],stage1_19[47],stage1_18[59]}
   );
   gpc606_5 gpc255 (
      {stage0_18[130], stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87]},
      {stage1_22[13],stage1_21[33],stage1_20[37],stage1_19[48],stage1_18[60]}
   );
   gpc606_5 gpc256 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141]},
      {stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93]},
      {stage1_22[14],stage1_21[34],stage1_20[38],stage1_19[49],stage1_18[61]}
   );
   gpc606_5 gpc257 (
      {stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[15],stage1_21[35],stage1_20[39],stage1_19[50]}
   );
   gpc606_5 gpc258 (
      {stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[16],stage1_21[36],stage1_20[40],stage1_19[51]}
   );
   gpc606_5 gpc259 (
      {stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[17],stage1_21[37],stage1_20[41],stage1_19[52]}
   );
   gpc606_5 gpc260 (
      {stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[18],stage1_21[38],stage1_20[42],stage1_19[53]}
   );
   gpc606_5 gpc261 (
      {stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[19],stage1_21[39],stage1_20[43],stage1_19[54]}
   );
   gpc606_5 gpc262 (
      {stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[20],stage1_21[40],stage1_20[44],stage1_19[55]}
   );
   gpc606_5 gpc263 (
      {stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[21],stage1_21[41],stage1_20[45],stage1_19[56]}
   );
   gpc606_5 gpc264 (
      {stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[22],stage1_21[42],stage1_20[46],stage1_19[57]}
   );
   gpc606_5 gpc265 (
      {stage0_19[148], stage0_19[149], stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[23],stage1_21[43],stage1_20[47],stage1_19[58]}
   );
   gpc606_5 gpc266 (
      {stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[9],stage1_22[24],stage1_21[44],stage1_20[48]}
   );
   gpc606_5 gpc267 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[10],stage1_22[25],stage1_21[45],stage1_20[49]}
   );
   gpc606_5 gpc268 (
      {stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[11],stage1_22[26],stage1_21[46],stage1_20[50]}
   );
   gpc615_5 gpc269 (
      {stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_21[54]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[12],stage1_22[27],stage1_21[47],stage1_20[51]}
   );
   gpc615_5 gpc270 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_21[55]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[13],stage1_22[28],stage1_21[48],stage1_20[52]}
   );
   gpc615_5 gpc271 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126]},
      {stage0_21[56]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[14],stage1_22[29],stage1_21[49],stage1_20[53]}
   );
   gpc615_5 gpc272 (
      {stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_21[57]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[15],stage1_22[30],stage1_21[50],stage1_20[54]}
   );
   gpc615_5 gpc273 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136]},
      {stage0_21[58]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[16],stage1_22[31],stage1_21[51],stage1_20[55]}
   );
   gpc615_5 gpc274 (
      {stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141]},
      {stage0_21[59]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[17],stage1_22[32],stage1_21[52],stage1_20[56]}
   );
   gpc615_5 gpc275 (
      {stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_21[60]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[18],stage1_22[33],stage1_21[53],stage1_20[57]}
   );
   gpc615_5 gpc276 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_21[61]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[19],stage1_22[34],stage1_21[54],stage1_20[58]}
   );
   gpc615_5 gpc277 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156]},
      {stage0_21[62]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[20],stage1_22[35],stage1_21[55],stage1_20[59]}
   );
   gpc615_5 gpc278 (
      {stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_21[63]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[21],stage1_22[36],stage1_21[56],stage1_20[60]}
   );
   gpc1163_5 gpc279 (
      {stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage0_23[0]},
      {stage0_24[0]},
      {stage1_25[0],stage1_24[13],stage1_23[22],stage1_22[37],stage1_21[57]}
   );
   gpc1163_5 gpc280 (
      {stage0_21[67], stage0_21[68], stage0_21[69]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage0_23[1]},
      {stage0_24[1]},
      {stage1_25[1],stage1_24[14],stage1_23[23],stage1_22[38],stage1_21[58]}
   );
   gpc1163_5 gpc281 (
      {stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage0_23[2]},
      {stage0_24[2]},
      {stage1_25[2],stage1_24[15],stage1_23[24],stage1_22[39],stage1_21[59]}
   );
   gpc1163_5 gpc282 (
      {stage0_21[73], stage0_21[74], stage0_21[75]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage0_23[3]},
      {stage0_24[3]},
      {stage1_25[3],stage1_24[16],stage1_23[25],stage1_22[40],stage1_21[60]}
   );
   gpc1163_5 gpc283 (
      {stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage0_23[4]},
      {stage0_24[4]},
      {stage1_25[4],stage1_24[17],stage1_23[26],stage1_22[41],stage1_21[61]}
   );
   gpc1163_5 gpc284 (
      {stage0_21[79], stage0_21[80], stage0_21[81]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage0_23[5]},
      {stage0_24[5]},
      {stage1_25[5],stage1_24[18],stage1_23[27],stage1_22[42],stage1_21[62]}
   );
   gpc1163_5 gpc285 (
      {stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage0_23[6]},
      {stage0_24[6]},
      {stage1_25[6],stage1_24[19],stage1_23[28],stage1_22[43],stage1_21[63]}
   );
   gpc1163_5 gpc286 (
      {stage0_21[85], stage0_21[86], stage0_21[87]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage0_23[7]},
      {stage0_24[7]},
      {stage1_25[7],stage1_24[20],stage1_23[29],stage1_22[44],stage1_21[64]}
   );
   gpc1163_5 gpc287 (
      {stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage0_23[8]},
      {stage0_24[8]},
      {stage1_25[8],stage1_24[21],stage1_23[30],stage1_22[45],stage1_21[65]}
   );
   gpc1163_5 gpc288 (
      {stage0_21[91], stage0_21[92], stage0_21[93]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage0_23[9]},
      {stage0_24[9]},
      {stage1_25[9],stage1_24[22],stage1_23[31],stage1_22[46],stage1_21[66]}
   );
   gpc606_5 gpc289 (
      {stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99]},
      {stage0_23[10], stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage1_25[10],stage1_24[23],stage1_23[32],stage1_22[47],stage1_21[67]}
   );
   gpc606_5 gpc290 (
      {stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105]},
      {stage0_23[16], stage0_23[17], stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21]},
      {stage1_25[11],stage1_24[24],stage1_23[33],stage1_22[48],stage1_21[68]}
   );
   gpc606_5 gpc291 (
      {stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111]},
      {stage0_23[22], stage0_23[23], stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27]},
      {stage1_25[12],stage1_24[25],stage1_23[34],stage1_22[49],stage1_21[69]}
   );
   gpc606_5 gpc292 (
      {stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117]},
      {stage0_23[28], stage0_23[29], stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33]},
      {stage1_25[13],stage1_24[26],stage1_23[35],stage1_22[50],stage1_21[70]}
   );
   gpc606_5 gpc293 (
      {stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123]},
      {stage0_23[34], stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage1_25[14],stage1_24[27],stage1_23[36],stage1_22[51],stage1_21[71]}
   );
   gpc606_5 gpc294 (
      {stage0_21[124], stage0_21[125], stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129]},
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45]},
      {stage1_25[15],stage1_24[28],stage1_23[37],stage1_22[52],stage1_21[72]}
   );
   gpc606_5 gpc295 (
      {stage0_21[130], stage0_21[131], stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135]},
      {stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51]},
      {stage1_25[16],stage1_24[29],stage1_23[38],stage1_22[53],stage1_21[73]}
   );
   gpc606_5 gpc296 (
      {stage0_21[136], stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_23[52], stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57]},
      {stage1_25[17],stage1_24[30],stage1_23[39],stage1_22[54],stage1_21[74]}
   );
   gpc606_5 gpc297 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147]},
      {stage0_23[58], stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63]},
      {stage1_25[18],stage1_24[31],stage1_23[40],stage1_22[55],stage1_21[75]}
   );
   gpc606_5 gpc298 (
      {stage0_21[148], stage0_21[149], stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153]},
      {stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69]},
      {stage1_25[19],stage1_24[32],stage1_23[41],stage1_22[56],stage1_21[76]}
   );
   gpc606_5 gpc299 (
      {stage0_21[154], stage0_21[155], stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159]},
      {stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75]},
      {stage1_25[20],stage1_24[33],stage1_23[42],stage1_22[57],stage1_21[77]}
   );
   gpc606_5 gpc300 (
      {stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[21],stage1_24[34],stage1_23[43]}
   );
   gpc606_5 gpc301 (
      {stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[22],stage1_24[35],stage1_23[44]}
   );
   gpc606_5 gpc302 (
      {stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[2],stage1_25[23],stage1_24[36],stage1_23[45]}
   );
   gpc606_5 gpc303 (
      {stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[3],stage1_25[24],stage1_24[37],stage1_23[46]}
   );
   gpc606_5 gpc304 (
      {stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[4],stage1_25[25],stage1_24[38],stage1_23[47]}
   );
   gpc606_5 gpc305 (
      {stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[5],stage1_25[26],stage1_24[39],stage1_23[48]}
   );
   gpc615_5 gpc306 (
      {stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage0_24[10]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[6],stage1_25[27],stage1_24[40],stage1_23[49]}
   );
   gpc615_5 gpc307 (
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121]},
      {stage0_24[11]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[7],stage1_25[28],stage1_24[41],stage1_23[50]}
   );
   gpc606_5 gpc308 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[8],stage1_26[8],stage1_25[29],stage1_24[42]}
   );
   gpc606_5 gpc309 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[9],stage1_26[9],stage1_25[30],stage1_24[43]}
   );
   gpc606_5 gpc310 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[10],stage1_26[10],stage1_25[31],stage1_24[44]}
   );
   gpc606_5 gpc311 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[11],stage1_26[11],stage1_25[32],stage1_24[45]}
   );
   gpc606_5 gpc312 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[12],stage1_26[12],stage1_25[33],stage1_24[46]}
   );
   gpc606_5 gpc313 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[13],stage1_26[13],stage1_25[34],stage1_24[47]}
   );
   gpc606_5 gpc314 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[14],stage1_26[14],stage1_25[35],stage1_24[48]}
   );
   gpc606_5 gpc315 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[15],stage1_26[15],stage1_25[36],stage1_24[49]}
   );
   gpc606_5 gpc316 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[16],stage1_26[16],stage1_25[37],stage1_24[50]}
   );
   gpc606_5 gpc317 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[17],stage1_26[17],stage1_25[38],stage1_24[51]}
   );
   gpc606_5 gpc318 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[18],stage1_26[18],stage1_25[39],stage1_24[52]}
   );
   gpc606_5 gpc319 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[19],stage1_26[19],stage1_25[40],stage1_24[53]}
   );
   gpc606_5 gpc320 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[20],stage1_26[20],stage1_25[41],stage1_24[54]}
   );
   gpc606_5 gpc321 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[21],stage1_26[21],stage1_25[42],stage1_24[55]}
   );
   gpc606_5 gpc322 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[22],stage1_26[22],stage1_25[43],stage1_24[56]}
   );
   gpc606_5 gpc323 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[23],stage1_26[23],stage1_25[44],stage1_24[57]}
   );
   gpc606_5 gpc324 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[24],stage1_26[24],stage1_25[45],stage1_24[58]}
   );
   gpc606_5 gpc325 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[25],stage1_26[25],stage1_25[46],stage1_24[59]}
   );
   gpc606_5 gpc326 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[26],stage1_26[26],stage1_25[47],stage1_24[60]}
   );
   gpc606_5 gpc327 (
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[27],stage1_26[27],stage1_25[48],stage1_24[61]}
   );
   gpc606_5 gpc328 (
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[28],stage1_26[28],stage1_25[49],stage1_24[62]}
   );
   gpc606_5 gpc329 (
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[29],stage1_26[29],stage1_25[50],stage1_24[63]}
   );
   gpc606_5 gpc330 (
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[30],stage1_26[30],stage1_25[51],stage1_24[64]}
   );
   gpc606_5 gpc331 (
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[31],stage1_26[31],stage1_25[52],stage1_24[65]}
   );
   gpc606_5 gpc332 (
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[32],stage1_26[32],stage1_25[53],stage1_24[66]}
   );
   gpc606_5 gpc333 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[25],stage1_27[33],stage1_26[33],stage1_25[54]}
   );
   gpc606_5 gpc334 (
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[26],stage1_27[34],stage1_26[34],stage1_25[55]}
   );
   gpc606_5 gpc335 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[27],stage1_27[35],stage1_26[35],stage1_25[56]}
   );
   gpc606_5 gpc336 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[28],stage1_27[36],stage1_26[36],stage1_25[57]}
   );
   gpc606_5 gpc337 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[29],stage1_27[37],stage1_26[37],stage1_25[58]}
   );
   gpc606_5 gpc338 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[30],stage1_27[38],stage1_26[38],stage1_25[59]}
   );
   gpc606_5 gpc339 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[31],stage1_27[39],stage1_26[39],stage1_25[60]}
   );
   gpc606_5 gpc340 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[32],stage1_27[40],stage1_26[40],stage1_25[61]}
   );
   gpc606_5 gpc341 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[33],stage1_27[41],stage1_26[41],stage1_25[62]}
   );
   gpc606_5 gpc342 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[34],stage1_27[42],stage1_26[42],stage1_25[63]}
   );
   gpc615_5 gpc343 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112]},
      {stage0_26[150]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[35],stage1_27[43],stage1_26[43],stage1_25[64]}
   );
   gpc615_5 gpc344 (
      {stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117]},
      {stage0_26[151]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[36],stage1_27[44],stage1_26[44],stage1_25[65]}
   );
   gpc615_5 gpc345 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122]},
      {stage0_26[152]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[37],stage1_27[45],stage1_26[45],stage1_25[66]}
   );
   gpc615_5 gpc346 (
      {stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_26[153]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[38],stage1_27[46],stage1_26[46],stage1_25[67]}
   );
   gpc615_5 gpc347 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132]},
      {stage0_26[154]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[39],stage1_27[47],stage1_26[47],stage1_25[68]}
   );
   gpc615_5 gpc348 (
      {stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_26[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[40],stage1_27[48],stage1_26[48],stage1_25[69]}
   );
   gpc615_5 gpc349 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142]},
      {stage0_26[156]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[41],stage1_27[49],stage1_26[49],stage1_25[70]}
   );
   gpc615_5 gpc350 (
      {stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_26[157]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[42],stage1_27[50],stage1_26[50],stage1_25[71]}
   );
   gpc615_5 gpc351 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152]},
      {stage0_26[158]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[43],stage1_27[51],stage1_26[51],stage1_25[72]}
   );
   gpc615_5 gpc352 (
      {stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_26[159]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[44],stage1_27[52],stage1_26[52],stage1_25[73]}
   );
   gpc615_5 gpc353 (
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[20],stage1_28[45],stage1_27[53]}
   );
   gpc615_5 gpc354 (
      {stage0_27[125], stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129]},
      {stage0_28[1]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[21],stage1_28[46],stage1_27[54]}
   );
   gpc615_5 gpc355 (
      {stage0_27[130], stage0_27[131], stage0_27[132], stage0_27[133], stage0_27[134]},
      {stage0_28[2]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[22],stage1_28[47],stage1_27[55]}
   );
   gpc615_5 gpc356 (
      {stage0_27[135], stage0_27[136], stage0_27[137], stage0_27[138], stage0_27[139]},
      {stage0_28[3]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[23],stage1_28[48],stage1_27[56]}
   );
   gpc615_5 gpc357 (
      {stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143], stage0_27[144]},
      {stage0_28[4]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[24],stage1_28[49],stage1_27[57]}
   );
   gpc615_5 gpc358 (
      {stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage0_28[5]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[25],stage1_28[50],stage1_27[58]}
   );
   gpc615_5 gpc359 (
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154]},
      {stage0_28[6]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[26],stage1_28[51],stage1_27[59]}
   );
   gpc2135_5 gpc360 (
      {stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_29[42], stage0_29[43], stage0_29[44]},
      {stage0_30[0]},
      {stage0_31[0], stage0_31[1]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[27],stage1_28[52]}
   );
   gpc606_5 gpc361 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[28],stage1_28[53]}
   );
   gpc606_5 gpc362 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[29],stage1_28[54]}
   );
   gpc606_5 gpc363 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[30],stage1_28[55]}
   );
   gpc606_5 gpc364 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[31],stage1_28[56]}
   );
   gpc606_5 gpc365 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[32],stage1_28[57]}
   );
   gpc606_5 gpc366 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[33],stage1_28[58]}
   );
   gpc606_5 gpc367 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[34],stage1_28[59]}
   );
   gpc606_5 gpc368 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[35],stage1_28[60]}
   );
   gpc606_5 gpc369 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[36],stage1_28[61]}
   );
   gpc606_5 gpc370 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[37],stage1_28[62]}
   );
   gpc606_5 gpc371 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[38],stage1_28[63]}
   );
   gpc606_5 gpc372 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[39],stage1_28[64]}
   );
   gpc606_5 gpc373 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[40],stage1_28[65]}
   );
   gpc606_5 gpc374 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[41],stage1_28[66]}
   );
   gpc606_5 gpc375 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89], stage0_30[90]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[42],stage1_28[67]}
   );
   gpc606_5 gpc376 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95], stage0_30[96]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[43],stage1_28[68]}
   );
   gpc606_5 gpc377 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101], stage0_30[102]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[44],stage1_28[69]}
   );
   gpc606_5 gpc378 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107], stage0_30[108]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[45],stage1_28[70]}
   );
   gpc606_5 gpc379 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113], stage0_30[114]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[46],stage1_28[71]}
   );
   gpc606_5 gpc380 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119], stage0_30[120]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[47],stage1_28[72]}
   );
   gpc606_5 gpc381 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125], stage0_30[126]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[48],stage1_28[73]}
   );
   gpc606_5 gpc382 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131], stage0_30[132]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[49],stage1_28[74]}
   );
   gpc606_5 gpc383 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137], stage0_30[138]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[50],stage1_28[75]}
   );
   gpc606_5 gpc384 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143], stage0_30[144]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[51],stage1_28[76]}
   );
   gpc606_5 gpc385 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149], stage0_30[150]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[52],stage1_28[77]}
   );
   gpc606_5 gpc386 (
      {stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49], stage0_29[50]},
      {stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage1_33[0],stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[53]}
   );
   gpc606_5 gpc387 (
      {stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55], stage0_29[56]},
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage1_33[1],stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[54]}
   );
   gpc606_5 gpc388 (
      {stage0_29[57], stage0_29[58], stage0_29[59], stage0_29[60], stage0_29[61], stage0_29[62]},
      {stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18], stage0_31[19]},
      {stage1_33[2],stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[55]}
   );
   gpc606_5 gpc389 (
      {stage0_29[63], stage0_29[64], stage0_29[65], stage0_29[66], stage0_29[67], stage0_29[68]},
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24], stage0_31[25]},
      {stage1_33[3],stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[56]}
   );
   gpc606_5 gpc390 (
      {stage0_29[69], stage0_29[70], stage0_29[71], stage0_29[72], stage0_29[73], stage0_29[74]},
      {stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30], stage0_31[31]},
      {stage1_33[4],stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[57]}
   );
   gpc606_5 gpc391 (
      {stage0_29[75], stage0_29[76], stage0_29[77], stage0_29[78], stage0_29[79], stage0_29[80]},
      {stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36], stage0_31[37]},
      {stage1_33[5],stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[58]}
   );
   gpc606_5 gpc392 (
      {stage0_29[81], stage0_29[82], stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86]},
      {stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42], stage0_31[43]},
      {stage1_33[6],stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[59]}
   );
   gpc606_5 gpc393 (
      {stage0_29[87], stage0_29[88], stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92]},
      {stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48], stage0_31[49]},
      {stage1_33[7],stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[60]}
   );
   gpc606_5 gpc394 (
      {stage0_29[93], stage0_29[94], stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98]},
      {stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54], stage0_31[55]},
      {stage1_33[8],stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[61]}
   );
   gpc606_5 gpc395 (
      {stage0_29[99], stage0_29[100], stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104]},
      {stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60], stage0_31[61]},
      {stage1_33[9],stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[62]}
   );
   gpc606_5 gpc396 (
      {stage0_29[105], stage0_29[106], stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110]},
      {stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67]},
      {stage1_33[10],stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[63]}
   );
   gpc606_5 gpc397 (
      {stage0_29[111], stage0_29[112], stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116]},
      {stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage1_33[11],stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[64]}
   );
   gpc606_5 gpc398 (
      {stage0_29[117], stage0_29[118], stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122]},
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78], stage0_31[79]},
      {stage1_33[12],stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[65]}
   );
   gpc606_5 gpc399 (
      {stage0_29[123], stage0_29[124], stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128]},
      {stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83], stage0_31[84], stage0_31[85]},
      {stage1_33[13],stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[66]}
   );
   gpc606_5 gpc400 (
      {stage0_29[129], stage0_29[130], stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134]},
      {stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89], stage0_31[90], stage0_31[91]},
      {stage1_33[14],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[67]}
   );
   gpc606_5 gpc401 (
      {stage0_29[135], stage0_29[136], stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140]},
      {stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97]},
      {stage1_33[15],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[68]}
   );
   gpc606_5 gpc402 (
      {stage0_29[141], stage0_29[142], stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146]},
      {stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage1_33[16],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[69]}
   );
   gpc606_5 gpc403 (
      {stage0_29[147], stage0_29[148], stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152]},
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108], stage0_31[109]},
      {stage1_33[17],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[70]}
   );
   gpc606_5 gpc404 (
      {stage0_29[153], stage0_29[154], stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158]},
      {stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113], stage0_31[114], stage0_31[115]},
      {stage1_33[18],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[71]}
   );
   gpc1_1 gpc405 (
      {stage0_0[144]},
      {stage1_0[32]}
   );
   gpc1_1 gpc406 (
      {stage0_0[145]},
      {stage1_0[33]}
   );
   gpc1_1 gpc407 (
      {stage0_0[146]},
      {stage1_0[34]}
   );
   gpc1_1 gpc408 (
      {stage0_0[147]},
      {stage1_0[35]}
   );
   gpc1_1 gpc409 (
      {stage0_0[148]},
      {stage1_0[36]}
   );
   gpc1_1 gpc410 (
      {stage0_0[149]},
      {stage1_0[37]}
   );
   gpc1_1 gpc411 (
      {stage0_0[150]},
      {stage1_0[38]}
   );
   gpc1_1 gpc412 (
      {stage0_0[151]},
      {stage1_0[39]}
   );
   gpc1_1 gpc413 (
      {stage0_0[152]},
      {stage1_0[40]}
   );
   gpc1_1 gpc414 (
      {stage0_0[153]},
      {stage1_0[41]}
   );
   gpc1_1 gpc415 (
      {stage0_0[154]},
      {stage1_0[42]}
   );
   gpc1_1 gpc416 (
      {stage0_0[155]},
      {stage1_0[43]}
   );
   gpc1_1 gpc417 (
      {stage0_0[156]},
      {stage1_0[44]}
   );
   gpc1_1 gpc418 (
      {stage0_0[157]},
      {stage1_0[45]}
   );
   gpc1_1 gpc419 (
      {stage0_0[158]},
      {stage1_0[46]}
   );
   gpc1_1 gpc420 (
      {stage0_0[159]},
      {stage1_0[47]}
   );
   gpc1_1 gpc421 (
      {stage0_0[160]},
      {stage1_0[48]}
   );
   gpc1_1 gpc422 (
      {stage0_0[161]},
      {stage1_0[49]}
   );
   gpc1_1 gpc423 (
      {stage0_1[144]},
      {stage1_1[38]}
   );
   gpc1_1 gpc424 (
      {stage0_1[145]},
      {stage1_1[39]}
   );
   gpc1_1 gpc425 (
      {stage0_1[146]},
      {stage1_1[40]}
   );
   gpc1_1 gpc426 (
      {stage0_1[147]},
      {stage1_1[41]}
   );
   gpc1_1 gpc427 (
      {stage0_1[148]},
      {stage1_1[42]}
   );
   gpc1_1 gpc428 (
      {stage0_1[149]},
      {stage1_1[43]}
   );
   gpc1_1 gpc429 (
      {stage0_1[150]},
      {stage1_1[44]}
   );
   gpc1_1 gpc430 (
      {stage0_1[151]},
      {stage1_1[45]}
   );
   gpc1_1 gpc431 (
      {stage0_1[152]},
      {stage1_1[46]}
   );
   gpc1_1 gpc432 (
      {stage0_1[153]},
      {stage1_1[47]}
   );
   gpc1_1 gpc433 (
      {stage0_1[154]},
      {stage1_1[48]}
   );
   gpc1_1 gpc434 (
      {stage0_1[155]},
      {stage1_1[49]}
   );
   gpc1_1 gpc435 (
      {stage0_1[156]},
      {stage1_1[50]}
   );
   gpc1_1 gpc436 (
      {stage0_1[157]},
      {stage1_1[51]}
   );
   gpc1_1 gpc437 (
      {stage0_1[158]},
      {stage1_1[52]}
   );
   gpc1_1 gpc438 (
      {stage0_1[159]},
      {stage1_1[53]}
   );
   gpc1_1 gpc439 (
      {stage0_1[160]},
      {stage1_1[54]}
   );
   gpc1_1 gpc440 (
      {stage0_1[161]},
      {stage1_1[55]}
   );
   gpc1_1 gpc441 (
      {stage0_3[155]},
      {stage1_3[69]}
   );
   gpc1_1 gpc442 (
      {stage0_3[156]},
      {stage1_3[70]}
   );
   gpc1_1 gpc443 (
      {stage0_3[157]},
      {stage1_3[71]}
   );
   gpc1_1 gpc444 (
      {stage0_3[158]},
      {stage1_3[72]}
   );
   gpc1_1 gpc445 (
      {stage0_3[159]},
      {stage1_3[73]}
   );
   gpc1_1 gpc446 (
      {stage0_3[160]},
      {stage1_3[74]}
   );
   gpc1_1 gpc447 (
      {stage0_3[161]},
      {stage1_3[75]}
   );
   gpc1_1 gpc448 (
      {stage0_4[139]},
      {stage1_4[72]}
   );
   gpc1_1 gpc449 (
      {stage0_4[140]},
      {stage1_4[73]}
   );
   gpc1_1 gpc450 (
      {stage0_4[141]},
      {stage1_4[74]}
   );
   gpc1_1 gpc451 (
      {stage0_4[142]},
      {stage1_4[75]}
   );
   gpc1_1 gpc452 (
      {stage0_4[143]},
      {stage1_4[76]}
   );
   gpc1_1 gpc453 (
      {stage0_4[144]},
      {stage1_4[77]}
   );
   gpc1_1 gpc454 (
      {stage0_4[145]},
      {stage1_4[78]}
   );
   gpc1_1 gpc455 (
      {stage0_4[146]},
      {stage1_4[79]}
   );
   gpc1_1 gpc456 (
      {stage0_4[147]},
      {stage1_4[80]}
   );
   gpc1_1 gpc457 (
      {stage0_4[148]},
      {stage1_4[81]}
   );
   gpc1_1 gpc458 (
      {stage0_4[149]},
      {stage1_4[82]}
   );
   gpc1_1 gpc459 (
      {stage0_4[150]},
      {stage1_4[83]}
   );
   gpc1_1 gpc460 (
      {stage0_4[151]},
      {stage1_4[84]}
   );
   gpc1_1 gpc461 (
      {stage0_4[152]},
      {stage1_4[85]}
   );
   gpc1_1 gpc462 (
      {stage0_4[153]},
      {stage1_4[86]}
   );
   gpc1_1 gpc463 (
      {stage0_4[154]},
      {stage1_4[87]}
   );
   gpc1_1 gpc464 (
      {stage0_4[155]},
      {stage1_4[88]}
   );
   gpc1_1 gpc465 (
      {stage0_4[156]},
      {stage1_4[89]}
   );
   gpc1_1 gpc466 (
      {stage0_4[157]},
      {stage1_4[90]}
   );
   gpc1_1 gpc467 (
      {stage0_4[158]},
      {stage1_4[91]}
   );
   gpc1_1 gpc468 (
      {stage0_4[159]},
      {stage1_4[92]}
   );
   gpc1_1 gpc469 (
      {stage0_4[160]},
      {stage1_4[93]}
   );
   gpc1_1 gpc470 (
      {stage0_4[161]},
      {stage1_4[94]}
   );
   gpc1_1 gpc471 (
      {stage0_6[124]},
      {stage1_6[68]}
   );
   gpc1_1 gpc472 (
      {stage0_6[125]},
      {stage1_6[69]}
   );
   gpc1_1 gpc473 (
      {stage0_6[126]},
      {stage1_6[70]}
   );
   gpc1_1 gpc474 (
      {stage0_6[127]},
      {stage1_6[71]}
   );
   gpc1_1 gpc475 (
      {stage0_6[128]},
      {stage1_6[72]}
   );
   gpc1_1 gpc476 (
      {stage0_6[129]},
      {stage1_6[73]}
   );
   gpc1_1 gpc477 (
      {stage0_6[130]},
      {stage1_6[74]}
   );
   gpc1_1 gpc478 (
      {stage0_6[131]},
      {stage1_6[75]}
   );
   gpc1_1 gpc479 (
      {stage0_6[132]},
      {stage1_6[76]}
   );
   gpc1_1 gpc480 (
      {stage0_6[133]},
      {stage1_6[77]}
   );
   gpc1_1 gpc481 (
      {stage0_6[134]},
      {stage1_6[78]}
   );
   gpc1_1 gpc482 (
      {stage0_6[135]},
      {stage1_6[79]}
   );
   gpc1_1 gpc483 (
      {stage0_6[136]},
      {stage1_6[80]}
   );
   gpc1_1 gpc484 (
      {stage0_6[137]},
      {stage1_6[81]}
   );
   gpc1_1 gpc485 (
      {stage0_6[138]},
      {stage1_6[82]}
   );
   gpc1_1 gpc486 (
      {stage0_6[139]},
      {stage1_6[83]}
   );
   gpc1_1 gpc487 (
      {stage0_6[140]},
      {stage1_6[84]}
   );
   gpc1_1 gpc488 (
      {stage0_6[141]},
      {stage1_6[85]}
   );
   gpc1_1 gpc489 (
      {stage0_6[142]},
      {stage1_6[86]}
   );
   gpc1_1 gpc490 (
      {stage0_6[143]},
      {stage1_6[87]}
   );
   gpc1_1 gpc491 (
      {stage0_6[144]},
      {stage1_6[88]}
   );
   gpc1_1 gpc492 (
      {stage0_6[145]},
      {stage1_6[89]}
   );
   gpc1_1 gpc493 (
      {stage0_6[146]},
      {stage1_6[90]}
   );
   gpc1_1 gpc494 (
      {stage0_6[147]},
      {stage1_6[91]}
   );
   gpc1_1 gpc495 (
      {stage0_6[148]},
      {stage1_6[92]}
   );
   gpc1_1 gpc496 (
      {stage0_6[149]},
      {stage1_6[93]}
   );
   gpc1_1 gpc497 (
      {stage0_6[150]},
      {stage1_6[94]}
   );
   gpc1_1 gpc498 (
      {stage0_6[151]},
      {stage1_6[95]}
   );
   gpc1_1 gpc499 (
      {stage0_6[152]},
      {stage1_6[96]}
   );
   gpc1_1 gpc500 (
      {stage0_6[153]},
      {stage1_6[97]}
   );
   gpc1_1 gpc501 (
      {stage0_6[154]},
      {stage1_6[98]}
   );
   gpc1_1 gpc502 (
      {stage0_6[155]},
      {stage1_6[99]}
   );
   gpc1_1 gpc503 (
      {stage0_6[156]},
      {stage1_6[100]}
   );
   gpc1_1 gpc504 (
      {stage0_6[157]},
      {stage1_6[101]}
   );
   gpc1_1 gpc505 (
      {stage0_6[158]},
      {stage1_6[102]}
   );
   gpc1_1 gpc506 (
      {stage0_6[159]},
      {stage1_6[103]}
   );
   gpc1_1 gpc507 (
      {stage0_6[160]},
      {stage1_6[104]}
   );
   gpc1_1 gpc508 (
      {stage0_6[161]},
      {stage1_6[105]}
   );
   gpc1_1 gpc509 (
      {stage0_7[158]},
      {stage1_7[62]}
   );
   gpc1_1 gpc510 (
      {stage0_7[159]},
      {stage1_7[63]}
   );
   gpc1_1 gpc511 (
      {stage0_7[160]},
      {stage1_7[64]}
   );
   gpc1_1 gpc512 (
      {stage0_7[161]},
      {stage1_7[65]}
   );
   gpc1_1 gpc513 (
      {stage0_9[152]},
      {stage1_9[67]}
   );
   gpc1_1 gpc514 (
      {stage0_9[153]},
      {stage1_9[68]}
   );
   gpc1_1 gpc515 (
      {stage0_9[154]},
      {stage1_9[69]}
   );
   gpc1_1 gpc516 (
      {stage0_9[155]},
      {stage1_9[70]}
   );
   gpc1_1 gpc517 (
      {stage0_9[156]},
      {stage1_9[71]}
   );
   gpc1_1 gpc518 (
      {stage0_9[157]},
      {stage1_9[72]}
   );
   gpc1_1 gpc519 (
      {stage0_9[158]},
      {stage1_9[73]}
   );
   gpc1_1 gpc520 (
      {stage0_9[159]},
      {stage1_9[74]}
   );
   gpc1_1 gpc521 (
      {stage0_9[160]},
      {stage1_9[75]}
   );
   gpc1_1 gpc522 (
      {stage0_9[161]},
      {stage1_9[76]}
   );
   gpc1_1 gpc523 (
      {stage0_10[141]},
      {stage1_10[72]}
   );
   gpc1_1 gpc524 (
      {stage0_10[142]},
      {stage1_10[73]}
   );
   gpc1_1 gpc525 (
      {stage0_10[143]},
      {stage1_10[74]}
   );
   gpc1_1 gpc526 (
      {stage0_10[144]},
      {stage1_10[75]}
   );
   gpc1_1 gpc527 (
      {stage0_10[145]},
      {stage1_10[76]}
   );
   gpc1_1 gpc528 (
      {stage0_10[146]},
      {stage1_10[77]}
   );
   gpc1_1 gpc529 (
      {stage0_10[147]},
      {stage1_10[78]}
   );
   gpc1_1 gpc530 (
      {stage0_10[148]},
      {stage1_10[79]}
   );
   gpc1_1 gpc531 (
      {stage0_10[149]},
      {stage1_10[80]}
   );
   gpc1_1 gpc532 (
      {stage0_10[150]},
      {stage1_10[81]}
   );
   gpc1_1 gpc533 (
      {stage0_10[151]},
      {stage1_10[82]}
   );
   gpc1_1 gpc534 (
      {stage0_10[152]},
      {stage1_10[83]}
   );
   gpc1_1 gpc535 (
      {stage0_10[153]},
      {stage1_10[84]}
   );
   gpc1_1 gpc536 (
      {stage0_10[154]},
      {stage1_10[85]}
   );
   gpc1_1 gpc537 (
      {stage0_10[155]},
      {stage1_10[86]}
   );
   gpc1_1 gpc538 (
      {stage0_10[156]},
      {stage1_10[87]}
   );
   gpc1_1 gpc539 (
      {stage0_10[157]},
      {stage1_10[88]}
   );
   gpc1_1 gpc540 (
      {stage0_10[158]},
      {stage1_10[89]}
   );
   gpc1_1 gpc541 (
      {stage0_10[159]},
      {stage1_10[90]}
   );
   gpc1_1 gpc542 (
      {stage0_10[160]},
      {stage1_10[91]}
   );
   gpc1_1 gpc543 (
      {stage0_10[161]},
      {stage1_10[92]}
   );
   gpc1_1 gpc544 (
      {stage0_11[155]},
      {stage1_11[60]}
   );
   gpc1_1 gpc545 (
      {stage0_11[156]},
      {stage1_11[61]}
   );
   gpc1_1 gpc546 (
      {stage0_11[157]},
      {stage1_11[62]}
   );
   gpc1_1 gpc547 (
      {stage0_11[158]},
      {stage1_11[63]}
   );
   gpc1_1 gpc548 (
      {stage0_11[159]},
      {stage1_11[64]}
   );
   gpc1_1 gpc549 (
      {stage0_11[160]},
      {stage1_11[65]}
   );
   gpc1_1 gpc550 (
      {stage0_11[161]},
      {stage1_11[66]}
   );
   gpc1_1 gpc551 (
      {stage0_13[144]},
      {stage1_13[68]}
   );
   gpc1_1 gpc552 (
      {stage0_13[145]},
      {stage1_13[69]}
   );
   gpc1_1 gpc553 (
      {stage0_13[146]},
      {stage1_13[70]}
   );
   gpc1_1 gpc554 (
      {stage0_13[147]},
      {stage1_13[71]}
   );
   gpc1_1 gpc555 (
      {stage0_13[148]},
      {stage1_13[72]}
   );
   gpc1_1 gpc556 (
      {stage0_13[149]},
      {stage1_13[73]}
   );
   gpc1_1 gpc557 (
      {stage0_13[150]},
      {stage1_13[74]}
   );
   gpc1_1 gpc558 (
      {stage0_13[151]},
      {stage1_13[75]}
   );
   gpc1_1 gpc559 (
      {stage0_13[152]},
      {stage1_13[76]}
   );
   gpc1_1 gpc560 (
      {stage0_13[153]},
      {stage1_13[77]}
   );
   gpc1_1 gpc561 (
      {stage0_13[154]},
      {stage1_13[78]}
   );
   gpc1_1 gpc562 (
      {stage0_13[155]},
      {stage1_13[79]}
   );
   gpc1_1 gpc563 (
      {stage0_13[156]},
      {stage1_13[80]}
   );
   gpc1_1 gpc564 (
      {stage0_13[157]},
      {stage1_13[81]}
   );
   gpc1_1 gpc565 (
      {stage0_13[158]},
      {stage1_13[82]}
   );
   gpc1_1 gpc566 (
      {stage0_13[159]},
      {stage1_13[83]}
   );
   gpc1_1 gpc567 (
      {stage0_13[160]},
      {stage1_13[84]}
   );
   gpc1_1 gpc568 (
      {stage0_13[161]},
      {stage1_13[85]}
   );
   gpc1_1 gpc569 (
      {stage0_14[161]},
      {stage1_14[68]}
   );
   gpc1_1 gpc570 (
      {stage0_16[111]},
      {stage1_16[56]}
   );
   gpc1_1 gpc571 (
      {stage0_16[112]},
      {stage1_16[57]}
   );
   gpc1_1 gpc572 (
      {stage0_16[113]},
      {stage1_16[58]}
   );
   gpc1_1 gpc573 (
      {stage0_16[114]},
      {stage1_16[59]}
   );
   gpc1_1 gpc574 (
      {stage0_16[115]},
      {stage1_16[60]}
   );
   gpc1_1 gpc575 (
      {stage0_16[116]},
      {stage1_16[61]}
   );
   gpc1_1 gpc576 (
      {stage0_16[117]},
      {stage1_16[62]}
   );
   gpc1_1 gpc577 (
      {stage0_16[118]},
      {stage1_16[63]}
   );
   gpc1_1 gpc578 (
      {stage0_16[119]},
      {stage1_16[64]}
   );
   gpc1_1 gpc579 (
      {stage0_16[120]},
      {stage1_16[65]}
   );
   gpc1_1 gpc580 (
      {stage0_16[121]},
      {stage1_16[66]}
   );
   gpc1_1 gpc581 (
      {stage0_16[122]},
      {stage1_16[67]}
   );
   gpc1_1 gpc582 (
      {stage0_16[123]},
      {stage1_16[68]}
   );
   gpc1_1 gpc583 (
      {stage0_16[124]},
      {stage1_16[69]}
   );
   gpc1_1 gpc584 (
      {stage0_16[125]},
      {stage1_16[70]}
   );
   gpc1_1 gpc585 (
      {stage0_16[126]},
      {stage1_16[71]}
   );
   gpc1_1 gpc586 (
      {stage0_16[127]},
      {stage1_16[72]}
   );
   gpc1_1 gpc587 (
      {stage0_16[128]},
      {stage1_16[73]}
   );
   gpc1_1 gpc588 (
      {stage0_16[129]},
      {stage1_16[74]}
   );
   gpc1_1 gpc589 (
      {stage0_16[130]},
      {stage1_16[75]}
   );
   gpc1_1 gpc590 (
      {stage0_16[131]},
      {stage1_16[76]}
   );
   gpc1_1 gpc591 (
      {stage0_16[132]},
      {stage1_16[77]}
   );
   gpc1_1 gpc592 (
      {stage0_16[133]},
      {stage1_16[78]}
   );
   gpc1_1 gpc593 (
      {stage0_16[134]},
      {stage1_16[79]}
   );
   gpc1_1 gpc594 (
      {stage0_16[135]},
      {stage1_16[80]}
   );
   gpc1_1 gpc595 (
      {stage0_16[136]},
      {stage1_16[81]}
   );
   gpc1_1 gpc596 (
      {stage0_16[137]},
      {stage1_16[82]}
   );
   gpc1_1 gpc597 (
      {stage0_16[138]},
      {stage1_16[83]}
   );
   gpc1_1 gpc598 (
      {stage0_16[139]},
      {stage1_16[84]}
   );
   gpc1_1 gpc599 (
      {stage0_16[140]},
      {stage1_16[85]}
   );
   gpc1_1 gpc600 (
      {stage0_16[141]},
      {stage1_16[86]}
   );
   gpc1_1 gpc601 (
      {stage0_16[142]},
      {stage1_16[87]}
   );
   gpc1_1 gpc602 (
      {stage0_16[143]},
      {stage1_16[88]}
   );
   gpc1_1 gpc603 (
      {stage0_16[144]},
      {stage1_16[89]}
   );
   gpc1_1 gpc604 (
      {stage0_16[145]},
      {stage1_16[90]}
   );
   gpc1_1 gpc605 (
      {stage0_16[146]},
      {stage1_16[91]}
   );
   gpc1_1 gpc606 (
      {stage0_16[147]},
      {stage1_16[92]}
   );
   gpc1_1 gpc607 (
      {stage0_16[148]},
      {stage1_16[93]}
   );
   gpc1_1 gpc608 (
      {stage0_16[149]},
      {stage1_16[94]}
   );
   gpc1_1 gpc609 (
      {stage0_16[150]},
      {stage1_16[95]}
   );
   gpc1_1 gpc610 (
      {stage0_16[151]},
      {stage1_16[96]}
   );
   gpc1_1 gpc611 (
      {stage0_16[152]},
      {stage1_16[97]}
   );
   gpc1_1 gpc612 (
      {stage0_16[153]},
      {stage1_16[98]}
   );
   gpc1_1 gpc613 (
      {stage0_16[154]},
      {stage1_16[99]}
   );
   gpc1_1 gpc614 (
      {stage0_16[155]},
      {stage1_16[100]}
   );
   gpc1_1 gpc615 (
      {stage0_16[156]},
      {stage1_16[101]}
   );
   gpc1_1 gpc616 (
      {stage0_16[157]},
      {stage1_16[102]}
   );
   gpc1_1 gpc617 (
      {stage0_16[158]},
      {stage1_16[103]}
   );
   gpc1_1 gpc618 (
      {stage0_16[159]},
      {stage1_16[104]}
   );
   gpc1_1 gpc619 (
      {stage0_16[160]},
      {stage1_16[105]}
   );
   gpc1_1 gpc620 (
      {stage0_16[161]},
      {stage1_16[106]}
   );
   gpc1_1 gpc621 (
      {stage0_18[142]},
      {stage1_18[62]}
   );
   gpc1_1 gpc622 (
      {stage0_18[143]},
      {stage1_18[63]}
   );
   gpc1_1 gpc623 (
      {stage0_18[144]},
      {stage1_18[64]}
   );
   gpc1_1 gpc624 (
      {stage0_18[145]},
      {stage1_18[65]}
   );
   gpc1_1 gpc625 (
      {stage0_18[146]},
      {stage1_18[66]}
   );
   gpc1_1 gpc626 (
      {stage0_18[147]},
      {stage1_18[67]}
   );
   gpc1_1 gpc627 (
      {stage0_18[148]},
      {stage1_18[68]}
   );
   gpc1_1 gpc628 (
      {stage0_18[149]},
      {stage1_18[69]}
   );
   gpc1_1 gpc629 (
      {stage0_18[150]},
      {stage1_18[70]}
   );
   gpc1_1 gpc630 (
      {stage0_18[151]},
      {stage1_18[71]}
   );
   gpc1_1 gpc631 (
      {stage0_18[152]},
      {stage1_18[72]}
   );
   gpc1_1 gpc632 (
      {stage0_18[153]},
      {stage1_18[73]}
   );
   gpc1_1 gpc633 (
      {stage0_18[154]},
      {stage1_18[74]}
   );
   gpc1_1 gpc634 (
      {stage0_18[155]},
      {stage1_18[75]}
   );
   gpc1_1 gpc635 (
      {stage0_18[156]},
      {stage1_18[76]}
   );
   gpc1_1 gpc636 (
      {stage0_18[157]},
      {stage1_18[77]}
   );
   gpc1_1 gpc637 (
      {stage0_18[158]},
      {stage1_18[78]}
   );
   gpc1_1 gpc638 (
      {stage0_18[159]},
      {stage1_18[79]}
   );
   gpc1_1 gpc639 (
      {stage0_18[160]},
      {stage1_18[80]}
   );
   gpc1_1 gpc640 (
      {stage0_18[161]},
      {stage1_18[81]}
   );
   gpc1_1 gpc641 (
      {stage0_19[154]},
      {stage1_19[59]}
   );
   gpc1_1 gpc642 (
      {stage0_19[155]},
      {stage1_19[60]}
   );
   gpc1_1 gpc643 (
      {stage0_19[156]},
      {stage1_19[61]}
   );
   gpc1_1 gpc644 (
      {stage0_19[157]},
      {stage1_19[62]}
   );
   gpc1_1 gpc645 (
      {stage0_19[158]},
      {stage1_19[63]}
   );
   gpc1_1 gpc646 (
      {stage0_19[159]},
      {stage1_19[64]}
   );
   gpc1_1 gpc647 (
      {stage0_19[160]},
      {stage1_19[65]}
   );
   gpc1_1 gpc648 (
      {stage0_19[161]},
      {stage1_19[66]}
   );
   gpc1_1 gpc649 (
      {stage0_21[160]},
      {stage1_21[78]}
   );
   gpc1_1 gpc650 (
      {stage0_21[161]},
      {stage1_21[79]}
   );
   gpc1_1 gpc651 (
      {stage0_22[138]},
      {stage1_22[58]}
   );
   gpc1_1 gpc652 (
      {stage0_22[139]},
      {stage1_22[59]}
   );
   gpc1_1 gpc653 (
      {stage0_22[140]},
      {stage1_22[60]}
   );
   gpc1_1 gpc654 (
      {stage0_22[141]},
      {stage1_22[61]}
   );
   gpc1_1 gpc655 (
      {stage0_22[142]},
      {stage1_22[62]}
   );
   gpc1_1 gpc656 (
      {stage0_22[143]},
      {stage1_22[63]}
   );
   gpc1_1 gpc657 (
      {stage0_22[144]},
      {stage1_22[64]}
   );
   gpc1_1 gpc658 (
      {stage0_22[145]},
      {stage1_22[65]}
   );
   gpc1_1 gpc659 (
      {stage0_22[146]},
      {stage1_22[66]}
   );
   gpc1_1 gpc660 (
      {stage0_22[147]},
      {stage1_22[67]}
   );
   gpc1_1 gpc661 (
      {stage0_22[148]},
      {stage1_22[68]}
   );
   gpc1_1 gpc662 (
      {stage0_22[149]},
      {stage1_22[69]}
   );
   gpc1_1 gpc663 (
      {stage0_22[150]},
      {stage1_22[70]}
   );
   gpc1_1 gpc664 (
      {stage0_22[151]},
      {stage1_22[71]}
   );
   gpc1_1 gpc665 (
      {stage0_22[152]},
      {stage1_22[72]}
   );
   gpc1_1 gpc666 (
      {stage0_22[153]},
      {stage1_22[73]}
   );
   gpc1_1 gpc667 (
      {stage0_22[154]},
      {stage1_22[74]}
   );
   gpc1_1 gpc668 (
      {stage0_22[155]},
      {stage1_22[75]}
   );
   gpc1_1 gpc669 (
      {stage0_22[156]},
      {stage1_22[76]}
   );
   gpc1_1 gpc670 (
      {stage0_22[157]},
      {stage1_22[77]}
   );
   gpc1_1 gpc671 (
      {stage0_22[158]},
      {stage1_22[78]}
   );
   gpc1_1 gpc672 (
      {stage0_22[159]},
      {stage1_22[79]}
   );
   gpc1_1 gpc673 (
      {stage0_22[160]},
      {stage1_22[80]}
   );
   gpc1_1 gpc674 (
      {stage0_22[161]},
      {stage1_22[81]}
   );
   gpc1_1 gpc675 (
      {stage0_23[122]},
      {stage1_23[51]}
   );
   gpc1_1 gpc676 (
      {stage0_23[123]},
      {stage1_23[52]}
   );
   gpc1_1 gpc677 (
      {stage0_23[124]},
      {stage1_23[53]}
   );
   gpc1_1 gpc678 (
      {stage0_23[125]},
      {stage1_23[54]}
   );
   gpc1_1 gpc679 (
      {stage0_23[126]},
      {stage1_23[55]}
   );
   gpc1_1 gpc680 (
      {stage0_23[127]},
      {stage1_23[56]}
   );
   gpc1_1 gpc681 (
      {stage0_23[128]},
      {stage1_23[57]}
   );
   gpc1_1 gpc682 (
      {stage0_23[129]},
      {stage1_23[58]}
   );
   gpc1_1 gpc683 (
      {stage0_23[130]},
      {stage1_23[59]}
   );
   gpc1_1 gpc684 (
      {stage0_23[131]},
      {stage1_23[60]}
   );
   gpc1_1 gpc685 (
      {stage0_23[132]},
      {stage1_23[61]}
   );
   gpc1_1 gpc686 (
      {stage0_23[133]},
      {stage1_23[62]}
   );
   gpc1_1 gpc687 (
      {stage0_23[134]},
      {stage1_23[63]}
   );
   gpc1_1 gpc688 (
      {stage0_23[135]},
      {stage1_23[64]}
   );
   gpc1_1 gpc689 (
      {stage0_23[136]},
      {stage1_23[65]}
   );
   gpc1_1 gpc690 (
      {stage0_23[137]},
      {stage1_23[66]}
   );
   gpc1_1 gpc691 (
      {stage0_23[138]},
      {stage1_23[67]}
   );
   gpc1_1 gpc692 (
      {stage0_23[139]},
      {stage1_23[68]}
   );
   gpc1_1 gpc693 (
      {stage0_23[140]},
      {stage1_23[69]}
   );
   gpc1_1 gpc694 (
      {stage0_23[141]},
      {stage1_23[70]}
   );
   gpc1_1 gpc695 (
      {stage0_23[142]},
      {stage1_23[71]}
   );
   gpc1_1 gpc696 (
      {stage0_23[143]},
      {stage1_23[72]}
   );
   gpc1_1 gpc697 (
      {stage0_23[144]},
      {stage1_23[73]}
   );
   gpc1_1 gpc698 (
      {stage0_23[145]},
      {stage1_23[74]}
   );
   gpc1_1 gpc699 (
      {stage0_23[146]},
      {stage1_23[75]}
   );
   gpc1_1 gpc700 (
      {stage0_23[147]},
      {stage1_23[76]}
   );
   gpc1_1 gpc701 (
      {stage0_23[148]},
      {stage1_23[77]}
   );
   gpc1_1 gpc702 (
      {stage0_23[149]},
      {stage1_23[78]}
   );
   gpc1_1 gpc703 (
      {stage0_23[150]},
      {stage1_23[79]}
   );
   gpc1_1 gpc704 (
      {stage0_23[151]},
      {stage1_23[80]}
   );
   gpc1_1 gpc705 (
      {stage0_23[152]},
      {stage1_23[81]}
   );
   gpc1_1 gpc706 (
      {stage0_23[153]},
      {stage1_23[82]}
   );
   gpc1_1 gpc707 (
      {stage0_23[154]},
      {stage1_23[83]}
   );
   gpc1_1 gpc708 (
      {stage0_23[155]},
      {stage1_23[84]}
   );
   gpc1_1 gpc709 (
      {stage0_23[156]},
      {stage1_23[85]}
   );
   gpc1_1 gpc710 (
      {stage0_23[157]},
      {stage1_23[86]}
   );
   gpc1_1 gpc711 (
      {stage0_23[158]},
      {stage1_23[87]}
   );
   gpc1_1 gpc712 (
      {stage0_23[159]},
      {stage1_23[88]}
   );
   gpc1_1 gpc713 (
      {stage0_23[160]},
      {stage1_23[89]}
   );
   gpc1_1 gpc714 (
      {stage0_23[161]},
      {stage1_23[90]}
   );
   gpc1_1 gpc715 (
      {stage0_25[158]},
      {stage1_25[74]}
   );
   gpc1_1 gpc716 (
      {stage0_25[159]},
      {stage1_25[75]}
   );
   gpc1_1 gpc717 (
      {stage0_25[160]},
      {stage1_25[76]}
   );
   gpc1_1 gpc718 (
      {stage0_25[161]},
      {stage1_25[77]}
   );
   gpc1_1 gpc719 (
      {stage0_26[160]},
      {stage1_26[53]}
   );
   gpc1_1 gpc720 (
      {stage0_26[161]},
      {stage1_26[54]}
   );
   gpc1_1 gpc721 (
      {stage0_27[155]},
      {stage1_27[60]}
   );
   gpc1_1 gpc722 (
      {stage0_27[156]},
      {stage1_27[61]}
   );
   gpc1_1 gpc723 (
      {stage0_27[157]},
      {stage1_27[62]}
   );
   gpc1_1 gpc724 (
      {stage0_27[158]},
      {stage1_27[63]}
   );
   gpc1_1 gpc725 (
      {stage0_27[159]},
      {stage1_27[64]}
   );
   gpc1_1 gpc726 (
      {stage0_27[160]},
      {stage1_27[65]}
   );
   gpc1_1 gpc727 (
      {stage0_27[161]},
      {stage1_27[66]}
   );
   gpc1_1 gpc728 (
      {stage0_29[159]},
      {stage1_29[72]}
   );
   gpc1_1 gpc729 (
      {stage0_29[160]},
      {stage1_29[73]}
   );
   gpc1_1 gpc730 (
      {stage0_29[161]},
      {stage1_29[74]}
   );
   gpc1_1 gpc731 (
      {stage0_30[151]},
      {stage1_30[52]}
   );
   gpc1_1 gpc732 (
      {stage0_30[152]},
      {stage1_30[53]}
   );
   gpc1_1 gpc733 (
      {stage0_30[153]},
      {stage1_30[54]}
   );
   gpc1_1 gpc734 (
      {stage0_30[154]},
      {stage1_30[55]}
   );
   gpc1_1 gpc735 (
      {stage0_30[155]},
      {stage1_30[56]}
   );
   gpc1_1 gpc736 (
      {stage0_30[156]},
      {stage1_30[57]}
   );
   gpc1_1 gpc737 (
      {stage0_30[157]},
      {stage1_30[58]}
   );
   gpc1_1 gpc738 (
      {stage0_30[158]},
      {stage1_30[59]}
   );
   gpc1_1 gpc739 (
      {stage0_30[159]},
      {stage1_30[60]}
   );
   gpc1_1 gpc740 (
      {stage0_30[160]},
      {stage1_30[61]}
   );
   gpc1_1 gpc741 (
      {stage0_30[161]},
      {stage1_30[62]}
   );
   gpc1_1 gpc742 (
      {stage0_31[116]},
      {stage1_31[52]}
   );
   gpc1_1 gpc743 (
      {stage0_31[117]},
      {stage1_31[53]}
   );
   gpc1_1 gpc744 (
      {stage0_31[118]},
      {stage1_31[54]}
   );
   gpc1_1 gpc745 (
      {stage0_31[119]},
      {stage1_31[55]}
   );
   gpc1_1 gpc746 (
      {stage0_31[120]},
      {stage1_31[56]}
   );
   gpc1_1 gpc747 (
      {stage0_31[121]},
      {stage1_31[57]}
   );
   gpc1_1 gpc748 (
      {stage0_31[122]},
      {stage1_31[58]}
   );
   gpc1_1 gpc749 (
      {stage0_31[123]},
      {stage1_31[59]}
   );
   gpc1_1 gpc750 (
      {stage0_31[124]},
      {stage1_31[60]}
   );
   gpc1_1 gpc751 (
      {stage0_31[125]},
      {stage1_31[61]}
   );
   gpc1_1 gpc752 (
      {stage0_31[126]},
      {stage1_31[62]}
   );
   gpc1_1 gpc753 (
      {stage0_31[127]},
      {stage1_31[63]}
   );
   gpc1_1 gpc754 (
      {stage0_31[128]},
      {stage1_31[64]}
   );
   gpc1_1 gpc755 (
      {stage0_31[129]},
      {stage1_31[65]}
   );
   gpc1_1 gpc756 (
      {stage0_31[130]},
      {stage1_31[66]}
   );
   gpc1_1 gpc757 (
      {stage0_31[131]},
      {stage1_31[67]}
   );
   gpc1_1 gpc758 (
      {stage0_31[132]},
      {stage1_31[68]}
   );
   gpc1_1 gpc759 (
      {stage0_31[133]},
      {stage1_31[69]}
   );
   gpc1_1 gpc760 (
      {stage0_31[134]},
      {stage1_31[70]}
   );
   gpc1_1 gpc761 (
      {stage0_31[135]},
      {stage1_31[71]}
   );
   gpc1_1 gpc762 (
      {stage0_31[136]},
      {stage1_31[72]}
   );
   gpc1_1 gpc763 (
      {stage0_31[137]},
      {stage1_31[73]}
   );
   gpc1_1 gpc764 (
      {stage0_31[138]},
      {stage1_31[74]}
   );
   gpc1_1 gpc765 (
      {stage0_31[139]},
      {stage1_31[75]}
   );
   gpc1_1 gpc766 (
      {stage0_31[140]},
      {stage1_31[76]}
   );
   gpc1_1 gpc767 (
      {stage0_31[141]},
      {stage1_31[77]}
   );
   gpc1_1 gpc768 (
      {stage0_31[142]},
      {stage1_31[78]}
   );
   gpc1_1 gpc769 (
      {stage0_31[143]},
      {stage1_31[79]}
   );
   gpc1_1 gpc770 (
      {stage0_31[144]},
      {stage1_31[80]}
   );
   gpc1_1 gpc771 (
      {stage0_31[145]},
      {stage1_31[81]}
   );
   gpc1_1 gpc772 (
      {stage0_31[146]},
      {stage1_31[82]}
   );
   gpc1_1 gpc773 (
      {stage0_31[147]},
      {stage1_31[83]}
   );
   gpc1_1 gpc774 (
      {stage0_31[148]},
      {stage1_31[84]}
   );
   gpc1_1 gpc775 (
      {stage0_31[149]},
      {stage1_31[85]}
   );
   gpc1_1 gpc776 (
      {stage0_31[150]},
      {stage1_31[86]}
   );
   gpc1_1 gpc777 (
      {stage0_31[151]},
      {stage1_31[87]}
   );
   gpc1_1 gpc778 (
      {stage0_31[152]},
      {stage1_31[88]}
   );
   gpc1_1 gpc779 (
      {stage0_31[153]},
      {stage1_31[89]}
   );
   gpc1_1 gpc780 (
      {stage0_31[154]},
      {stage1_31[90]}
   );
   gpc1_1 gpc781 (
      {stage0_31[155]},
      {stage1_31[91]}
   );
   gpc1_1 gpc782 (
      {stage0_31[156]},
      {stage1_31[92]}
   );
   gpc1_1 gpc783 (
      {stage0_31[157]},
      {stage1_31[93]}
   );
   gpc1_1 gpc784 (
      {stage0_31[158]},
      {stage1_31[94]}
   );
   gpc1_1 gpc785 (
      {stage0_31[159]},
      {stage1_31[95]}
   );
   gpc1_1 gpc786 (
      {stage0_31[160]},
      {stage1_31[96]}
   );
   gpc1_1 gpc787 (
      {stage0_31[161]},
      {stage1_31[97]}
   );
   gpc1163_5 gpc788 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc789 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc790 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc791 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc792 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[18]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc793 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[19]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc794 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[20]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc795 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[21]},
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc796 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[22]},
      {stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc797 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[23]},
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc798 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[24]},
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc799 (
      {stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc800 (
      {stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc801 (
      {stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc802 (
      {stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48]},
      {stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc803 (
      {stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54]},
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage2_5[4],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc615_5 gpc804 (
      {stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_3[33]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[5],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc805 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[6]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc806 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[7]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc807 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[8]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc808 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[9],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc809 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[10]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[10],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc810 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[11]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[6],stage2_5[11],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc811 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[6],stage2_6[7],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc812 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[7],stage2_6[8],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc813 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[8],stage2_6[9],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc814 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[9],stage2_6[10],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc815 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[10],stage2_6[11],stage2_5[16],stage2_4[27]}
   );
   gpc606_5 gpc816 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[11],stage2_6[12],stage2_5[17],stage2_4[28]}
   );
   gpc606_5 gpc817 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[12],stage2_6[13],stage2_5[18],stage2_4[29]}
   );
   gpc606_5 gpc818 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[13],stage2_6[14],stage2_5[19],stage2_4[30]}
   );
   gpc606_5 gpc819 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[14],stage2_6[15],stage2_5[20],stage2_4[31]}
   );
   gpc606_5 gpc820 (
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[15],stage2_6[16],stage2_5[21],stage2_4[32]}
   );
   gpc606_5 gpc821 (
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[16],stage2_6[17],stage2_5[22],stage2_4[33]}
   );
   gpc606_5 gpc822 (
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[17],stage2_6[18],stage2_5[23],stage2_4[34]}
   );
   gpc606_5 gpc823 (
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[18],stage2_6[19],stage2_5[24],stage2_4[35]}
   );
   gpc606_5 gpc824 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[13],stage2_7[19],stage2_6[20],stage2_5[25]}
   );
   gpc606_5 gpc825 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[14],stage2_7[20],stage2_6[21],stage2_5[26]}
   );
   gpc606_5 gpc826 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[15],stage2_7[21],stage2_6[22],stage2_5[27]}
   );
   gpc606_5 gpc827 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[16],stage2_7[22],stage2_6[23]}
   );
   gpc606_5 gpc828 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[17],stage2_7[23],stage2_6[24]}
   );
   gpc606_5 gpc829 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[18],stage2_7[24],stage2_6[25]}
   );
   gpc606_5 gpc830 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[19],stage2_7[25],stage2_6[26]}
   );
   gpc606_5 gpc831 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[20],stage2_7[26]}
   );
   gpc606_5 gpc832 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[5],stage2_9[8],stage2_8[21],stage2_7[27]}
   );
   gpc606_5 gpc833 (
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[6],stage2_9[9],stage2_8[22],stage2_7[28]}
   );
   gpc606_5 gpc834 (
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[7],stage2_9[10],stage2_8[23],stage2_7[29]}
   );
   gpc606_5 gpc835 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[8],stage2_9[11],stage2_8[24],stage2_7[30]}
   );
   gpc606_5 gpc836 (
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[9],stage2_9[12],stage2_8[25],stage2_7[31]}
   );
   gpc606_5 gpc837 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[10],stage2_9[13],stage2_8[26],stage2_7[32]}
   );
   gpc606_5 gpc838 (
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[11],stage2_9[14],stage2_8[27],stage2_7[33]}
   );
   gpc606_5 gpc839 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[8],stage2_10[12],stage2_9[15],stage2_8[28]}
   );
   gpc606_5 gpc840 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[9],stage2_10[13],stage2_9[16],stage2_8[29]}
   );
   gpc606_5 gpc841 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[10],stage2_10[14],stage2_9[17],stage2_8[30]}
   );
   gpc606_5 gpc842 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[11],stage2_10[15],stage2_9[18],stage2_8[31]}
   );
   gpc606_5 gpc843 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[12],stage2_10[16],stage2_9[19],stage2_8[32]}
   );
   gpc606_5 gpc844 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[13],stage2_10[17],stage2_9[20]}
   );
   gpc615_5 gpc845 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58]},
      {stage1_10[30]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[14],stage2_10[18],stage2_9[21]}
   );
   gpc615_5 gpc846 (
      {stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63]},
      {stage1_10[31]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[15],stage2_10[19],stage2_9[22]}
   );
   gpc615_5 gpc847 (
      {stage1_9[64], stage1_9[65], stage1_9[66], stage1_9[67], stage1_9[68]},
      {stage1_10[32]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[16],stage2_10[20],stage2_9[23]}
   );
   gpc606_5 gpc848 (
      {stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37], stage1_10[38]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[17],stage2_10[21]}
   );
   gpc606_5 gpc849 (
      {stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[18],stage2_10[22]}
   );
   gpc606_5 gpc850 (
      {stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[19],stage2_10[23]}
   );
   gpc606_5 gpc851 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[20],stage2_10[24]}
   );
   gpc606_5 gpc852 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[21],stage2_10[25]}
   );
   gpc606_5 gpc853 (
      {stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[22],stage2_10[26]}
   );
   gpc606_5 gpc854 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73], stage1_10[74]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[23],stage2_10[27]}
   );
   gpc606_5 gpc855 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[24]}
   );
   gpc606_5 gpc856 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[25]}
   );
   gpc606_5 gpc857 (
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[26]}
   );
   gpc606_5 gpc858 (
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[27]}
   );
   gpc615_5 gpc859 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[42]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[28]}
   );
   gpc615_5 gpc860 (
      {stage1_11[53], stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57]},
      {stage1_12[43]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[29]}
   );
   gpc606_5 gpc861 (
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[13],stage2_13[17],stage2_12[22]}
   );
   gpc606_5 gpc862 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54], stage1_12[55]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[14],stage2_13[18],stage2_12[23]}
   );
   gpc1415_5 gpc863 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40]},
      {stage1_14[12]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3]},
      {stage1_16[0]},
      {stage2_17[0],stage2_16[2],stage2_15[8],stage2_14[15],stage2_13[19]}
   );
   gpc615_5 gpc864 (
      {stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45]},
      {stage1_14[13]},
      {stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage2_17[1],stage2_16[3],stage2_15[9],stage2_14[16],stage2_13[20]}
   );
   gpc615_5 gpc865 (
      {stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage1_14[14]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15]},
      {stage2_17[2],stage2_16[4],stage2_15[10],stage2_14[17],stage2_13[21]}
   );
   gpc615_5 gpc866 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55]},
      {stage1_14[15]},
      {stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21]},
      {stage2_17[3],stage2_16[5],stage2_15[11],stage2_14[18],stage2_13[22]}
   );
   gpc615_5 gpc867 (
      {stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60]},
      {stage1_14[16]},
      {stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage2_17[4],stage2_16[6],stage2_15[12],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc868 (
      {stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_14[17]},
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage2_17[5],stage2_16[7],stage2_15[13],stage2_14[20],stage2_13[24]}
   );
   gpc606_5 gpc869 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[0],stage2_17[6],stage2_16[8],stage2_15[14],stage2_14[21]}
   );
   gpc606_5 gpc870 (
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[1],stage2_17[7],stage2_16[9],stage2_15[15],stage2_14[22]}
   );
   gpc606_5 gpc871 (
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage2_18[2],stage2_17[8],stage2_16[10],stage2_15[16],stage2_14[23]}
   );
   gpc606_5 gpc872 (
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage2_18[3],stage2_17[9],stage2_16[11],stage2_15[17],stage2_14[24]}
   );
   gpc606_5 gpc873 (
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30]},
      {stage2_18[4],stage2_17[10],stage2_16[12],stage2_15[18],stage2_14[25]}
   );
   gpc606_5 gpc874 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36]},
      {stage2_18[5],stage2_17[11],stage2_16[13],stage2_15[19],stage2_14[26]}
   );
   gpc606_5 gpc875 (
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42]},
      {stage2_18[6],stage2_17[12],stage2_16[14],stage2_15[20],stage2_14[27]}
   );
   gpc1406_5 gpc876 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[15],stage2_15[21]}
   );
   gpc615_5 gpc877 (
      {stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43], stage1_15[44]},
      {stage1_16[43]},
      {stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[16],stage2_15[22]}
   );
   gpc615_5 gpc878 (
      {stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_16[44]},
      {stage1_17[10], stage1_17[11], stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[17],stage2_15[23]}
   );
   gpc615_5 gpc879 (
      {stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_17[16]},
      {stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6]},
      {stage2_20[0],stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[18]}
   );
   gpc615_5 gpc880 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54]},
      {stage1_17[17]},
      {stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12]},
      {stage2_20[1],stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[19]}
   );
   gpc615_5 gpc881 (
      {stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_17[18]},
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18]},
      {stage2_20[2],stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[20]}
   );
   gpc615_5 gpc882 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_17[19]},
      {stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24]},
      {stage2_20[3],stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[21]}
   );
   gpc615_5 gpc883 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69]},
      {stage1_17[20]},
      {stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30]},
      {stage2_20[4],stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[22]}
   );
   gpc615_5 gpc884 (
      {stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74]},
      {stage1_17[21]},
      {stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage2_20[5],stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[23]}
   );
   gpc615_5 gpc885 (
      {stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_17[22]},
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42]},
      {stage2_20[6],stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[24]}
   );
   gpc615_5 gpc886 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84]},
      {stage1_17[23]},
      {stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48]},
      {stage2_20[7],stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[25]}
   );
   gpc615_5 gpc887 (
      {stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_17[24]},
      {stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54]},
      {stage2_20[8],stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[26]}
   );
   gpc606_5 gpc888 (
      {stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[9],stage2_19[12],stage2_18[19],stage2_17[25]}
   );
   gpc606_5 gpc889 (
      {stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[10],stage2_19[13],stage2_18[20],stage2_17[26]}
   );
   gpc606_5 gpc890 (
      {stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41], stage1_17[42]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[11],stage2_19[14],stage2_18[21],stage2_17[27]}
   );
   gpc615_5 gpc891 (
      {stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_18[55]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[12],stage2_19[15],stage2_18[22],stage2_17[28]}
   );
   gpc615_5 gpc892 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52]},
      {stage1_18[56]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[13],stage2_19[16],stage2_18[23],stage2_17[29]}
   );
   gpc615_5 gpc893 (
      {stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage1_18[57]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[14],stage2_19[17],stage2_18[24],stage2_17[30]}
   );
   gpc606_5 gpc894 (
      {stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[15],stage2_19[18],stage2_18[25]}
   );
   gpc606_5 gpc895 (
      {stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[16],stage2_19[19],stage2_18[26]}
   );
   gpc606_5 gpc896 (
      {stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[8],stage2_20[17],stage2_19[20],stage2_18[27]}
   );
   gpc606_5 gpc897 (
      {stage1_18[76], stage1_18[77], stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[9],stage2_20[18],stage2_19[21],stage2_18[28]}
   );
   gpc606_5 gpc898 (
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[10],stage2_20[19],stage2_19[22]}
   );
   gpc606_5 gpc899 (
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[11],stage2_20[20],stage2_19[23]}
   );
   gpc606_5 gpc900 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[12],stage2_20[21],stage2_19[24]}
   );
   gpc606_5 gpc901 (
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[13],stage2_20[22],stage2_19[25]}
   );
   gpc606_5 gpc902 (
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[14],stage2_20[23],stage2_19[26]}
   );
   gpc606_5 gpc903 (
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[9],stage2_21[15],stage2_20[24]}
   );
   gpc606_5 gpc904 (
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[10],stage2_21[16],stage2_20[25]}
   );
   gpc606_5 gpc905 (
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[11],stage2_21[17],stage2_20[26]}
   );
   gpc615_5 gpc906 (
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46]},
      {stage1_21[30]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[8],stage2_22[12],stage2_21[18],stage2_20[27]}
   );
   gpc615_5 gpc907 (
      {stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_21[31]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[9],stage2_22[13],stage2_21[19],stage2_20[28]}
   );
   gpc606_5 gpc908 (
      {stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[5],stage2_23[10],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc909 (
      {stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[6],stage2_23[11],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc910 (
      {stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[7],stage2_23[12],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc911 (
      {stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[8],stage2_23[13],stage2_22[17],stage2_21[23]}
   );
   gpc606_5 gpc912 (
      {stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[9],stage2_23[14],stage2_22[18],stage2_21[24]}
   );
   gpc606_5 gpc913 (
      {stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[10],stage2_23[15],stage2_22[19],stage2_21[25]}
   );
   gpc606_5 gpc914 (
      {stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[11],stage2_23[16],stage2_22[20],stage2_21[26]}
   );
   gpc606_5 gpc915 (
      {stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[12],stage2_23[17],stage2_22[21],stage2_21[27]}
   );
   gpc606_5 gpc916 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[8],stage2_24[13],stage2_23[18],stage2_22[22]}
   );
   gpc606_5 gpc917 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[9],stage2_24[14],stage2_23[19],stage2_22[23]}
   );
   gpc606_5 gpc918 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[10],stage2_24[15],stage2_23[20],stage2_22[24]}
   );
   gpc606_5 gpc919 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[11],stage2_24[16],stage2_23[21],stage2_22[25]}
   );
   gpc606_5 gpc920 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[12],stage2_24[17],stage2_23[22],stage2_22[26]}
   );
   gpc606_5 gpc921 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[13],stage2_24[18],stage2_23[23],stage2_22[27]}
   );
   gpc606_5 gpc922 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[14],stage2_24[19],stage2_23[24],stage2_22[28]}
   );
   gpc606_5 gpc923 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[15],stage2_24[20],stage2_23[25],stage2_22[29]}
   );
   gpc606_5 gpc924 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[16],stage2_24[21],stage2_23[26]}
   );
   gpc606_5 gpc925 (
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[17],stage2_24[22],stage2_23[27]}
   );
   gpc606_5 gpc926 (
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[18],stage2_24[23],stage2_23[28]}
   );
   gpc606_5 gpc927 (
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[19],stage2_24[24],stage2_23[29]}
   );
   gpc606_5 gpc928 (
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[20],stage2_24[25],stage2_23[30]}
   );
   gpc606_5 gpc929 (
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[13],stage2_25[21],stage2_24[26]}
   );
   gpc606_5 gpc930 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[14],stage2_25[22],stage2_24[27]}
   );
   gpc606_5 gpc931 (
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[15],stage2_25[23]}
   );
   gpc606_5 gpc932 (
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[16],stage2_25[24]}
   );
   gpc606_5 gpc933 (
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[17],stage2_25[25]}
   );
   gpc606_5 gpc934 (
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[18],stage2_25[26]}
   );
   gpc606_5 gpc935 (
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[6],stage2_27[11],stage2_26[19],stage2_25[27]}
   );
   gpc606_5 gpc936 (
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[7],stage2_27[12],stage2_26[20],stage2_25[28]}
   );
   gpc606_5 gpc937 (
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[8],stage2_27[13],stage2_26[21],stage2_25[29]}
   );
   gpc606_5 gpc938 (
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[9],stage2_27[14],stage2_26[22],stage2_25[30]}
   );
   gpc606_5 gpc939 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[8],stage2_28[10],stage2_27[15],stage2_26[23]}
   );
   gpc606_5 gpc940 (
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[9],stage2_28[11],stage2_27[16],stage2_26[24]}
   );
   gpc606_5 gpc941 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[10],stage2_28[12],stage2_27[17],stage2_26[25]}
   );
   gpc606_5 gpc942 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[11],stage2_28[13],stage2_27[18],stage2_26[26]}
   );
   gpc606_5 gpc943 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[12],stage2_28[14],stage2_27[19],stage2_26[27]}
   );
   gpc606_5 gpc944 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[13],stage2_28[15],stage2_27[20],stage2_26[28]}
   );
   gpc606_5 gpc945 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[14],stage2_28[16],stage2_27[21],stage2_26[29]}
   );
   gpc615_5 gpc946 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[15],stage2_28[17],stage2_27[22]}
   );
   gpc615_5 gpc947 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[16],stage2_28[18],stage2_27[23]}
   );
   gpc606_5 gpc948 (
      {stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[2],stage2_30[9],stage2_29[17],stage2_28[19]}
   );
   gpc606_5 gpc949 (
      {stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[3],stage2_30[10],stage2_29[18],stage2_28[20]}
   );
   gpc606_5 gpc950 (
      {stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[4],stage2_30[11],stage2_29[19],stage2_28[21]}
   );
   gpc615_5 gpc951 (
      {stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66]},
      {stage1_29[12]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[5],stage2_30[12],stage2_29[20],stage2_28[22]}
   );
   gpc615_5 gpc952 (
      {stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_29[13]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[6],stage2_30[13],stage2_29[21],stage2_28[23]}
   );
   gpc606_5 gpc953 (
      {stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[5],stage2_31[7],stage2_30[14],stage2_29[22]}
   );
   gpc606_5 gpc954 (
      {stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[6],stage2_31[8],stage2_30[15],stage2_29[23]}
   );
   gpc606_5 gpc955 (
      {stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[7],stage2_31[9],stage2_30[16],stage2_29[24]}
   );
   gpc606_5 gpc956 (
      {stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[8],stage2_31[10],stage2_30[17],stage2_29[25]}
   );
   gpc606_5 gpc957 (
      {stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[9],stage2_31[11],stage2_30[18],stage2_29[26]}
   );
   gpc606_5 gpc958 (
      {stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[10],stage2_31[12],stage2_30[19],stage2_29[27]}
   );
   gpc615_5 gpc959 (
      {stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53], stage1_29[54]},
      {stage1_30[30]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[11],stage2_31[13],stage2_30[20],stage2_29[28]}
   );
   gpc615_5 gpc960 (
      {stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_30[31]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[12],stage2_31[14],stage2_30[21],stage2_29[29]}
   );
   gpc615_5 gpc961 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64]},
      {stage1_30[32]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[13],stage2_31[15],stage2_30[22],stage2_29[30]}
   );
   gpc615_5 gpc962 (
      {stage1_29[65], stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69]},
      {stage1_30[33]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[14],stage2_31[16],stage2_30[23],stage2_29[31]}
   );
   gpc615_5 gpc963 (
      {stage1_29[70], stage1_29[71], stage1_29[72], stage1_29[73], stage1_29[74]},
      {stage1_30[34]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[15],stage2_31[17],stage2_30[24],stage2_29[32]}
   );
   gpc615_5 gpc964 (
      {stage1_30[35], stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39]},
      {stage1_31[66]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[11],stage2_32[16],stage2_31[18],stage2_30[25]}
   );
   gpc615_5 gpc965 (
      {stage1_30[40], stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44]},
      {stage1_31[67]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[12],stage2_32[17],stage2_31[19],stage2_30[26]}
   );
   gpc615_5 gpc966 (
      {stage1_30[45], stage1_30[46], stage1_30[47], stage1_30[48], stage1_30[49]},
      {stage1_31[68]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[13],stage2_32[18],stage2_31[20],stage2_30[27]}
   );
   gpc615_5 gpc967 (
      {stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_31[69]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[14],stage2_32[19],stage2_31[21],stage2_30[28]}
   );
   gpc135_4 gpc968 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[24], stage1_32[25], stage1_32[26]},
      {stage1_33[0]},
      {stage2_34[4],stage2_33[15],stage2_32[20],stage2_31[22]}
   );
   gpc606_5 gpc969 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[0],stage2_34[5],stage2_33[16],stage2_32[21],stage2_31[23]}
   );
   gpc606_5 gpc970 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[1],stage2_34[6],stage2_33[17],stage2_32[22],stage2_31[24]}
   );
   gpc1_1 gpc971 (
      {stage1_1[55]},
      {stage2_1[16]}
   );
   gpc1_1 gpc972 (
      {stage1_3[64]},
      {stage2_3[23]}
   );
   gpc1_1 gpc973 (
      {stage1_3[65]},
      {stage2_3[24]}
   );
   gpc1_1 gpc974 (
      {stage1_3[66]},
      {stage2_3[25]}
   );
   gpc1_1 gpc975 (
      {stage1_3[67]},
      {stage2_3[26]}
   );
   gpc1_1 gpc976 (
      {stage1_3[68]},
      {stage2_3[27]}
   );
   gpc1_1 gpc977 (
      {stage1_3[69]},
      {stage2_3[28]}
   );
   gpc1_1 gpc978 (
      {stage1_3[70]},
      {stage2_3[29]}
   );
   gpc1_1 gpc979 (
      {stage1_3[71]},
      {stage2_3[30]}
   );
   gpc1_1 gpc980 (
      {stage1_3[72]},
      {stage2_3[31]}
   );
   gpc1_1 gpc981 (
      {stage1_3[73]},
      {stage2_3[32]}
   );
   gpc1_1 gpc982 (
      {stage1_3[74]},
      {stage2_3[33]}
   );
   gpc1_1 gpc983 (
      {stage1_3[75]},
      {stage2_3[34]}
   );
   gpc1_1 gpc984 (
      {stage1_4[90]},
      {stage2_4[36]}
   );
   gpc1_1 gpc985 (
      {stage1_4[91]},
      {stage2_4[37]}
   );
   gpc1_1 gpc986 (
      {stage1_4[92]},
      {stage2_4[38]}
   );
   gpc1_1 gpc987 (
      {stage1_4[93]},
      {stage2_4[39]}
   );
   gpc1_1 gpc988 (
      {stage1_4[94]},
      {stage2_4[40]}
   );
   gpc1_1 gpc989 (
      {stage1_6[102]},
      {stage2_6[27]}
   );
   gpc1_1 gpc990 (
      {stage1_6[103]},
      {stage2_6[28]}
   );
   gpc1_1 gpc991 (
      {stage1_6[104]},
      {stage2_6[29]}
   );
   gpc1_1 gpc992 (
      {stage1_6[105]},
      {stage2_6[30]}
   );
   gpc1_1 gpc993 (
      {stage1_9[69]},
      {stage2_9[24]}
   );
   gpc1_1 gpc994 (
      {stage1_9[70]},
      {stage2_9[25]}
   );
   gpc1_1 gpc995 (
      {stage1_9[71]},
      {stage2_9[26]}
   );
   gpc1_1 gpc996 (
      {stage1_9[72]},
      {stage2_9[27]}
   );
   gpc1_1 gpc997 (
      {stage1_9[73]},
      {stage2_9[28]}
   );
   gpc1_1 gpc998 (
      {stage1_9[74]},
      {stage2_9[29]}
   );
   gpc1_1 gpc999 (
      {stage1_9[75]},
      {stage2_9[30]}
   );
   gpc1_1 gpc1000 (
      {stage1_9[76]},
      {stage2_9[31]}
   );
   gpc1_1 gpc1001 (
      {stage1_10[75]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1002 (
      {stage1_10[76]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1003 (
      {stage1_10[77]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1004 (
      {stage1_10[78]},
      {stage2_10[31]}
   );
   gpc1_1 gpc1005 (
      {stage1_10[79]},
      {stage2_10[32]}
   );
   gpc1_1 gpc1006 (
      {stage1_10[80]},
      {stage2_10[33]}
   );
   gpc1_1 gpc1007 (
      {stage1_10[81]},
      {stage2_10[34]}
   );
   gpc1_1 gpc1008 (
      {stage1_10[82]},
      {stage2_10[35]}
   );
   gpc1_1 gpc1009 (
      {stage1_10[83]},
      {stage2_10[36]}
   );
   gpc1_1 gpc1010 (
      {stage1_10[84]},
      {stage2_10[37]}
   );
   gpc1_1 gpc1011 (
      {stage1_10[85]},
      {stage2_10[38]}
   );
   gpc1_1 gpc1012 (
      {stage1_10[86]},
      {stage2_10[39]}
   );
   gpc1_1 gpc1013 (
      {stage1_10[87]},
      {stage2_10[40]}
   );
   gpc1_1 gpc1014 (
      {stage1_10[88]},
      {stage2_10[41]}
   );
   gpc1_1 gpc1015 (
      {stage1_10[89]},
      {stage2_10[42]}
   );
   gpc1_1 gpc1016 (
      {stage1_10[90]},
      {stage2_10[43]}
   );
   gpc1_1 gpc1017 (
      {stage1_10[91]},
      {stage2_10[44]}
   );
   gpc1_1 gpc1018 (
      {stage1_10[92]},
      {stage2_10[45]}
   );
   gpc1_1 gpc1019 (
      {stage1_11[58]},
      {stage2_11[30]}
   );
   gpc1_1 gpc1020 (
      {stage1_11[59]},
      {stage2_11[31]}
   );
   gpc1_1 gpc1021 (
      {stage1_11[60]},
      {stage2_11[32]}
   );
   gpc1_1 gpc1022 (
      {stage1_11[61]},
      {stage2_11[33]}
   );
   gpc1_1 gpc1023 (
      {stage1_11[62]},
      {stage2_11[34]}
   );
   gpc1_1 gpc1024 (
      {stage1_11[63]},
      {stage2_11[35]}
   );
   gpc1_1 gpc1025 (
      {stage1_11[64]},
      {stage2_11[36]}
   );
   gpc1_1 gpc1026 (
      {stage1_11[65]},
      {stage2_11[37]}
   );
   gpc1_1 gpc1027 (
      {stage1_11[66]},
      {stage2_11[38]}
   );
   gpc1_1 gpc1028 (
      {stage1_13[66]},
      {stage2_13[25]}
   );
   gpc1_1 gpc1029 (
      {stage1_13[67]},
      {stage2_13[26]}
   );
   gpc1_1 gpc1030 (
      {stage1_13[68]},
      {stage2_13[27]}
   );
   gpc1_1 gpc1031 (
      {stage1_13[69]},
      {stage2_13[28]}
   );
   gpc1_1 gpc1032 (
      {stage1_13[70]},
      {stage2_13[29]}
   );
   gpc1_1 gpc1033 (
      {stage1_13[71]},
      {stage2_13[30]}
   );
   gpc1_1 gpc1034 (
      {stage1_13[72]},
      {stage2_13[31]}
   );
   gpc1_1 gpc1035 (
      {stage1_13[73]},
      {stage2_13[32]}
   );
   gpc1_1 gpc1036 (
      {stage1_13[74]},
      {stage2_13[33]}
   );
   gpc1_1 gpc1037 (
      {stage1_13[75]},
      {stage2_13[34]}
   );
   gpc1_1 gpc1038 (
      {stage1_13[76]},
      {stage2_13[35]}
   );
   gpc1_1 gpc1039 (
      {stage1_13[77]},
      {stage2_13[36]}
   );
   gpc1_1 gpc1040 (
      {stage1_13[78]},
      {stage2_13[37]}
   );
   gpc1_1 gpc1041 (
      {stage1_13[79]},
      {stage2_13[38]}
   );
   gpc1_1 gpc1042 (
      {stage1_13[80]},
      {stage2_13[39]}
   );
   gpc1_1 gpc1043 (
      {stage1_13[81]},
      {stage2_13[40]}
   );
   gpc1_1 gpc1044 (
      {stage1_13[82]},
      {stage2_13[41]}
   );
   gpc1_1 gpc1045 (
      {stage1_13[83]},
      {stage2_13[42]}
   );
   gpc1_1 gpc1046 (
      {stage1_13[84]},
      {stage2_13[43]}
   );
   gpc1_1 gpc1047 (
      {stage1_13[85]},
      {stage2_13[44]}
   );
   gpc1_1 gpc1048 (
      {stage1_14[60]},
      {stage2_14[28]}
   );
   gpc1_1 gpc1049 (
      {stage1_14[61]},
      {stage2_14[29]}
   );
   gpc1_1 gpc1050 (
      {stage1_14[62]},
      {stage2_14[30]}
   );
   gpc1_1 gpc1051 (
      {stage1_14[63]},
      {stage2_14[31]}
   );
   gpc1_1 gpc1052 (
      {stage1_14[64]},
      {stage2_14[32]}
   );
   gpc1_1 gpc1053 (
      {stage1_14[65]},
      {stage2_14[33]}
   );
   gpc1_1 gpc1054 (
      {stage1_14[66]},
      {stage2_14[34]}
   );
   gpc1_1 gpc1055 (
      {stage1_14[67]},
      {stage2_14[35]}
   );
   gpc1_1 gpc1056 (
      {stage1_14[68]},
      {stage2_14[36]}
   );
   gpc1_1 gpc1057 (
      {stage1_15[50]},
      {stage2_15[24]}
   );
   gpc1_1 gpc1058 (
      {stage1_15[51]},
      {stage2_15[25]}
   );
   gpc1_1 gpc1059 (
      {stage1_15[52]},
      {stage2_15[26]}
   );
   gpc1_1 gpc1060 (
      {stage1_15[53]},
      {stage2_15[27]}
   );
   gpc1_1 gpc1061 (
      {stage1_15[54]},
      {stage2_15[28]}
   );
   gpc1_1 gpc1062 (
      {stage1_15[55]},
      {stage2_15[29]}
   );
   gpc1_1 gpc1063 (
      {stage1_15[56]},
      {stage2_15[30]}
   );
   gpc1_1 gpc1064 (
      {stage1_15[57]},
      {stage2_15[31]}
   );
   gpc1_1 gpc1065 (
      {stage1_15[58]},
      {stage2_15[32]}
   );
   gpc1_1 gpc1066 (
      {stage1_15[59]},
      {stage2_15[33]}
   );
   gpc1_1 gpc1067 (
      {stage1_16[90]},
      {stage2_16[27]}
   );
   gpc1_1 gpc1068 (
      {stage1_16[91]},
      {stage2_16[28]}
   );
   gpc1_1 gpc1069 (
      {stage1_16[92]},
      {stage2_16[29]}
   );
   gpc1_1 gpc1070 (
      {stage1_16[93]},
      {stage2_16[30]}
   );
   gpc1_1 gpc1071 (
      {stage1_16[94]},
      {stage2_16[31]}
   );
   gpc1_1 gpc1072 (
      {stage1_16[95]},
      {stage2_16[32]}
   );
   gpc1_1 gpc1073 (
      {stage1_16[96]},
      {stage2_16[33]}
   );
   gpc1_1 gpc1074 (
      {stage1_16[97]},
      {stage2_16[34]}
   );
   gpc1_1 gpc1075 (
      {stage1_16[98]},
      {stage2_16[35]}
   );
   gpc1_1 gpc1076 (
      {stage1_16[99]},
      {stage2_16[36]}
   );
   gpc1_1 gpc1077 (
      {stage1_16[100]},
      {stage2_16[37]}
   );
   gpc1_1 gpc1078 (
      {stage1_16[101]},
      {stage2_16[38]}
   );
   gpc1_1 gpc1079 (
      {stage1_16[102]},
      {stage2_16[39]}
   );
   gpc1_1 gpc1080 (
      {stage1_16[103]},
      {stage2_16[40]}
   );
   gpc1_1 gpc1081 (
      {stage1_16[104]},
      {stage2_16[41]}
   );
   gpc1_1 gpc1082 (
      {stage1_16[105]},
      {stage2_16[42]}
   );
   gpc1_1 gpc1083 (
      {stage1_16[106]},
      {stage2_16[43]}
   );
   gpc1_1 gpc1084 (
      {stage1_17[58]},
      {stage2_17[31]}
   );
   gpc1_1 gpc1085 (
      {stage1_17[59]},
      {stage2_17[32]}
   );
   gpc1_1 gpc1086 (
      {stage1_17[60]},
      {stage2_17[33]}
   );
   gpc1_1 gpc1087 (
      {stage1_17[61]},
      {stage2_17[34]}
   );
   gpc1_1 gpc1088 (
      {stage1_17[62]},
      {stage2_17[35]}
   );
   gpc1_1 gpc1089 (
      {stage1_17[63]},
      {stage2_17[36]}
   );
   gpc1_1 gpc1090 (
      {stage1_19[66]},
      {stage2_19[27]}
   );
   gpc1_1 gpc1091 (
      {stage1_20[52]},
      {stage2_20[29]}
   );
   gpc1_1 gpc1092 (
      {stage1_20[53]},
      {stage2_20[30]}
   );
   gpc1_1 gpc1093 (
      {stage1_20[54]},
      {stage2_20[31]}
   );
   gpc1_1 gpc1094 (
      {stage1_20[55]},
      {stage2_20[32]}
   );
   gpc1_1 gpc1095 (
      {stage1_20[56]},
      {stage2_20[33]}
   );
   gpc1_1 gpc1096 (
      {stage1_20[57]},
      {stage2_20[34]}
   );
   gpc1_1 gpc1097 (
      {stage1_20[58]},
      {stage2_20[35]}
   );
   gpc1_1 gpc1098 (
      {stage1_20[59]},
      {stage2_20[36]}
   );
   gpc1_1 gpc1099 (
      {stage1_20[60]},
      {stage2_20[37]}
   );
   gpc1_1 gpc1100 (
      {stage1_22[78]},
      {stage2_22[30]}
   );
   gpc1_1 gpc1101 (
      {stage1_22[79]},
      {stage2_22[31]}
   );
   gpc1_1 gpc1102 (
      {stage1_22[80]},
      {stage2_22[32]}
   );
   gpc1_1 gpc1103 (
      {stage1_22[81]},
      {stage2_22[33]}
   );
   gpc1_1 gpc1104 (
      {stage1_23[78]},
      {stage2_23[31]}
   );
   gpc1_1 gpc1105 (
      {stage1_23[79]},
      {stage2_23[32]}
   );
   gpc1_1 gpc1106 (
      {stage1_23[80]},
      {stage2_23[33]}
   );
   gpc1_1 gpc1107 (
      {stage1_23[81]},
      {stage2_23[34]}
   );
   gpc1_1 gpc1108 (
      {stage1_23[82]},
      {stage2_23[35]}
   );
   gpc1_1 gpc1109 (
      {stage1_23[83]},
      {stage2_23[36]}
   );
   gpc1_1 gpc1110 (
      {stage1_23[84]},
      {stage2_23[37]}
   );
   gpc1_1 gpc1111 (
      {stage1_23[85]},
      {stage2_23[38]}
   );
   gpc1_1 gpc1112 (
      {stage1_23[86]},
      {stage2_23[39]}
   );
   gpc1_1 gpc1113 (
      {stage1_23[87]},
      {stage2_23[40]}
   );
   gpc1_1 gpc1114 (
      {stage1_23[88]},
      {stage2_23[41]}
   );
   gpc1_1 gpc1115 (
      {stage1_23[89]},
      {stage2_23[42]}
   );
   gpc1_1 gpc1116 (
      {stage1_23[90]},
      {stage2_23[43]}
   );
   gpc1_1 gpc1117 (
      {stage1_24[60]},
      {stage2_24[28]}
   );
   gpc1_1 gpc1118 (
      {stage1_24[61]},
      {stage2_24[29]}
   );
   gpc1_1 gpc1119 (
      {stage1_24[62]},
      {stage2_24[30]}
   );
   gpc1_1 gpc1120 (
      {stage1_24[63]},
      {stage2_24[31]}
   );
   gpc1_1 gpc1121 (
      {stage1_24[64]},
      {stage2_24[32]}
   );
   gpc1_1 gpc1122 (
      {stage1_24[65]},
      {stage2_24[33]}
   );
   gpc1_1 gpc1123 (
      {stage1_24[66]},
      {stage2_24[34]}
   );
   gpc1_1 gpc1124 (
      {stage1_26[54]},
      {stage2_26[30]}
   );
   gpc1_1 gpc1125 (
      {stage1_27[58]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1126 (
      {stage1_27[59]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1127 (
      {stage1_27[60]},
      {stage2_27[26]}
   );
   gpc1_1 gpc1128 (
      {stage1_27[61]},
      {stage2_27[27]}
   );
   gpc1_1 gpc1129 (
      {stage1_27[62]},
      {stage2_27[28]}
   );
   gpc1_1 gpc1130 (
      {stage1_27[63]},
      {stage2_27[29]}
   );
   gpc1_1 gpc1131 (
      {stage1_27[64]},
      {stage2_27[30]}
   );
   gpc1_1 gpc1132 (
      {stage1_27[65]},
      {stage2_27[31]}
   );
   gpc1_1 gpc1133 (
      {stage1_27[66]},
      {stage2_27[32]}
   );
   gpc1_1 gpc1134 (
      {stage1_28[72]},
      {stage2_28[24]}
   );
   gpc1_1 gpc1135 (
      {stage1_28[73]},
      {stage2_28[25]}
   );
   gpc1_1 gpc1136 (
      {stage1_28[74]},
      {stage2_28[26]}
   );
   gpc1_1 gpc1137 (
      {stage1_28[75]},
      {stage2_28[27]}
   );
   gpc1_1 gpc1138 (
      {stage1_28[76]},
      {stage2_28[28]}
   );
   gpc1_1 gpc1139 (
      {stage1_28[77]},
      {stage2_28[29]}
   );
   gpc1_1 gpc1140 (
      {stage1_30[55]},
      {stage2_30[29]}
   );
   gpc1_1 gpc1141 (
      {stage1_30[56]},
      {stage2_30[30]}
   );
   gpc1_1 gpc1142 (
      {stage1_30[57]},
      {stage2_30[31]}
   );
   gpc1_1 gpc1143 (
      {stage1_30[58]},
      {stage2_30[32]}
   );
   gpc1_1 gpc1144 (
      {stage1_30[59]},
      {stage2_30[33]}
   );
   gpc1_1 gpc1145 (
      {stage1_30[60]},
      {stage2_30[34]}
   );
   gpc1_1 gpc1146 (
      {stage1_30[61]},
      {stage2_30[35]}
   );
   gpc1_1 gpc1147 (
      {stage1_30[62]},
      {stage2_30[36]}
   );
   gpc1_1 gpc1148 (
      {stage1_31[87]},
      {stage2_31[25]}
   );
   gpc1_1 gpc1149 (
      {stage1_31[88]},
      {stage2_31[26]}
   );
   gpc1_1 gpc1150 (
      {stage1_31[89]},
      {stage2_31[27]}
   );
   gpc1_1 gpc1151 (
      {stage1_31[90]},
      {stage2_31[28]}
   );
   gpc1_1 gpc1152 (
      {stage1_31[91]},
      {stage2_31[29]}
   );
   gpc1_1 gpc1153 (
      {stage1_31[92]},
      {stage2_31[30]}
   );
   gpc1_1 gpc1154 (
      {stage1_31[93]},
      {stage2_31[31]}
   );
   gpc1_1 gpc1155 (
      {stage1_31[94]},
      {stage2_31[32]}
   );
   gpc1_1 gpc1156 (
      {stage1_31[95]},
      {stage2_31[33]}
   );
   gpc1_1 gpc1157 (
      {stage1_31[96]},
      {stage2_31[34]}
   );
   gpc1_1 gpc1158 (
      {stage1_31[97]},
      {stage2_31[35]}
   );
   gpc1_1 gpc1159 (
      {stage1_32[27]},
      {stage2_32[23]}
   );
   gpc1_1 gpc1160 (
      {stage1_32[28]},
      {stage2_32[24]}
   );
   gpc1_1 gpc1161 (
      {stage1_32[29]},
      {stage2_32[25]}
   );
   gpc1_1 gpc1162 (
      {stage1_32[30]},
      {stage2_32[26]}
   );
   gpc1_1 gpc1163 (
      {stage1_32[31]},
      {stage2_32[27]}
   );
   gpc1_1 gpc1164 (
      {stage1_32[32]},
      {stage2_32[28]}
   );
   gpc1_1 gpc1165 (
      {stage1_32[33]},
      {stage2_32[29]}
   );
   gpc1_1 gpc1166 (
      {stage1_32[34]},
      {stage2_32[30]}
   );
   gpc1_1 gpc1167 (
      {stage1_32[35]},
      {stage2_32[31]}
   );
   gpc1_1 gpc1168 (
      {stage1_32[36]},
      {stage2_32[32]}
   );
   gpc1_1 gpc1169 (
      {stage1_32[37]},
      {stage2_32[33]}
   );
   gpc1_1 gpc1170 (
      {stage1_32[38]},
      {stage2_32[34]}
   );
   gpc1_1 gpc1171 (
      {stage1_32[39]},
      {stage2_32[35]}
   );
   gpc1_1 gpc1172 (
      {stage1_32[40]},
      {stage2_32[36]}
   );
   gpc1_1 gpc1173 (
      {stage1_32[41]},
      {stage2_32[37]}
   );
   gpc1_1 gpc1174 (
      {stage1_32[42]},
      {stage2_32[38]}
   );
   gpc1_1 gpc1175 (
      {stage1_32[43]},
      {stage2_32[39]}
   );
   gpc1_1 gpc1176 (
      {stage1_32[44]},
      {stage2_32[40]}
   );
   gpc1_1 gpc1177 (
      {stage1_33[13]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1178 (
      {stage1_33[14]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1179 (
      {stage1_33[15]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1180 (
      {stage1_33[16]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1181 (
      {stage1_33[17]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1182 (
      {stage1_33[18]},
      {stage2_33[23]}
   );
   gpc135_4 gpc1183 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1184 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc1185 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1186 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[3],stage3_2[3]}
   );
   gpc1163_5 gpc1187 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[4]}
   );
   gpc1163_5 gpc1188 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[5]}
   );
   gpc1163_5 gpc1189 (
      {stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage2_5[2]},
      {stage2_6[2]},
      {stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5],stage3_3[6]}
   );
   gpc623_5 gpc1190 (
      {stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_4[30], stage2_4[31]},
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage3_7[3],stage3_6[5],stage3_5[6],stage3_4[6],stage3_3[7]}
   );
   gpc615_5 gpc1191 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[9]},
      {stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage3_8[0],stage3_7[4],stage3_6[6],stage3_5[7],stage3_4[7]}
   );
   gpc615_5 gpc1192 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], 1'b0},
      {stage2_5[10]},
      {stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14]},
      {stage3_8[1],stage3_7[5],stage3_6[7],stage3_5[8],stage3_4[8]}
   );
   gpc606_5 gpc1193 (
      {stage2_5[11], stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc1194 (
      {stage2_5[17], stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[7],stage3_6[9],stage3_5[10]}
   );
   gpc606_5 gpc1195 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], 1'b0},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[4],stage3_7[8],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc1196 (
      {stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[5],stage3_7[9],stage3_6[11]}
   );
   gpc606_5 gpc1197 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[4],stage3_8[6],stage3_7[10],stage3_6[12]}
   );
   gpc615_5 gpc1198 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[5],stage3_8[7],stage3_7[11]}
   );
   gpc615_5 gpc1199 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[6],stage3_8[8],stage3_7[12]}
   );
   gpc606_5 gpc1200 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[4],stage3_9[7],stage3_8[9]}
   );
   gpc606_5 gpc1201 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[5],stage3_9[8],stage3_8[10]}
   );
   gpc1343_5 gpc1202 (
      {stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15]},
      {stage2_11[0], stage2_11[1], stage2_11[2]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[4],stage3_10[6],stage3_9[9]}
   );
   gpc1343_5 gpc1203 (
      {stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[3],stage3_11[5],stage3_10[7],stage3_9[10]}
   );
   gpc1343_5 gpc1204 (
      {stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[4],stage3_11[6],stage3_10[8],stage3_9[11]}
   );
   gpc1343_5 gpc1205 (
      {stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27]},
      {stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[5],stage3_11[7],stage3_10[9],stage3_9[12]}
   );
   gpc1343_5 gpc1206 (
      {stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31]},
      {stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[4]},
      {stage3_13[4],stage3_12[6],stage3_11[8],stage3_10[10],stage3_9[13]}
   );
   gpc606_5 gpc1207 (
      {stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37]},
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage3_14[0],stage3_13[5],stage3_12[7],stage3_11[9],stage3_10[11]}
   );
   gpc606_5 gpc1208 (
      {stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43]},
      {stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16]},
      {stage3_14[1],stage3_13[6],stage3_12[8],stage3_11[10],stage3_10[12]}
   );
   gpc606_5 gpc1209 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[7],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc1210 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[8],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc1211 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[9],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc1212 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[10],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc1213 (
      {stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[6],stage3_13[11],stage3_12[13]}
   );
   gpc606_5 gpc1214 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[5],stage3_14[7],stage3_13[12]}
   );
   gpc606_5 gpc1215 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[2],stage3_15[6],stage3_14[8],stage3_13[13]}
   );
   gpc606_5 gpc1216 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[3],stage3_15[7],stage3_14[9],stage3_13[14]}
   );
   gpc615_5 gpc1217 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[18]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[4],stage3_15[8],stage3_14[10]}
   );
   gpc615_5 gpc1218 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[19]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[4],stage3_16[5],stage3_15[9],stage3_14[11]}
   );
   gpc615_5 gpc1219 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[20]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[5],stage3_16[6],stage3_15[10],stage3_14[12]}
   );
   gpc615_5 gpc1220 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[21]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[6],stage3_16[7],stage3_15[11],stage3_14[13]}
   );
   gpc615_5 gpc1221 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[22]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[7],stage3_16[8],stage3_15[12],stage3_14[14]}
   );
   gpc615_5 gpc1222 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[23]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[8],stage3_16[9],stage3_15[13],stage3_14[15]}
   );
   gpc615_5 gpc1223 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[9],stage3_16[10],stage3_15[14]}
   );
   gpc615_5 gpc1224 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[37]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[7],stage3_17[10],stage3_16[11],stage3_15[15]}
   );
   gpc606_5 gpc1225 (
      {stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41], stage2_16[42], stage2_16[43]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[8],stage3_17[11],stage3_16[12]}
   );
   gpc606_5 gpc1226 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[9],stage3_17[12]}
   );
   gpc606_5 gpc1227 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[10],stage3_17[13]}
   );
   gpc606_5 gpc1228 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[5],stage3_18[11],stage3_17[14]}
   );
   gpc606_5 gpc1229 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[6],stage3_18[12],stage3_17[15]}
   );
   gpc606_5 gpc1230 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[4],stage3_20[5],stage3_19[7],stage3_18[13]}
   );
   gpc606_5 gpc1231 (
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[5],stage3_20[6],stage3_19[8],stage3_18[14]}
   );
   gpc606_5 gpc1232 (
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[6],stage3_20[7],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc1233 (
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28]},
      {stage2_19[24]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[7],stage3_20[8],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc1234 (
      {stage2_19[25], stage2_19[26], stage2_19[27], 1'b0, 1'b0},
      {stage2_20[24]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[4],stage3_21[8],stage3_20[9],stage3_19[11]}
   );
   gpc606_5 gpc1235 (
      {stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[1],stage3_22[5],stage3_21[9],stage3_20[10]}
   );
   gpc615_5 gpc1236 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10]},
      {stage2_22[6]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[2],stage3_22[6],stage3_21[10]}
   );
   gpc615_5 gpc1237 (
      {stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage2_22[7]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[3],stage3_22[7],stage3_21[11]}
   );
   gpc615_5 gpc1238 (
      {stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20]},
      {stage2_22[8]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[3],stage3_23[4],stage3_22[8],stage3_21[12]}
   );
   gpc615_5 gpc1239 (
      {stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24], stage2_21[25]},
      {stage2_22[9]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[4],stage3_23[5],stage3_22[9],stage3_21[13]}
   );
   gpc615_5 gpc1240 (
      {stage2_21[26], stage2_21[27], 1'b0, 1'b0, 1'b0},
      {stage2_22[10]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[5],stage3_23[6],stage3_22[10],stage3_21[14]}
   );
   gpc207_4 gpc1241 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[0], stage2_24[1]},
      {stage3_25[5],stage3_24[6],stage3_23[7],stage3_22[11]}
   );
   gpc606_5 gpc1242 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7]},
      {stage3_26[0],stage3_25[6],stage3_24[7],stage3_23[8],stage3_22[12]}
   );
   gpc606_5 gpc1243 (
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[1],stage3_25[7],stage3_24[8],stage3_23[9]}
   );
   gpc606_5 gpc1244 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[2],stage3_25[8],stage3_24[9],stage3_23[10]}
   );
   gpc606_5 gpc1245 (
      {stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[2],stage3_26[3],stage3_25[9],stage3_24[10]}
   );
   gpc606_5 gpc1246 (
      {stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[3],stage3_26[4],stage3_25[10],stage3_24[11]}
   );
   gpc606_5 gpc1247 (
      {stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[4],stage3_26[5],stage3_25[11],stage3_24[12]}
   );
   gpc606_5 gpc1248 (
      {stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[5],stage3_26[6],stage3_25[12],stage3_24[13]}
   );
   gpc606_5 gpc1249 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[4],stage3_27[6],stage3_26[7],stage3_25[13]}
   );
   gpc606_5 gpc1250 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[5],stage3_27[7],stage3_26[8],stage3_25[14]}
   );
   gpc606_5 gpc1251 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[6],stage3_27[8],stage3_26[9],stage3_25[15]}
   );
   gpc606_5 gpc1252 (
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[3],stage3_28[7],stage3_27[9],stage3_26[10]}
   );
   gpc615_5 gpc1253 (
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22]},
      {stage2_28[6]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[1],stage3_29[4],stage3_28[8],stage3_27[10]}
   );
   gpc615_5 gpc1254 (
      {stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27]},
      {stage2_28[7]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[2],stage3_29[5],stage3_28[9],stage3_27[11]}
   );
   gpc615_5 gpc1255 (
      {stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[8]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[3],stage3_29[6],stage3_28[10],stage3_27[12]}
   );
   gpc135_4 gpc1256 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[18], stage2_29[19], stage2_29[20]},
      {stage2_30[0]},
      {stage3_31[3],stage3_30[4],stage3_29[7],stage3_28[11]}
   );
   gpc606_5 gpc1257 (
      {stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19]},
      {stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5], stage2_30[6]},
      {stage3_32[0],stage3_31[4],stage3_30[5],stage3_29[8],stage3_28[12]}
   );
   gpc606_5 gpc1258 (
      {stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24], stage2_29[25], stage2_29[26]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[1],stage3_31[5],stage3_30[6],stage3_29[9]}
   );
   gpc606_5 gpc1259 (
      {stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[2],stage3_31[6],stage3_30[7],stage3_29[10]}
   );
   gpc615_5 gpc1260 (
      {stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[3],stage3_31[7],stage3_30[8]}
   );
   gpc615_5 gpc1261 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[4],stage3_31[8],stage3_30[9]}
   );
   gpc615_5 gpc1262 (
      {stage2_30[17], stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21]},
      {stage2_31[14]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[4],stage3_32[5],stage3_31[9],stage3_30[10]}
   );
   gpc615_5 gpc1263 (
      {stage2_30[22], stage2_30[23], stage2_30[24], stage2_30[25], stage2_30[26]},
      {stage2_31[15]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[5],stage3_32[6],stage3_31[10],stage3_30[11]}
   );
   gpc615_5 gpc1264 (
      {stage2_30[27], stage2_30[28], stage2_30[29], stage2_30[30], stage2_30[31]},
      {stage2_31[16]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[6],stage3_32[7],stage3_31[11],stage3_30[12]}
   );
   gpc615_5 gpc1265 (
      {stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35], stage2_30[36]},
      {stage2_31[17]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[7],stage3_32[8],stage3_31[12],stage3_30[13]}
   );
   gpc606_5 gpc1266 (
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[6],stage3_33[8],stage3_32[9],stage3_31[13]}
   );
   gpc606_5 gpc1267 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[7],stage3_33[9],stage3_32[10],stage3_31[14]}
   );
   gpc615_5 gpc1268 (
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage2_32[36]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[8],stage3_33[10],stage3_32[11],stage3_31[15]}
   );
   gpc1_1 gpc1269 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1270 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1271 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1272 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1273 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1274 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1275 (
      {stage2_1[9]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1276 (
      {stage2_1[10]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_1[11]},
      {stage3_1[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_1[12]},
      {stage3_1[5]}
   );
   gpc1_1 gpc1279 (
      {stage2_1[13]},
      {stage3_1[6]}
   );
   gpc1_1 gpc1280 (
      {stage2_1[14]},
      {stage3_1[7]}
   );
   gpc1_1 gpc1281 (
      {stage2_1[15]},
      {stage3_1[8]}
   );
   gpc1_1 gpc1282 (
      {stage2_1[16]},
      {stage3_1[9]}
   );
   gpc1_1 gpc1283 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1284 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc1285 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc1286 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc1287 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc1288 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc1289 (
      {stage2_3[20]},
      {stage3_3[8]}
   );
   gpc1_1 gpc1290 (
      {stage2_3[21]},
      {stage3_3[9]}
   );
   gpc1_1 gpc1291 (
      {stage2_3[22]},
      {stage3_3[10]}
   );
   gpc1_1 gpc1292 (
      {stage2_3[23]},
      {stage3_3[11]}
   );
   gpc1_1 gpc1293 (
      {stage2_3[24]},
      {stage3_3[12]}
   );
   gpc1_1 gpc1294 (
      {stage2_3[25]},
      {stage3_3[13]}
   );
   gpc1_1 gpc1295 (
      {stage2_3[26]},
      {stage3_3[14]}
   );
   gpc1_1 gpc1296 (
      {stage2_3[27]},
      {stage3_3[15]}
   );
   gpc1_1 gpc1297 (
      {stage2_3[28]},
      {stage3_3[16]}
   );
   gpc1_1 gpc1298 (
      {stage2_3[29]},
      {stage3_3[17]}
   );
   gpc1_1 gpc1299 (
      {stage2_3[30]},
      {stage3_3[18]}
   );
   gpc1_1 gpc1300 (
      {stage2_3[31]},
      {stage3_3[19]}
   );
   gpc1_1 gpc1301 (
      {stage2_3[32]},
      {stage3_3[20]}
   );
   gpc1_1 gpc1302 (
      {stage2_3[33]},
      {stage3_3[21]}
   );
   gpc1_1 gpc1303 (
      {stage2_3[34]},
      {stage3_3[22]}
   );
   gpc1_1 gpc1304 (
      {stage2_6[27]},
      {stage3_6[13]}
   );
   gpc1_1 gpc1305 (
      {stage2_6[28]},
      {stage3_6[14]}
   );
   gpc1_1 gpc1306 (
      {stage2_6[29]},
      {stage3_6[15]}
   );
   gpc1_1 gpc1307 (
      {stage2_6[30]},
      {stage3_6[16]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[28]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[29]},
      {stage3_7[14]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[30]},
      {stage3_7[15]}
   );
   gpc1_1 gpc1311 (
      {stage2_7[31]},
      {stage3_7[16]}
   );
   gpc1_1 gpc1312 (
      {stage2_7[32]},
      {stage3_7[17]}
   );
   gpc1_1 gpc1313 (
      {stage2_7[33]},
      {stage3_7[18]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc1315 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc1316 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc1317 (
      {stage2_8[29]},
      {stage3_8[14]}
   );
   gpc1_1 gpc1318 (
      {stage2_8[30]},
      {stage3_8[15]}
   );
   gpc1_1 gpc1319 (
      {stage2_8[31]},
      {stage3_8[16]}
   );
   gpc1_1 gpc1320 (
      {stage2_8[32]},
      {stage3_8[17]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[27]},
      {stage3_9[14]}
   );
   gpc1_1 gpc1322 (
      {stage2_9[28]},
      {stage3_9[15]}
   );
   gpc1_1 gpc1323 (
      {stage2_9[29]},
      {stage3_9[16]}
   );
   gpc1_1 gpc1324 (
      {stage2_9[30]},
      {stage3_9[17]}
   );
   gpc1_1 gpc1325 (
      {stage2_9[31]},
      {stage3_9[18]}
   );
   gpc1_1 gpc1326 (
      {stage2_10[44]},
      {stage3_10[13]}
   );
   gpc1_1 gpc1327 (
      {stage2_10[45]},
      {stage3_10[14]}
   );
   gpc1_1 gpc1328 (
      {stage2_12[23]},
      {stage3_12[14]}
   );
   gpc1_1 gpc1329 (
      {stage2_13[42]},
      {stage3_13[15]}
   );
   gpc1_1 gpc1330 (
      {stage2_13[43]},
      {stage3_13[16]}
   );
   gpc1_1 gpc1331 (
      {stage2_13[44]},
      {stage3_13[17]}
   );
   gpc1_1 gpc1332 (
      {stage2_14[36]},
      {stage3_14[16]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[36]},
      {stage3_17[16]}
   );
   gpc1_1 gpc1334 (
      {stage2_20[31]},
      {stage3_20[11]}
   );
   gpc1_1 gpc1335 (
      {stage2_20[32]},
      {stage3_20[12]}
   );
   gpc1_1 gpc1336 (
      {stage2_20[33]},
      {stage3_20[13]}
   );
   gpc1_1 gpc1337 (
      {stage2_20[34]},
      {stage3_20[14]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[35]},
      {stage3_20[15]}
   );
   gpc1_1 gpc1339 (
      {stage2_20[36]},
      {stage3_20[16]}
   );
   gpc1_1 gpc1340 (
      {stage2_20[37]},
      {stage3_20[17]}
   );
   gpc1_1 gpc1341 (
      {stage2_22[24]},
      {stage3_22[13]}
   );
   gpc1_1 gpc1342 (
      {stage2_22[25]},
      {stage3_22[14]}
   );
   gpc1_1 gpc1343 (
      {stage2_22[26]},
      {stage3_22[15]}
   );
   gpc1_1 gpc1344 (
      {stage2_22[27]},
      {stage3_22[16]}
   );
   gpc1_1 gpc1345 (
      {stage2_22[28]},
      {stage3_22[17]}
   );
   gpc1_1 gpc1346 (
      {stage2_22[29]},
      {stage3_22[18]}
   );
   gpc1_1 gpc1347 (
      {stage2_22[30]},
      {stage3_22[19]}
   );
   gpc1_1 gpc1348 (
      {stage2_22[31]},
      {stage3_22[20]}
   );
   gpc1_1 gpc1349 (
      {stage2_22[32]},
      {stage3_22[21]}
   );
   gpc1_1 gpc1350 (
      {stage2_22[33]},
      {stage3_22[22]}
   );
   gpc1_1 gpc1351 (
      {stage2_23[42]},
      {stage3_23[11]}
   );
   gpc1_1 gpc1352 (
      {stage2_23[43]},
      {stage3_23[12]}
   );
   gpc1_1 gpc1353 (
      {stage2_24[32]},
      {stage3_24[14]}
   );
   gpc1_1 gpc1354 (
      {stage2_24[33]},
      {stage3_24[15]}
   );
   gpc1_1 gpc1355 (
      {stage2_24[34]},
      {stage3_24[16]}
   );
   gpc1_1 gpc1356 (
      {stage2_25[30]},
      {stage3_25[16]}
   );
   gpc1_1 gpc1357 (
      {stage2_26[30]},
      {stage3_26[11]}
   );
   gpc1_1 gpc1358 (
      {stage2_28[20]},
      {stage3_28[13]}
   );
   gpc1_1 gpc1359 (
      {stage2_28[21]},
      {stage3_28[14]}
   );
   gpc1_1 gpc1360 (
      {stage2_28[22]},
      {stage3_28[15]}
   );
   gpc1_1 gpc1361 (
      {stage2_28[23]},
      {stage3_28[16]}
   );
   gpc1_1 gpc1362 (
      {stage2_28[24]},
      {stage3_28[17]}
   );
   gpc1_1 gpc1363 (
      {stage2_28[25]},
      {stage3_28[18]}
   );
   gpc1_1 gpc1364 (
      {stage2_28[26]},
      {stage3_28[19]}
   );
   gpc1_1 gpc1365 (
      {stage2_28[27]},
      {stage3_28[20]}
   );
   gpc1_1 gpc1366 (
      {stage2_28[28]},
      {stage3_28[21]}
   );
   gpc1_1 gpc1367 (
      {stage2_28[29]},
      {stage3_28[22]}
   );
   gpc1_1 gpc1368 (
      {stage2_31[35]},
      {stage3_31[16]}
   );
   gpc1_1 gpc1369 (
      {stage2_32[37]},
      {stage3_32[12]}
   );
   gpc1_1 gpc1370 (
      {stage2_32[38]},
      {stage3_32[13]}
   );
   gpc1_1 gpc1371 (
      {stage2_32[39]},
      {stage3_32[14]}
   );
   gpc1_1 gpc1372 (
      {stage2_32[40]},
      {stage3_32[15]}
   );
   gpc1_1 gpc1373 (
      {stage2_33[18]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1374 (
      {stage2_33[19]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1375 (
      {stage2_33[20]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1376 (
      {stage2_33[21]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1377 (
      {stage2_33[22]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1378 (
      {stage2_33[23]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1379 (
      {stage2_34[0]},
      {stage3_34[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_34[1]},
      {stage3_34[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_34[2]},
      {stage3_34[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_34[3]},
      {stage3_34[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_34[4]},
      {stage3_34[13]}
   );
   gpc1_1 gpc1384 (
      {stage2_34[5]},
      {stage3_34[14]}
   );
   gpc1_1 gpc1385 (
      {stage2_34[6]},
      {stage3_34[15]}
   );
   gpc1_1 gpc1386 (
      {stage2_35[0]},
      {stage3_35[3]}
   );
   gpc1_1 gpc1387 (
      {stage2_35[1]},
      {stage3_35[4]}
   );
   gpc606_5 gpc1388 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1389 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1390 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc1391 (
      {stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage3_4[1]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc1392 (
      {stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6], stage3_4[7]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc1393 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[3]}
   );
   gpc615_5 gpc1394 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[4]}
   );
   gpc1406_5 gpc1395 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc1396 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[4],stage4_7[6]}
   );
   gpc615_5 gpc1397 (
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18]},
      {stage3_8[12]},
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage4_11[2],stage4_10[4],stage4_9[4],stage4_8[5],stage4_7[7]}
   );
   gpc615_5 gpc1398 (
      {stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_9[16]},
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[5],stage4_8[6]}
   );
   gpc7_3 gpc1399 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[4],stage4_10[6]}
   );
   gpc606_5 gpc1400 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[2],stage4_11[5]}
   );
   gpc606_5 gpc1401 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[1],stage4_13[1],stage4_12[3],stage4_11[6]}
   );
   gpc606_5 gpc1402 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[2],stage4_13[2],stage4_12[4]}
   );
   gpc606_5 gpc1403 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[3],stage4_13[3],stage4_12[5]}
   );
   gpc606_5 gpc1404 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[2],stage4_15[4],stage4_14[4],stage4_13[4]}
   );
   gpc615_5 gpc1405 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[3],stage4_15[5],stage4_14[5]}
   );
   gpc606_5 gpc1406 (
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[2],stage4_16[4],stage4_15[6]}
   );
   gpc606_5 gpc1407 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[1],stage4_18[2],stage4_17[3],stage4_16[5]}
   );
   gpc1163_5 gpc1408 (
      {stage3_17[6], stage3_17[7], stage3_17[8]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[1],stage4_19[2],stage4_18[3],stage4_17[4]}
   );
   gpc1343_5 gpc1409 (
      {stage3_19[1], stage3_19[2], stage3_19[3]},
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[0], stage3_21[1], stage3_21[2]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[1],stage4_20[2],stage4_19[3]}
   );
   gpc606_5 gpc1410 (
      {stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[2],stage4_20[3]}
   );
   gpc606_5 gpc1411 (
      {stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16]},
      {stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[3],stage4_20[4]}
   );
   gpc606_5 gpc1412 (
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[4]}
   );
   gpc606_5 gpc1413 (
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[5]}
   );
   gpc207_4 gpc1414 (
      {stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[2],stage4_24[4],stage4_23[5],stage4_22[5]}
   );
   gpc2135_5 gpc1415 (
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1]},
      {stage4_28[0],stage4_27[0],stage4_26[0],stage4_25[3],stage4_24[5]}
   );
   gpc2135_5 gpc1416 (
      {stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage3_26[1]},
      {stage3_27[2], stage3_27[3]},
      {stage4_28[1],stage4_27[1],stage4_26[1],stage4_25[4],stage4_24[6]}
   );
   gpc2135_5 gpc1417 (
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16]},
      {stage3_25[6], stage3_25[7], stage3_25[8]},
      {stage3_26[2]},
      {stage3_27[4], stage3_27[5]},
      {stage4_28[2],stage4_27[2],stage4_26[2],stage4_25[5],stage4_24[7]}
   );
   gpc606_5 gpc1418 (
      {stage3_25[9], stage3_25[10], stage3_25[11], stage3_25[12], stage3_25[13], stage3_25[14]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[0],stage4_28[3],stage4_27[3],stage4_26[3],stage4_25[6]}
   );
   gpc615_5 gpc1419 (
      {stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7]},
      {stage3_27[12]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[1],stage4_28[4],stage4_27[4],stage4_26[4]}
   );
   gpc2135_5 gpc1420 (
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[2],stage4_28[5]}
   );
   gpc2135_5 gpc1421 (
      {stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15]},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[3],stage4_28[6]}
   );
   gpc606_5 gpc1422 (
      {stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7]},
      {stage4_32[2],stage4_31[2],stage4_30[3],stage4_29[4],stage4_28[7]}
   );
   gpc615_5 gpc1423 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10]},
      {stage3_30[8]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[0],stage4_32[3],stage4_31[3],stage4_30[4],stage4_29[5]}
   );
   gpc615_5 gpc1424 (
      {stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13]},
      {stage3_31[10]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[4],stage4_31[4],stage4_30[5]}
   );
   gpc606_5 gpc1425 (
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[2],stage4_32[5],stage4_31[5]}
   );
   gpc606_5 gpc1426 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[1],stage4_34[2],stage4_33[3],stage4_32[6]}
   );
   gpc1163_5 gpc1427 (
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage3_35[0]},
      {1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1428 (
      {stage3_33[9], stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], 1'b0, 1'b0},
      {stage4_37[1],stage4_36[2],stage4_35[3],stage4_34[4],stage4_33[5]}
   );
   gpc1_1 gpc1429 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1430 (
      {stage3_1[6]},
      {stage4_1[2]}
   );
   gpc1_1 gpc1431 (
      {stage3_1[7]},
      {stage4_1[3]}
   );
   gpc1_1 gpc1432 (
      {stage3_1[8]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1433 (
      {stage3_1[9]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1434 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1435 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc1436 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1437 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1438 (
      {stage3_3[16]},
      {stage4_3[4]}
   );
   gpc1_1 gpc1439 (
      {stage3_3[17]},
      {stage4_3[5]}
   );
   gpc1_1 gpc1440 (
      {stage3_3[18]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1441 (
      {stage3_3[19]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1442 (
      {stage3_3[20]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1443 (
      {stage3_3[21]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1444 (
      {stage3_3[22]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1445 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1446 (
      {stage3_6[16]},
      {stage4_6[5]}
   );
   gpc1_1 gpc1447 (
      {stage3_9[17]},
      {stage4_9[6]}
   );
   gpc1_1 gpc1448 (
      {stage3_9[18]},
      {stage4_9[7]}
   );
   gpc1_1 gpc1449 (
      {stage3_10[14]},
      {stage4_10[7]}
   );
   gpc1_1 gpc1450 (
      {stage3_11[12]},
      {stage4_11[7]}
   );
   gpc1_1 gpc1451 (
      {stage3_11[13]},
      {stage4_11[8]}
   );
   gpc1_1 gpc1452 (
      {stage3_11[14]},
      {stage4_11[9]}
   );
   gpc1_1 gpc1453 (
      {stage3_12[12]},
      {stage4_12[6]}
   );
   gpc1_1 gpc1454 (
      {stage3_12[13]},
      {stage4_12[7]}
   );
   gpc1_1 gpc1455 (
      {stage3_12[14]},
      {stage4_12[8]}
   );
   gpc1_1 gpc1456 (
      {stage3_15[13]},
      {stage4_15[7]}
   );
   gpc1_1 gpc1457 (
      {stage3_15[14]},
      {stage4_15[8]}
   );
   gpc1_1 gpc1458 (
      {stage3_15[15]},
      {stage4_15[9]}
   );
   gpc1_1 gpc1459 (
      {stage3_16[12]},
      {stage4_16[6]}
   );
   gpc1_1 gpc1460 (
      {stage3_17[9]},
      {stage4_17[5]}
   );
   gpc1_1 gpc1461 (
      {stage3_17[10]},
      {stage4_17[6]}
   );
   gpc1_1 gpc1462 (
      {stage3_17[11]},
      {stage4_17[7]}
   );
   gpc1_1 gpc1463 (
      {stage3_17[12]},
      {stage4_17[8]}
   );
   gpc1_1 gpc1464 (
      {stage3_17[13]},
      {stage4_17[9]}
   );
   gpc1_1 gpc1465 (
      {stage3_17[14]},
      {stage4_17[10]}
   );
   gpc1_1 gpc1466 (
      {stage3_17[15]},
      {stage4_17[11]}
   );
   gpc1_1 gpc1467 (
      {stage3_17[16]},
      {stage4_17[12]}
   );
   gpc1_1 gpc1468 (
      {stage3_18[12]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1469 (
      {stage3_18[13]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1470 (
      {stage3_18[14]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1471 (
      {stage3_18[15]},
      {stage4_18[7]}
   );
   gpc1_1 gpc1472 (
      {stage3_18[16]},
      {stage4_18[8]}
   );
   gpc1_1 gpc1473 (
      {stage3_19[4]},
      {stage4_19[4]}
   );
   gpc1_1 gpc1474 (
      {stage3_19[5]},
      {stage4_19[5]}
   );
   gpc1_1 gpc1475 (
      {stage3_19[6]},
      {stage4_19[6]}
   );
   gpc1_1 gpc1476 (
      {stage3_19[7]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1477 (
      {stage3_19[8]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1478 (
      {stage3_19[9]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1479 (
      {stage3_19[10]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1480 (
      {stage3_19[11]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1481 (
      {stage3_20[17]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1482 (
      {stage3_22[20]},
      {stage4_22[6]}
   );
   gpc1_1 gpc1483 (
      {stage3_22[21]},
      {stage4_22[7]}
   );
   gpc1_1 gpc1484 (
      {stage3_22[22]},
      {stage4_22[8]}
   );
   gpc1_1 gpc1485 (
      {stage3_23[12]},
      {stage4_23[6]}
   );
   gpc1_1 gpc1486 (
      {stage3_25[15]},
      {stage4_25[7]}
   );
   gpc1_1 gpc1487 (
      {stage3_25[16]},
      {stage4_25[8]}
   );
   gpc1_1 gpc1488 (
      {stage3_26[8]},
      {stage4_26[5]}
   );
   gpc1_1 gpc1489 (
      {stage3_26[9]},
      {stage4_26[6]}
   );
   gpc1_1 gpc1490 (
      {stage3_26[10]},
      {stage4_26[7]}
   );
   gpc1_1 gpc1491 (
      {stage3_26[11]},
      {stage4_26[8]}
   );
   gpc1_1 gpc1492 (
      {stage3_28[22]},
      {stage4_28[8]}
   );
   gpc1_1 gpc1493 (
      {stage3_32[12]},
      {stage4_32[7]}
   );
   gpc1_1 gpc1494 (
      {stage3_32[13]},
      {stage4_32[8]}
   );
   gpc1_1 gpc1495 (
      {stage3_32[14]},
      {stage4_32[9]}
   );
   gpc1_1 gpc1496 (
      {stage3_32[15]},
      {stage4_32[10]}
   );
   gpc1_1 gpc1497 (
      {stage3_33[15]},
      {stage4_33[6]}
   );
   gpc1_1 gpc1498 (
      {stage3_33[16]},
      {stage4_33[7]}
   );
   gpc1_1 gpc1499 (
      {stage3_34[12]},
      {stage4_34[5]}
   );
   gpc1_1 gpc1500 (
      {stage3_34[13]},
      {stage4_34[6]}
   );
   gpc1_1 gpc1501 (
      {stage3_34[14]},
      {stage4_34[7]}
   );
   gpc1_1 gpc1502 (
      {stage3_34[15]},
      {stage4_34[8]}
   );
   gpc623_5 gpc1503 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1163_5 gpc1504 (
      {stage4_3[6], stage4_3[7], stage4_3[8]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1415_5 gpc1505 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1]}
   );
   gpc223_4 gpc1506 (
      {stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[4], stage4_8[5]},
      {stage4_9[1], stage4_9[2]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[2]}
   );
   gpc2135_5 gpc1507 (
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc615_5 gpc1508 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc615_5 gpc1509 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[8]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], 1'b0},
      {stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2],stage5_11[2]}
   );
   gpc1163_5 gpc1510 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc606_5 gpc1511 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc615_5 gpc1512 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_18[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[2],stage5_17[2]}
   );
   gpc615_5 gpc1513 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10]},
      {stage4_18[7]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[2],stage5_19[2],stage5_18[3],stage5_17[3]}
   );
   gpc606_5 gpc1514 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[2],stage5_20[3]}
   );
   gpc135_4 gpc1515 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[0]},
      {stage5_24[1],stage5_23[1],stage5_22[1],stage5_21[3]}
   );
   gpc615_5 gpc1516 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[2],stage5_23[2]}
   );
   gpc2135_5 gpc1517 (
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_26[0]},
      {stage4_27[0], stage4_27[1]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[3]}
   );
   gpc2223_5 gpc1518 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[2]}
   );
   gpc615_5 gpc1519 (
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8]},
      {stage4_27[4]},
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[3],stage5_26[3]}
   );
   gpc606_5 gpc1520 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[2]}
   );
   gpc606_5 gpc1521 (
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[1],stage5_33[1],stage5_32[1],stage5_31[1]}
   );
   gpc606_5 gpc1522 (
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], 1'b0},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[1],stage5_34[2],stage5_33[2],stage5_32[2]}
   );
   gpc2116_5 gpc1523 (
      {stage4_34[6], stage4_34[7], stage4_34[8], 1'b0, 1'b0, 1'b0},
      {stage4_35[0]},
      {stage4_36[0]},
      {stage4_37[0], stage4_37[1]},
      {stage5_38[0],stage5_37[0],stage5_36[1],stage5_35[2],stage5_34[3]}
   );
   gpc1_1 gpc1524 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1525 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1526 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1527 (
      {stage4_1[4]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1528 (
      {stage4_1[5]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1529 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc1530 (
      {stage4_2[3]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1531 (
      {stage4_2[4]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1532 (
      {stage4_2[5]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1533 (
      {stage4_3[9]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1534 (
      {stage4_3[10]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1535 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc1536 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc1537 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc1538 (
      {stage4_7[4]},
      {stage5_7[3]}
   );
   gpc1_1 gpc1539 (
      {stage4_7[5]},
      {stage5_7[4]}
   );
   gpc1_1 gpc1540 (
      {stage4_7[6]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1541 (
      {stage4_7[7]},
      {stage5_7[6]}
   );
   gpc1_1 gpc1542 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc1543 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc1544 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc1545 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc1546 (
      {stage4_14[3]},
      {stage5_14[3]}
   );
   gpc1_1 gpc1547 (
      {stage4_14[4]},
      {stage5_14[4]}
   );
   gpc1_1 gpc1548 (
      {stage4_14[5]},
      {stage5_14[5]}
   );
   gpc1_1 gpc1549 (
      {stage4_15[6]},
      {stage5_15[2]}
   );
   gpc1_1 gpc1550 (
      {stage4_15[7]},
      {stage5_15[3]}
   );
   gpc1_1 gpc1551 (
      {stage4_15[8]},
      {stage5_15[4]}
   );
   gpc1_1 gpc1552 (
      {stage4_15[9]},
      {stage5_15[5]}
   );
   gpc1_1 gpc1553 (
      {stage4_17[11]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1554 (
      {stage4_17[12]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1555 (
      {stage4_18[8]},
      {stage5_18[4]}
   );
   gpc1_1 gpc1556 (
      {stage4_21[5]},
      {stage5_21[4]}
   );
   gpc1_1 gpc1557 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc1558 (
      {stage4_24[6]},
      {stage5_24[4]}
   );
   gpc1_1 gpc1559 (
      {stage4_24[7]},
      {stage5_24[5]}
   );
   gpc1_1 gpc1560 (
      {stage4_28[8]},
      {stage5_28[3]}
   );
   gpc1_1 gpc1561 (
      {stage4_29[2]},
      {stage5_29[2]}
   );
   gpc1_1 gpc1562 (
      {stage4_29[3]},
      {stage5_29[3]}
   );
   gpc1_1 gpc1563 (
      {stage4_29[4]},
      {stage5_29[4]}
   );
   gpc1_1 gpc1564 (
      {stage4_29[5]},
      {stage5_29[5]}
   );
   gpc1_1 gpc1565 (
      {stage4_33[6]},
      {stage5_33[3]}
   );
   gpc1_1 gpc1566 (
      {stage4_33[7]},
      {stage5_33[4]}
   );
   gpc1_1 gpc1567 (
      {stage4_35[1]},
      {stage5_35[3]}
   );
   gpc1_1 gpc1568 (
      {stage4_35[2]},
      {stage5_35[4]}
   );
   gpc1_1 gpc1569 (
      {stage4_35[3]},
      {stage5_35[5]}
   );
   gpc1_1 gpc1570 (
      {stage4_36[1]},
      {stage5_36[2]}
   );
   gpc1_1 gpc1571 (
      {stage4_36[2]},
      {stage5_36[3]}
   );
   gpc1343_5 gpc1572 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc1573 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1]}
   );
   gpc1343_5 gpc1574 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc135_4 gpc1575 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1163_5 gpc1576 (
      {stage5_13[1], stage5_13[2], 1'b0},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc615_5 gpc1577 (
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage5_16[1]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc135_4 gpc1578 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[1]}
   );
   gpc1163_5 gpc1579 (
      {stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], 1'b0},
      {stage5_22[0]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[0],stage6_22[0],stage6_21[1],stage6_20[1]}
   );
   gpc1163_5 gpc1580 (
      {stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_25[0]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[1],stage6_23[1]}
   );
   gpc1343_5 gpc1581 (
      {stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[1]}
   );
   gpc2135_5 gpc1582 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage5_30[0], stage5_30[1], stage5_30[2]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc1583 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], 1'b0},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1]}
   );
   gpc1415_5 gpc1584 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {1'b0},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3]},
      {stage5_37[0]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[1]}
   );
   gpc1_1 gpc1585 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc1586 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc1587 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1588 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1589 (
      {stage5_3[3]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1590 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1591 (
      {stage5_6[1]},
      {stage6_6[1]}
   );
   gpc1_1 gpc1592 (
      {stage5_7[6]},
      {stage6_7[1]}
   );
   gpc1_1 gpc1593 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc1594 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc1595 (
      {stage5_25[1]},
      {stage6_25[1]}
   );
   gpc1_1 gpc1596 (
      {stage5_28[3]},
      {stage6_28[1]}
   );
   gpc1_1 gpc1597 (
      {stage5_31[1]},
      {stage6_31[1]}
   );
   gpc1_1 gpc1598 (
      {stage5_32[2]},
      {stage6_32[1]}
   );
   gpc1_1 gpc1599 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor_CLA162_32 compressor_CLA162_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h6fb9645655650f464a6acc231c3bd81367467361d5e65f3cb2e6dcb99e02d803ce463cdcb059a52d76528d126eeb8c0403fafa7c7725e5748f2c5b856539abdf88cbf6836738cd346a8c80ae1c587ba5bb99009f632c830643ef825eea6bc99ba4f48e8cd099dd982478c4b566c74b8dd4437528cadfb996d44400af9dc2bc559cce51e9793cdb61386854e371cf6bc131d094bd75cfca05464f426775b90049381b7b7c958428177599d84e7affeb314829c43a3e667abb3d4f754ee81f92d16ff8d52bc6e43a53867960449dddb0fab132722a33fe901c0f8191a76eec364c237aeb797d34cb1022146ee9641840d7451477f5327dd438256aa5d6a169c4a240e048bee9bc073f86d7c8e304f812852759f31890e4c4c8de6d6a1ec0256a8474030f31da88df3b21e97d14f551a70ddc76c2219eaa35797834cf630e4e18ab28b11ae84a55baa4a4606b64f6a4ca9a85bdd2524f55ca7540aeef622e4c375e620d9f58737c3d62210d607bb3754bf547c46561c6c59f20ba6f748481c65c9dde462cc59b93dd4d81c6578e337a8eb228c20b777ba10815597cf0d55b93e1661789e73e19690883566f3db2956df0ad53fb17448631700f37ab511baf37732399035918ee4bdc12146da02d279c5d986980cb6c82c6f6d9da76ae470ead2d7a3473170e3e9df1b72004c09adc9f23b754c764672565c96375e181ef50edb37a4b8eea5e88043388bbf7e2f49e856f315672d44efa65f81577e08bda84c40c43396f0aa78d6b6d84f5934e2a557ac1ed97afec30dd3b8f9ca8dd430c5f84878e295b9f0124ebd661a03566011d941972c5de72b4ff5003275ecee26e683d4bfca020710e9cb8593517f34c93a933b9a3b3a8eb75f4e8f3ff113cd445e666e6bbdbd1b92d3e0362f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha01cda59555b8c4863314120aa81abc9121a1168122b9f3293750130a2c4429eb059e81c63c6f94de36568f797c424b4129a748679ba56058a70f0153c193ed2e7730ee659170aa13c377be5cfe667ebdd7919d960e8939245ada62f96faf5e5f21422fb731160669be6e3677db3b2d98f1b7605580770472fe2c7212c8362fe9d07223481b6f67ef55c057ed86ae75d1f5f42867bb6c7ab9177f1bc7e42317c4515a5ced3fdf4da7f51db88a2a3b750b511afd669942ad1d1d80614f4ac1a5f1fe242989fa4fa7aa8d558d130cf5a84045c84c49cb2bdd833a2f739ac5b2aa153f3373ea869830b958e14f65507dcbb96320950f7564bb05564c9f50cb9db34d99a34e2e31da29389438c908ef51beb7bfa4fd45ee43ba21786ead2410f415674db8065cda2efdda8980dfc0d3144ea021f50e1574bb6ed9b86639c5157f311a8b17e4976bd298befa29c9e6338ba7843e14b544fe23a1ad86c571cf0e3f36a071ec3adfb51ca60a9c12d2d5b82c19feb02b5b752ed0d1e1c9405502294d96376ce9ebc466f198b61c401f29b2521d97f426c24ada3cd502c6e0a6e81037e148deba9f3c53b849df2d632ca9d9ed4a5c000832a238974b8f28797811e0c55bb599e0cb26f16681e9550b42910123ed8678f35175084ff81d0f9b0913513b4cc91f1a13b78f54bf1796cceed77dc292993c5e81950f56d5ecf1646e73a559e80daa3c54f2b4dd9ee846dfa896ed7237a944351f17be3e1b5cc5eb258a7b2a0f0420dd25ef627d511e1f628f7369b4f959b99fc5faf512d38e647dfba91d92af8cbc359bcb4b5a0daba8dc04b1e8a4968c3c903e408aa26ebc4ed984631ab3f0ca389d40510fb2a64cf0841bdba25aacbce2c11da6e8fc1ad66d5ae396edf71a1345b121302414845;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h94fd7bfb2a6448a7fdd8d799481133d36d9bdc709de3659b948ac290703cdb1eb6db040e9e331caf0300afdd5ed46909930a1ee8ea031bf19922cdc2d26e72b07dd002539267927992ae2df45bcf3ebc688948b872c407fc9f1176e84eb6c6cd8eba7aacbf57b9ce68f1bf5309e7eb067bd9eb4d57eb981b1e72eeb12fc35cbe84310ff60d27d83e11ccadd96af559d4f7ce2dc0b9d1db488d5c00c9497921af3dcd9d44d8f9f1e61512ecb6b91212847cd51dca8af0ff25788b091181cd7094025613ee52abd2da74547c15292e499c5420ee2e2ed576487a7d5a8cf38d4170aed6d50281a08666bd8d9f4b159f29f4f2ee75151fe5cfbea9508785c86f4aa9f7b849104447fd6b7ed65586c490cffad97168b48130333ec8c536bd12e0c0dd9d346156d08d792d35cb79dfe7e089127c7e3ae6c499cbaaf7faa43e2261a5003ddfc84d3bf475f17717326c0c9d05a0b4f7a7bd5506bfa9cdbd0cdee218a13604e7c94ab1cb06acec080389c2ff89eac09912439a679cf7eb8a7b107fe718001f2490afa4ab1e3ac991efb2ade7a5898b51259f032e9ffa5c5e8fda7f39855e8282223ac49980e017bafae0ad02035779690f414f61c7bdf9391796d00127e57aac92b20c53658ce230d6af199234f395e0e4b81ac6044cfc632b705ef4067254df77cb94b87f4682340cb453ee3ea4dda28e07142c7a13e72c4e7142055485bcd1f17d3352847c9e2d0b7bd3b7b72a88f65105c1f865d80c237dad550af12fd61a9f9e6afddfb0925a31dfcf26c0ff3eba8a0f17ccfdc0bce9cccf55be9803180b3c94e9a99db1afe3a8e30ae9efdb65d8711d681c08b3ab05ea1e7b15d3f446ad6f6fa141f4bbb8f45f3263b16216965b13ab07e89c4a59c3a4d2e5f6592cdba3c2374adc7048;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9fe9c6ad18a057d2c9f62b0d7c6160198a531cbd3846c53a8db86b2d208614c71896c6de710975d1d74279619811888125e085a293a209a36678589c57faa37317cfff5958a293df952b28afd48625b41b7b19f01b0f4a93c9c2d560c8c922d5618eae93b17e27b746f0d45ad11ebd04c84c29c6f735d76a7b9a5689b7981c0266ee85cc06765f512af5ad3da4ebcd487117e7652e52bdd691dcbd2849123cace7ab81611eb19a0d1629d2eff7a1c8907cd7d75ce981edd0c99fab9f43513c37b9543870404009a61f970dc2fb2cc89eb20a5454bb1e19dfe116e3cf46ef159949ccf2f91c823439180e3176bae215010acdf40abaf971eab4ecdfb5aa3a5476e7e3d64000290dab7333736f3401dd65dbf8ec0ae3907a2a648091a2e56fb43b8a803fc4174d82fb567c7de2e7b4a4a38f65077268521f5926ac706c01320b84002b340227c1c5faf4c8045ab51f1273860aa4fc9ef497e49fab3ee479ac0d7f4568d01afb0f3a654ddcdc9eef4c427798152c5430c4a46f8fdc98425e76e6dadfa68c0e90cd3d552dd3f17356b65ed52f3d157b601d1686b297d1854e5f9196ac24f4ce2714a70dd1f4e15e09bea5918755ce437254ce278880d0f1385c0518f0fad826de32f7ecf7187747ed2618173eec530b26b344172589a8e2cac495361e087223ffed71ce0dd25452c846524336faeacf9cc97a138abdb5050ea012cd97f3165d0a49e399d792b325ee94a176487ecf89fe7ff6df822be11e3c2adc9fa665070ca71570994867073cc2c606f91c0bc410b0532c815c3f40f37978cbb91e92bbcb44dafb63fc9508d90b862d4a572ceebdf41b83af0b748d47a806cd00d2492c23911405eb13a5c9616db2aa7c7d504bd6b435ebf3727bc856eb06d22ae8b2d974dbcad396;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hff35e1120bc8db945a208d05049c010e29f3f84d54860f7f17c5b92639fe39693343ca61a74ddd75d70eb9183f3edcf3d321df17a9fd38d7c392406157cf1c1b6bf552425dd51b4c98c82da0e9a486f04a54465dca865059c736d8e2258723bb98135d8204bfb50258f5e25fb55be5d8bc3be990ad649cccd5d78e8b5087a306b8a810a6b5371261b2bcd6131dc69e9df9684b703dfa405162d1334b89d7c5a739a96e89e6e88179cc7b09dd82bdae91419e298ea0849cbcf2d16bad2b123641f38ffd673a7e80c09cc0733f6cf94b8adaeb4c860afb4354be1e8c5d1c1709549fc2efe08f5ac75427bb16c721a2b97a2c2052547c39b5f71154f2cc3cf38d853b366d417ab47f4be4f0f5018f340f5ad3da3e23678fd8d307a2270c99e989e57b5eb8cde8baf1a95e5fee551fb0592390c24e36946fb7cbb24592ade30e12fd948f829f73043ebbdd5d49a517ffa3f7147f395d1b817892b619bb2ddb47c39a7a9a606d1cfba803f99c75a15e56aad321cb42e094ef526eff01f6638c9392c7d2c52ea4e79c218ec91099699060d674933416cd773e2aeae0e53e006e47989254a320494c2065ce28340908dad7feea172813918d5e7981064a62a9357a7fb52152fc7da4957f491a07f75930521e70033c76e1c885a7768e3611b7d3fc320bdbfddb1d79c2c9d1631c73ea0418a022e8b599d731faf745bf241e7e68618eeb08b8650156414f715cae30182df4b9f4e1a47c00d9b8f6e78160ce27628bd854ae6ffde527f2e12f1ebeb9a5fe40d5859bcb0833b476a353954bee6cb6d3474748dd42113fa2675b8be1f34d0b7454286dc3225138ac4321c3a95f56285194b42d7e20b0a3fa26c7c5d2456a89c36bda4495df71bad42133ba4f28716cd08d8a32ceceebec5271b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4a0312577b0fe11a3dcc470b582bb9da276f79eabfe1dad3ec7f176be4fe133029a8d5839559242e09a543609e20fe6ab4c7e27a4aa6dbc07e7c781fbca2f405cb5860c57ea0b70a7e20ef18df05677ce6445c94ac37d482a0a908df073a0314deabb8b0ed8c90369198800fd7da71464c46326012941f5fe343787cd520515dd62242206bffa4a8b09b26d7c56cddc87782e67e16fd055669830187a13bdf9326504d175ffd5129882b3dfab268588841863e99bbb4766ff672e9d5d556108339e201918142e0bff4fe347a73ad842d47ad3b28845773b4fad49a5eecca3a89e63c9abe96bf082f9ec6ee3fcd77e055dc1b55932873db94508cbf14f74a483c4c6c6d57f06ab0132119c71fe240ede022a1b7fe217a1252a9b70d406c89f9b341a875e891b9fc3d0fd65dec7e732171829840ddeb801b57445825687790f7657bd83d026a5fb144de279646c9a4987de39c199471adb00050341e305d33d466aa3b991cfa5c13c0fff849920cedd88eae28d81a3a3ff4027f71145d977c814861f3538f08e8fdcbd5a693852cccf13db535643476fa6bee23b0c1bed1f4b870e220ecb91366fd29f0d69c8c934f6e9f068c1fdb658413eb284e378476dc9f5646fc9566cd3c63d2a96625ec90b08fc54f2d25158e5c57c7732bdb057086f5e1b3b4a38bd5bce804879cf492584e49d035e2cabacb6ed77ae6a730e2dec4606599a30b47b69e2132f8fdf0c74f4cf25e65ff28d0ea8a5826f4ba5775ab3c3e597fc2759a9cb4af67f41f6c0b0addf2e581ab98d79ade3cb1a0d6b060894adfc5f53fc291e8ef08b9051930756afe1244a45b8c646f1ea283bd7702ee1bf93bf3468509560961d2efb4483808d797a77e1495db76d58ea2258f699cbdc42a9bb30e79d16d54e290cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb8914549ddb21792d4e2bae1a5b0dc07e3da9364ef8938beef8d4174c3ab7aa25ca3fb3d9ebb4fab9cd9286c446b3e8869d1b6e0c531bd4462db5e427174f74f03ae51c0aebeca6e9210ba3e2f787bf958df76c32e36d94e362c55dc4c914d377ae4fa7f0a5f2ce1e6028c5504a3bd0d81414327fe39ff15711fc8a9db6d104a03db926339c3aba7607db06dc6f858c60421b4effcfe0a8b4e7304bba827947f49ba6b8ed3f8b4783ab28399f040a640fa1f22ebbf30d9dfd94b86d3e43ed2f6833cbdee989aa0bdc15033a9bf58837989554a4e770ea9d004b360ae439c969025ac235157fdd9417609da3598a3c969ba1d24e46b115a272f85d7c88dd6cd40a3888ab6d7811da2cef039abd602ba0c2f86f2f1cf1e3033f1818a7f7f7bc6016840c2486667d7160e1565b4a85a1ae5540bf3c2f9a044b5e2f095dca2fce254a0841b141acb48a0a34082aebde0a4c489d27f9ddaa4be1ddf6a2f96c5eac2a97b93fb3457d1b10ca1eb7244b8983ce5eaf27e40788645b0cfa7203f5dfcce03d09d0ac6cb48e1ade8583e5269117e52351a6c2f2f10c147993ad743b5c9817499cf19365f3a74662d4e52baa4124e87297a7ec24038cb0389ba1d09bca1a4d70639cf34129c7c1863e4afb89ad96ceba173cc74c83327754dec3d5c39b054dd1b2d79dfa6b5b830883f617af54aa2d22556ab63b417581661ff89fcebdb120dface89bc20eaeacc8d9315388d4437205f6048cf7645fc0ac7fcba08fa18c7491e60fc472ef157590b5db0d3220c21280e17f45d477dad6ac7c93dd047afcf5aabe2365503b503b5dc6e2d99eba15088f7f63a5891ca5fa770c3dbe51b029b59dd3f940e4705bad2bf333dee2ba5dfc4036989e14700dc9727334a816f522a6179e843127ceb6a0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4ec647620cd690addd439c60f40cbb5db4dcc719a90e57e7553f8f28bba222485a8777d8807e07526cba72e6d3482d09c24f8b796bfc2dfd8df7a5a1a121ad46fdafeeb83e23d1b76a67460152f2c4ee1c2513c78ac24826c42e67dfe5ecddfd42de8a38932813ac8b55856f590f530d4bf89be5b341f1a3a3198954b262bb0647012982829ad1e19024db8a58244cc73b6addd8a781148a546c14339834362cf56806a49bead27153c047beff9ed80c03e6f7d0edc964c2baeaf4183dac8316a94922ea61f004134adee7d52996913a92d6232e04298c751d644e2e2a8a464b4b59a34e50d72cb1aa3d5d84cecbaa4a0e11d51dc3d998a8da651801dc7ff2c21f8371b08515d25dee931862e44519ef3f0b59d7f6a137cd9aa75ff6f4afe0a04c52a7b78e51de4f072c7e6b748a093d1432afb7708e88cb98a867ebc618dd250b1282cc7409a19a4cf0fec98a355c9bc95e9d60941e30b4a922602e9d7cafe996f58dfa2455ed29deba39c9caf98cae2334f675a54cc3ae25499833a0f3f96c1eee265b843628622e15d94fbc446be3e7e2ec0ee0c930e3b60a00009f28525dd013b16ec71a92e58a0635d2915d1ab496f6edf1c70852621582abdbb60b0031955b2c1d0adefd738cd826d1aea352dd77d755210346f66b5c9ed1225aa58122d85f444e75a38dbe228a7ffee47e18597233b0386f05572df5c9a2efc794edad252cb557128b08b0d813eaf417e2720dbe9d387fbdd614160752bd1d4e512f267ac29f22baacfff98b97b956b37a0e359f092b3dab57248514ebb2644e0345767ff53113963feea85e9b073e91780b58045b836d887eea986eeca161cd2199e027d3c2c666826b43652470e73f2dd19481bab23ad4030de02ddc3275a3fa2ca8883986228d04fb36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h10e6e434f0d05d4be788df468d164da81ab6caa5b3e230b2d3af0f998c4a6a93b9d8ea70a80632992f3f43befeb50d3c31cd4e0b18a38f5b74c1930b5934f470e85972af81a6ecaddf7cfac4fb858bb9624c0f89ecd2179c02d772936987048f67ee0356fb5ed4f33b2476d88b7a3e527da7fe9d2e3fb4a99a1b7b35021fc25029a1c9ec9829e715506c977650fe42386f704a7658a9a46cbff714a123fcfbd60c920ce5f925c4c3c280266164af02cb67150be90e4c5c17280fd97a736308f0b7fefbc13bc361cf699b3614174920018907bbcaa1f45b3cd792e9fbab68172c2b6b356ed0ca9bce6efbf775bb30d9c8cc38fc1fc77159e77b3045adfc8fd6b65bb7f2975007c9ccb1354209671f189bb0b6ca05642781eb12aec6c1628b09a6470b62379c85f828360fb3dbdfd57f96c43412af3b1825413381c84cd60f0c010d3c2cf15eb8ebc9ffa6d5934abc0822a549937ceb2fea8a1c3fbafd88cc6c2d92e79032773823085e166a12f3ce8027b57b52e28a2e3661906c8db74d97a27d493d4abea7db7306f79169dc5e44e2cc9bc18d8e155eb4996ec4562104da42c83508c80c72dbd85bdd2deb358dd79fe485a48ee6d72d3071bf3bcaec780c2b56b84d074b1a4dc019864ca4d4a99de531495237a4fbd1cd63c06312f4807a650cae6418ee8fa7394878e79a4626fab3654e913e28faed62851ce4542df4a78a2d99c5c9ff28b008dda2f11dd8ca2d7e5c3151601d6c7f199a08efe70d677922bdd707937df7429bb4c030fe752664914876a982752928c3701300371012cdc8256350f1a5f74e222c8b69de5697bf97c8489c91c07c8db530ac9146313d30adce1894f94a8bdea8af7da7a1f60f9f4ee23d4b8ccebab77a6cc7be61dc9556ae21e6799bfea058b1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h983f1549a337681565c9bb1de7b3c2fbf1c6f7d65d0297544646df147a03755fcd02521f36d023c74fa04f775c9cc9f955dd9db99c5186fe8ab1092beac8818629db6331b7ff711c4640b0d48637513f75b8f85195960477206b1b804542c8744fe8cbb19dcaff67fcbb6b41e2c4b22f1b75d339093ebd15ddf464d446cda9c09a8b7368e147661a2e8d878a62d6fb9abea2e56a46b0d0ebfef7b788f897a17420058ccaf0194fd758bf9f72013ce9f0e35e0e9762487b58a4054177464c43ce6ef13b91c81902bcf8b88802e31cac6db21bf71e818f30eb2cb1d2e47b423fb5b81fd0132b38008d331acf49eb183262d4e51a6b7dfbd7ac26054c09297c376d8e3560c6626253f8e13a6ed309bbc78c546844f660e0672a0765de9e62648690a00a979ec958aeddcfe3a10c7889408b19b47aac1a229fb81127d915938213dcadedd4f23d96f3fb23de8889261f1bdf7de12e10e89718a11b8c1180b4ef9bb79cd174d21702eebea8153aeabc34a3ff6d60209557046b6bc94f02233cae5e0ada12f95de735d19a31fc3a5c1bbeb252dc7d0053c50381c76df0180c307c10bd8b6781aa138c362ef23afe50ab113e39d1c54f3cda01b14f05b594b46300368b0bc154733d8f93159f6d88dc3ca3468269672fb0eed38b47330b045690a77d39507b2a5e22890238828761cd869545c1a734dd28033cebf07d1a393f1b060c513ac18dc346324739bef54c458d2baa55bdddbee6af117092803b458806d70f057e5410c686bd5778918381c90e413ae7db9ba9fc1256c5a1707f5a08e319ada4c306124e1d6bd36843af7e09f8001c4c0ae5d8fd75c3283d93577cff9b6e4efa201e60c809af8881046fe83a679fc4a612fc1cfd7906b2415d9462d5d36c1e5d4c1d3161a2365459;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1facb63fdcb31a85fbeb4f8b4a1753ad669e05f357e83466a57dcfcc6ed8dc6149dc5b09afd21f5a949cb8989207ccd606b8577aabf34027548d7d509e7768a6bc41198269d13580ef12284b9757c95911a74787b7bf7064c146ce877d83bee5ec26c7d63e2603918f6bb233ccee627163d923b46e7ca372170b90d073ba90914756a5ba3cf9416e773897d1824268492497cf6e00f9e0b007205f755537b2ea5d412f60be793d12823ac4039bb5895c8472ffdce5c5ca6196b0d2a5f74c79b5f6ebdd8112509f31200145fe474bb628c82383815eb43c54c5f9c6372d575cbf0d7fdb1f0a2e939ce461da63889ce16ad5a12c27f40d5162fb9fff0e2a9e8f519a58b0d1df0e69d31643172dede6ead14e90c1cec3a32fc4fd154049220cb1f4f36fbf0eb927df8c836f090db8e9b9ce7f8c239b1764fc847133ccbfdd87c87c3d516efa268c70401f42232955e6a4d39ba8bc6f76099434ca8fe620121e9fefdbf120f3b50b4110ce65c10f85010b3bd9253ff817b870697c314b2f3689ef83924088fa69aa124feaa2a5399c1f747e825d1f62004c84e4d8f1c2a073006a4681e26eb8e54bb1fe9c20a8e6aa3384348ae26acfb03e7a1b34f4b5b50112b48fa5706186b906376154ae64da407e73549448e9e074b4f6c17ea0b50e92c3e40994a6a4b657c1c409a362b3f4d97202ff918eccb6eff02ae3285ecb3786348ee3721852deba2ae9eb39d5195d56ad16ba7f3d234852779cea7666dd1b32d1a1bd6b683a8cde3e09904231dfc8e0291b7263099c5ad89cfb6b26b601f4f35290eefc3768637f9c121e0b415879ba2b6f90a34061aeb8b076e42bcadc08e29e8d66661ecb6bcaf8b2697efe0e16ef7d84a5307244c3556712769d5ddbdc51b7f5be5c5d7173f6e185ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfe018404400475486a5e63bd879732e93ca0b56bdc17158e615059c3148221f1882bc50a39eb81b893287fd3e3f78490d16f7ee61c385255d6f90679c61d6f4124baf766961472cf3e46965ca21add35557c724b28d6a9145de49e8fb29d1d38081864e20a22c3b7cfd8a6c4c2526bc934d6aad07186dd317586d67551c623e08b1e5271f8e4df1015206cd6a6c3a2894dc86e9525a7dea94be76ba924b2090d8c966a2190b4ddf8b830a7de7d9ebf9b312ae57706b29ece4ac106191dfc337000d84a958f646c4e7bbe61979bba65397a2925fd11196fdb97389769450991e47537f6cee496cffe6fdd5fc0f40d7e7527afa16dedd9a8e0446fb0b764626866f1fb494b7c0b94279d01d7f4f10ca3584142f6df68805897119004721e6cdc4de0a9ec8ae038a212dda7c6db3fb7093d599fd526f4fb07c280cc0732d1ba0de6b4212da631c29d150c98b1ec0662f27c5cd54f1e3baf93302ea1ae58010b9cd018eb3d5cdd16a91dd4a5548690b0528637393b3029692733c71aff48c08513edb460d2c7871bcb5edbffafaf76b51e622c32e8c6ad6e866a50a88818dc52c8cbce686b5b7cedb949f31533b221de0ea33547a9a9934978ee45ee57df4adf026f6ed2e6aa192a25d386b55cd3a3c9f8d9cbb84051f304e1775e7c1f0467816c86d53e7f642469f9ab4200dcbac05c769bc2c8c9c50ad2d7157a1e13c399d0a18306f850bd0dcc99b8e4264db04597183b939b894766f6fd5f8935e16d8d204a71a59ab4c0463084cb1bc45d449fccce44a8493e506d15fea0274d1b624150cdb210ba7287b3af4dd6e58f5ad97abe2438bfe71d0f78946cadd1a95ce90a74f7ccddedd0255e5780d369b9d9c07e8970404d2c4d9544ef77d85dbae12e05143fc8aaf83d8a00fdc60f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5fcd8265750b75c9fa87242150c21c0fe0f29ef291ed84b773fb2c61af23de78b70febeffe15bec3ea6a078e230b8fa3f92900fedde0b495e2be4ebc58f7b6b2466ecf46beafcbd44ef6f070b32f997e2ddb3458949d08370aaeff19321a5d447899016051ad1f1e6d34a9e2d9ff8c5691f3a95f1f8f388cf8b232ace41f793fac8ad1a92000ec39f90ce00562d4f00728d5d85276e2b94fc39dcaddd64e346608d6f0759b7307e597a8516c1a9cbd1f87dd2df73d748d52f598c23b3890844776002116d0f9d595bb4a6c3764f5bbb5317949d0e5e80ea224c8a8d59bb738c4c52d162a5acb6dc9eb676aa9c1be2ac3c267c9931a5561aee21870c0b93b88d9e7ebcdad89ae092fb96171c74e5b58fc551ae8896e48649200a72749819eb08510139b5c33a288813eba036ed0d7717506412b8b194634c68de89ce8e555fcfd22be044cc57bab35c8f19646241a7969d1de12922f92e9d42f307475655ffbeaa138924745c33748b95f565105c03ddb0432a2b415c979c402a332809fc8cf1ec02aeebf9ec94651339adbf7f24db5e374ee16520338ca1f78faf53e9b12f491b5b60fd748d4303218f0c96acd27265e7132b06cb8268eba8f58d6cd1804907cb743d08736a9b867daa0535a6d20904f6e5c98ba7ef0f52a2a44563ed69bf4bb86437cc23940130daed5df960cc0ccac172323e43206665a92bab72247a8463c451eaf706c63d617d235e939b4642279f0ee55a75371471f8d851a7bd2423d1b339a825834bc8749cbfcd0fc040b9b6d0dd95c477df17393ec6a9edce72e2f90df44d66d062e14238d159e54a35bb7ab9d646113628c959d369c4ce476fcce9d0a0bc2670d1bb033ca7bed58c546f59c59f2fd50da070034d274cf903f332443c5d748bc3db21273;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h887ea628cf2a61d5d708edbecc1ea4c497e32819f1e44432adb0030ddaae190956875c3cb968066d026505bdd7a4c451d0628db8ff384c1cf61a6fb6bbe768eaf755b106dec8b8fb3399d24ea4a4a96acba1095013704c38ee1ca0f3b05cf0b1972601793bf0f3a36be1deddab63ec3c5c6f44dad4cd69164bde709f3c0a6b6e7b40195a5b9ceade50f26d30628d8788c414e0d7091a51e71d97b78e0096af283d6c2e1cfc35dbd1ef7e580ee9c8b2e305db923f7d4537e84abeaaba167a5b19e59c45bf3d73c709eb4281a7f8fd74551a05e182dbd628a85957b787977bd29020f2590d1c8e6ce9ed6a1e0940805fc8a215fd8cc97e51bacc2d839a25f64f39040d9f0c719539d49d8cb604d5e783d99f32bd5ed23507b7a75a197cd5df7e86ec7b129c7e23efb8986628481414a45c809bd1955fb516e5cd1a96a83b989b090740f1c712e0d3a44571a885c333c3f1b61db3927fe287e25204b8d97c36b598dffd322a453505dcca7095c70fa3e0546a5415004e29d2ec350ae8f1e0a078014d3faf56a7d4dd330348ea495415f1b8f3b96fa90572edebb8fb080054844cce78ac872d6a46a3450f56bd50a865c6c19ce1e667b42a5e7dca009a82ffbbc6cfe828e126746c367326f2ef4d60f2e85ecb7d4603274753f5f1b0cb701669ad0ef13dfa6c81d3731d7d87586d5251e1fd7e9431bf52d3d9d870ed550aef269117633ef5172b4fd48643e60024a67dcb7bb4750b26a8fa1ad27dc300fa03a3b95b9a91cf20848c638df80ea074b5cf8b754b36203063e7af8cbcead3017b76c7d9f86cbee188dcaa12ce80b4371e85b906d0447f793a4c62df7d0c9ba5e1c8661e463734d7bcb40487ee89d0a5c8262d725f7675a03bf6f7c4e19fef6ff910b4d807c7d50d39544fd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3a0647acf471681fb30252aea9317fe314f0a6291134adacad812cec7581401f3b727707b7090e27dc956e048c9517c06c67b826d6a3a604feacdae23325f087d3fa6b22e8d46d837d29d5665eb174300093813384d2328a573b4a4e6f594b3c752ab1d53efab4408f06c81c1209ee44a65216e1c29a5e8b3fea8b858f51cebd8f1e6348167493bcc9a739945892ba5ff4332dda0e4c0532ae909cb95e3615e83f06f87e0fe5087734387e74bc61094046c4d42088822b793925bcfdd6ce397dcc327fba9842db6f7e2dfebb896bc0614407e8f588d7737b73791338fcbac72df8e7d807444739601193a51f3bb2ddc5da0fb48536d368140356c2f135440c6574857d69f64c333582cdaa9ce052fe24ca689c52d1beb8ea49eef12d3e89789b6ac1c2e89560e1f672cde203f92492a1180c490fc590bdda535185b300fd3440c606403fa30163a21f48efa9163f67521c05eb3d475d4322ce38a35c21703741315b0d5af275ab328fef17a11ceef8aadf2e833d0aee3469795458b6d5d755e60c382ac70d95b88bcc5052168ac2eef87c86002487e2cf4ee2c0523401919d54dcca2397b0f7ddb1c2b27b371f607bca684b84fc7220ec81a9acee29bf1205b30bcac543858ae77cee52e6d9676a6640ce68fde74458c6afae3a1c571d053bef7303788ed102ada9fb98b46d3342e37493e344d55ebf32738e011a9918c8580fca51f9f0624e6eec7f51c0cbe21f7869c12fcd4270c875de205eaa3bf954a3893224e2a7b3d2d5763e7857696d9046cbc1dcd2f05a534f072086c3aebf551a5bab3dbe9b65b566a1d5ab2b8942d60bf33a1c219d4e1a1ccb17d546ed17c3b92fe1a1f9fb7c4003409ade64cfd009863e1abe629de1aa598845060cba5e22b3b6a91a2a7ad5c8e7a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb456783b7498aa7ad20d89aa14f94869be726944d394bde18f3acdf6ce7b6f59ba20d8cba22ee5f6c5a2e1e75f5fdb922856b363a6bf49820b4c962900bfb914259ce02de28722f2cd88ee7923563612a4f6b32dff9e370660ec347dd3db54ed0134464089eebff810431e8bd055ade23d6713906bac0f98c115187de531af42dc09ada86ea9a44fd1da8b57cd07c1356113c976d6e0a821619932df41c62261321067f9a86abae0543eb9c5391482c286539ff1162745fe789fd0adbe2020ad617ce85c01ace9595736a91102e96e3152bf4cd6a2c2cf5f58077e7ec46e3fa0aac927526c7fa48078ecd729126a5f839f33c87bb554eb52c3e8e8bd201b8bdfba2d676e8af2e1d64e6428146b93e30c6074031388d4a1a0be1e2c442e1cf3221782326debb732002f36258dfe06a97c00545e81bb48e76ab1237f445c297a5abaaf2781b5ad310a2788b1338348db137a3118569d95cd71f1b0d8b5c8d6a94f60bbe30417a92af040792245799ffbe796c34675ea92927aa8c8d4318929ea669661749162a23b7e88df5a836d4407dc68c3efcb3134f71a473710c9976423fbf0bfcdfb4817dbced5e02ceb980dca9a5b68f7b402754b92013144f1569838196a69cefd02618f4ddc27bec888d8dbe1c2e18c82129ab8a1faf53f68b8b6e36c639b1574fab0a02dcaeec7a4cc5aa2119eccd6452ad2655e98966c413a039d56f043b2cd7aad0d09ad5f381552355fda3751069512fcc1911be6c77affd69ef6f900112c1fa1c5798e0ccf68afbf7fdc0bd98d1a31b910256c89fcdb9efc2a53910322d129292edbec584aedfd150f1acd5a17701d2a5d70e76265ac52a0c05e588eb4accb057ae5486d555b99ccbb65cabe7b2809ed99062aeceec6d74f12d3b277b622f202ec2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5ca164c14a7a94a46a27b4c6172b21bcd0845dd4b74da98c492015b56c5a4549bf869ff834bf2840195c54ead4c41bd7d5516dcb92deeed5f21b123ec61c7bf167efbe6b8b5a0881e65f476ba268ae0e72168e1c9258bdff5a86fe06401c4ee824cc599db93661195917f3601415a045e599a02bfdbdbd0465576201153ca98a17ea7a6ff0b31e525f8927f0c26326918dc623e69ae9c52d1c9c55f7bcd8bde57544a37a2a371b47d26e1006d62cf9a9d0dde57aa4282a2b59b03c8d7b647b585d3949a6f5e01b7ba19b0c0a17c9999bd885c857c0f91f6164d53520efaabe2c745dffbcb225081f356324a98d8eed853b3d9f06adfcf2eb95885d93bb8474c28e23a8ab524b8d0b960f009ec56d82e8624b8864483c8e50527899c52633e717f9e999426e9e76a08b9ab3c62f3e30f107e23be43acf4d997f0b02b511287f5dcaa68f27479283f2f766176105cbb6c7d082bb0187f910ddd20b8e3720ddb91db79075d1c8b045b3ce5f3a114fd5c5416a193fddc3b2c6a1e44b87ab63866e70073fb82c2aae7c1496cac4d978c9212e32c569b1be430c48373f3de90a7c443ed2e0424272f997cfd0590f525ed881033b01050e831921da6524212df382bddbb6b1efb19020dd8801950baee4014dad839daa46909ef5545791ac305e7a57c0632a95614d8098449e855fc04a3007ccc76659c19e044ec5325aa201eebb9942ff7a7561b50718ae6af944688583019426fe767fe33e8355251bd82e508bcb8b854d46091dc2e9ae78244b6143b021f222b2ba09c8e4f8bd94826f4a801996c36973bf55b9006d3d44ae0719b2679a676b3ec46da89b15e97aae223a2e11f7083173c2fe5d7222241b5e6ab3a695024a240e7d49f8fa9150879739b9d0405fba8c93b80a436c46e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc831022852242be49aab2702c3759d808d18a352cab33ed7b7e2423309957963f2ec0c9e7a6898af325f6d9d42e752a8518df57e949e9516d524659d6132bbae8e06c49256830af84cd98ef7e96b4c185393aa26d4f8a5d2e575d1b643d1dd0808ffffde94afc30fbe401513e8d665cf233e333dc2caed36af568adb644cb189a0cd9a3558aad4f1806ac035c0881cfcec6300146296d06e246a7d456a7b1cfd875ec9d7ee6e8e926f8c627ce3ad4f7c8d3d1182b5060e86f91c813032a6c3cf0e3463629d6c6ebc9fe2c584420519127d4b0e4fdde88a46e5b1e6a7d17d74af20dc3bed8b4ae6e36082ca16aa92d9a7874fc5c0abe0bbe5994c749ff8b6e0b1015010213ffabe71fee31663154bf799ee32866220d5a6823970f56e0d33d17a2e594042f0f87e6b8836756181672b16086255fba65eaf1a852366b54dcc63ffc8ea089a3aed3b11ceec5b918044b8aa83c8babb0b0aaeb0e0adffb091946ad689685a1b7e7cc58e1514f0e70d43919ded585d7bf4c280886c7a3f7b527486d4fbce2f2d4fccb9c190a4377658dd416a5ee3c0ddde99e3e30d363189098671458596595af9c2c9e26bd1c1f31deeb98bfad09f159323739eae036828f21fd90255d127dd292ff3dc72dc3405260be2e593396c4ad1dada9b7fe0b4211e8ecd1acf08917645c7a0b6ede1768537fb5837c47c21403567c105020e3a7d4fcc905325f99fee17ae11a0465fcb1a9aea45fa28907cf3f6a05dcc1e4d7593e8fe6867f3af0cb1fc191fccdc367e79ac0433702271ec224c63638f9b7607da8938efa041ceeaedb5f32528a8f21390fbcc59a52b3f147369a23bd191720f4b78f51949eefa289f6ab27825f4b72c1d805d9eb57bdbd019bad9d6e2e161e57d1d024806d581ef0a5a9fcac5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h54cd7f3d40ad3f2384f18f1551916d2162de7191edf55e804c9eaa006504280832b05f6f81b5dd4359c24b82a74a6e3437f5a8ff718b2941fb584eb6faccce56b35cb50f2acf1d54724b640f6a7fb87c05137a475aa20529421b84a3a2aec3a9114999c0490e7982ea711218c3c67ffb74b3468a2f54ce906405a0f48e6ab26d44b24f82f7d763af8acae3cdf9f27647127fa8892687e79ec7dbc434c02e339b09c3450f403f2f372a49b10e14c033b15d03de1fe68c0db4206df29a8f37eb5343d3a8283ed8d456fa28782d3377236bb24e99994fab7414c11f5521b22f228fca7602338f722437fdf6a1eab57a5096dd0855196ed9b57e5680e0bf723c4288be0f7d490d63e360e3f7d87851596e894d8e87d023acb0946c8b895a9a2237c232e4b3ada739ac2f1cd68f45e4869385242dd56d4c8bfef7316cc34d7129fc217a9baa81dae409bd3791306133d3db00f2f8d66add8efae715519bdedb6b3d6c610812087797f7f926b8cd145b4940a0d1502b5e8bfd8dbee7d6836e01213f37d24a918ccd20fbd93eccefe0039e4995e15fd60687244d292abc848d69f826e688962d920327f665512297539a9f5ea1ea730285778df12127eeeb80fba833f70934ddddc6d11d207bbb8e0991754c25123495f42d91d90958743b6e52b182c4943223130be84881a28fea4bafd49fb0b3c68faf73ab80205031a3de56cd8a7b7e740214f92b4b6c4164f7064a4df36697af2891a8e0c6146fd9448c7ac4fcb2800d503fb6e69142decc5455b8bede2cdce0b63905e181e8cae4aea253092c5340c12eff82c3a0526123666a50e58df616d2a8d1ba0d2ebc4d310df2de4965eb96e5d561669f27d742d74bbaa826b20ff787dbcbf90214e632668bf8657eaa49fc6df3026a150a9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h51679df854d331d0e5489fb8019f89bce18f35c336290d4890a66164ec6197b6c750ab486f40dc55621a154c71d3b75988ccd7cf9c438ea757d0ed813de0c509b6b2a09136fce778ed7737de8585446614852f8d7c9829e4792862e04873e353dc953f485a7bd68204aeb4a919aac9e7fc20f17d67e427aa2fd7d798835b2234ba50fd2d0b898f79d34b6e7ca8950472e159ff4da14b75e081bdc017a09031f0aa61a0672953bc7f6c4e391987bf91cad2a5f08875f533bf5abefa3174c68e8c87c680893cc2cc459adec726b495a9e83544d29f1b7c72028b92f58582f3ab55212888616e8930a048f60a5efe014f8b76291b504433800cb1b8ee115f19d1d90a473cf7f59194c48362666b9fbdc9f53e42b91ba5fdb153e0565dabdce2797d1aa6889e20513cc9f1ae1faee447eb6945d77b0e4482b8073821ef2067d29812693a31c18bfb4fd277f0704032f0ff1f2148394fc81f5f558e30736ab8fd18dd43db2c26e8dcd28e621a6e473ca18f484a5bbef223b717313ac5459e3ce97c019d8fd79629d73d1df120ba9e52065b221d7fbcadd812f42e81d6ab0059f6b5da5b386694b4d6f1f095a28957f862c27bec943b7700abef4570bfdc509b1f12c65f7ce903cd1de10fb332b388a8934a098cdef99c8040b4d18410c378152299362c116ab434c0323a4a4a00aa27ddfa52ac4f5efd4ee121716d5c020e3860284e4bc587246064fc1493c390bbfbc3e87cb59780c152b668e90680f167918fb0ea4d58a8f95c2e86b125b977e355438b1ef00eef449b50b5f5477df218ac73ecb3026d9aff7088be62a22ccce2683073b3cfbc931a5ae7e70690b41d844fd8b85a13d24978ee7c06b32c00e94d40793649d018485522d57b825ce57eb7a7bb13663caf9a5ba85284de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h496e4c33c3fbf7a196448c5ccb60ff5b96aedec919e5a81814d8553a411963cf68db380b019dd8156dbcf36b235707f60b5fb88514ebf25d24e4f95db6751db5ac2255904d786b5b8a8415cfb8f3be3009774fc9ff4e46c49d27ed0bea8313624e202814118ed61f51a4ed7085d2a750de675c009c3116db11576d55bffd67a2a13d49a34b732a0b5541b1900c6a3daa0c8edc6644c17e31fa0f2299a33e90d4a90ce4e334380a17c9aa617d5f2f247a97161bedb5665b993178d3eb8dfb64c506c24d9bedb5368fa373e1f9ed33d354d96cac72874d7598b7db987f0d67836642d13c69e5c4ef42ff93d793175e7023cbf7818d1d1143ff286f0862ac53d31a2613c0602c5626f08f697931c0a65c58123101984f376f0bf40d478a6df8f12cb04b7c6b5863954bfc5c1455f34f2c51c7c14227dfc34329ba6d93d16e298c2b5bdae00c450b3a3f07bc5e9bed4fd87136cd67d7407bf4abde3220753d38e402e95c04e3927980e1e750e03b0597991b4ab7dc6314d1c8a0686a9190470ca76cae92132495aa597b351152ee7ddd46a6eea9f96de5126765721570560c95c9b502ee500bafedcea75cad581a43a67bc977abf7a8f0c810982e0a6f7e0fbb54609416b08519492ff9e765e3871eb12ab78d2ef7038249df2f52c6e204652dc851d3d78314ddc50b4b45ad64e20b07288e95247d61e96d534299dfb9f1cc0e8441a78872e49926af50ef89916a5691b7c6ccf70cd2f35cd67726fe7132b222ff6fcdf1f0808b56213967771959bbfbe063205d7305ea9cecfc69378badd383828637993bdb935d6e9280238cf227aa2b975235a8739245289510592724c4a7095d93dc8893ba022f7c1558622709da2e26686dea5a17c339160e073aef8a4e6c89989bec5a0f548137;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h884a6c322e938efa84af7c21ff01732c3a08d9b1f7f3338aef6bf383408498bcf44568cc113a1603461a22c554049ecb2bd6d2684da9ebbfc3c10cc98faa0118d8a76a3d36a3b892ee9e9f6dd74d217e6cab55be1c7ec83ed0fadd00ae51d698717937783bc83d9c0f6c031223d6e03458f393bb99994e45089b57759df42328cc73a9bb408b010152c17a46a06290f7d8f6a2f7db5f1e653bcba06158faf803ae9db244752545f5e13ba1b662dc7b8a242b112221d4205e549cb46f9120f50a6a98cd64db32d55ca254db4d4651ff633235a1a38812f2e6998231d7a3d4c14732692bebf7143dffba40623e7a8cc0948aeb794c609513b64e0e90b804fc2b1b2dbb574af2e42edf8778520a598459e507807b756b9fb971f5f7a3067c231f847df21ec69e6d844b4a3b1b0c89496a602d3c41f5fd92e4fba463f5d694b8ed99f142d21f4f5b693961240b36c6e77259106237402150925d88974ce55adca9aaef793ccce2b355dc3ff98ec986c2971e7d1814392bda5fc69711b58fd3390dc6e225a7a67da59470766ee4bb687a6f5e52aa6307311af83e4fc6e0c006ba340353ddf7ce2224a7e38540b7f54121532d6fef071a09fe6b9f42e6caa552ba5d333876d7cf60858c57e3928649e47638579ad5b7c0addf535a2189dcda7f0fffc202913ed03c585b663d0439f74057f1033493cd1bbf315a35ec324d5406d3f6b19b79aca9bc959d3fe4d79be0e96f8910f2ed4195f722c4effe706567d74301c2bca0d396d376a529eba5954fc17bc58adf34fab293e52904de746cb3002e39bfccae1ce68c12430b8856ca56031eb1789cdfca5d4280fa9981602a93e349999439e2fcea2424c7fe86844c064024ffd5927aad7a7838f139512a3a3cd208657b1bd102732e901b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h54d0da6191586a7452fcfb627ae8749b019211d1fdb06509bc7c3ed7a0f671b6c856517614f4e57e313fef661ea29882e3d612b541dc66d25b74e82ac3c94a1ab5b737b6cd1b5055261755886b1d789c1d45d1e555127c8418e464e7babfe23c783d198b649c0e413a19ac7b58df9721939ea0c09d4e30279cd08b6c8cdb695f49602ed5dbad4552179a7dd1808db9ea888d64a83126353951a645325132b9c26bf1f1dfa0b6e77988329336302cef19f4cb8f0e700923e5c0b0efc2cc56eebaf2022d69db1a1a7a4e5c47c2b62d9dfc7896e7b4db21a23f9f139eb5eabb7a2896bb1eba5b0ac4108c53c34e2b58e20cfae2c2ffa3a51f86f4fd429131d81c1ca4be7e66f87308b0afdfd5c0d72b157265fcdc31a630352871526d7526543d7e0ff4da9b892b51e7460e843f1bf8edf731dd1d3cec815fca1806bb4f33dd589fbd57c13511861be8ebe77346199132691b06b070322eaa8c043d262f50beea5f97c401c6aa833c1fd59b0d96b915991d1fa30e0f3e4ae45770370c09e25e2f969108d176f48379e55b91736a8127ece6516345a43deb46d6cd3d96e8cfc4cba3232094ee07f4ac1a34c232dca318c3bec40f23b7cc40dbd9515aa014b3e3ca82e112eb91e341bb21d8cd9a4f5d3715308552dfe8ace72e6643351a78ed398290527cc49b819760118d1d6a14ab6f68653a7bff3f880dee4f7366601dbf6dc0d6fd417d7a2d8c5a953adc5da20d2c6d01b44c714905f717ca635a59bfe1d786e19863604a810cbe425b0e57bc90de2b9edbf16c79991f745142eb129c9887470c071bb909ff66b7e9402193826ac81c9d49598062b8d107f021c1b002bdc58327f8d1bbddcc87fb07dd1a60582585fc1cbc96480763ac996b4c85c60ea57079a76f21b2c0e7700fd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h526321a337fbe16e99625091050f6d1d64e83f9b9f92988826141f28e03ba0c9831c864e749beb5b58f901c79535dd6eaa10cff5d5450991d3cec82eb3e75815e281ceadff4f3fc080f210d231421604952ef540435e73c8c77098df1f8796069c095ac85a07e7dcc35d136a0c680847814c57cdf0c994ea0011312914defa074aa553628f9884cc368a018a45d91ba7c88dda97cf79a36142e2ee99fa8c6ad1396abfb4dccc11037668fc9d6cfca480a20f8da6890c9d2bd541e1f7cb200150eae6e13540be1402958d281624e016b877dac98f79dd35f56159537da7c786604e5d6849e90247308cf355f43d7fe23f9a3066d1472adf96a6020552aeed8c1e2311be27d733dd65e85daaa2bef20f85d14795a85bea58702ed4f5ea1a13e4ec019b5d9322d2ceb1bf8f900742b0743dd1f0893aa827514d2fd6d4591bf65e8b42a79f6d042a542ca3dee16f394e29f000e81ca7e81cf4ce2517d824a557c11d5a396ac3cddf9f8b4d583cf5ac7282ebfbe592bb1ab0a8ad71f9801ca88a0e366cf42dc75d4c2b720e412f812d842307fe3b65a82fc758e10eb625d20b55f92c44ba19ca94520b00273c80d83fc415749b0ed94c2086d77a7914f8712e8dabf1bc3c623548f5575930f99a06ee4d6c77b54c28b1d9455f6d10e5f0c99ad3d580e4660fec6443aa55e00a95b1021313cb619bbcc8db731d11c71949819474673a9635771a7c34752129bd3d2c9a525d4094e306e5a2ff4018c9e67a02d470fceb5be222130018423a84b24e6db25ea72455a706317b4c5a6747f664c54238948e86206c2c77bcd003f4787bf07ce1f1fd74458fe41fbc52c04ab611b91bab7f4744b8c5d85eef160bf90a43e24d43c8b68d323a26aadcd837b721c78b45cd6762a4c6fb8de6398c00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9822b93c7a28ad4f3dc4bc2421d8fa1f92ebb67a67f002d766d9771fe9a778ef355eacb22813644a3d5e82e2f23d82bcc00a41a18e1203f7edf41b21a50b7a233c6647d8ca10e848d9f2b69db08d1e00030ba57478619d2a2c919bb1c70e4fcc23f8eb1dccecb4af86e3a5d0915ea54faeabcc05b86601ad26b45bec8773b7907474007cf0d21bb50ba706da4656f9c83691bd370ed9ada1b68963c79f8de6216c51f3efe60f89410b369d73e00caff71750872435c97166b9b04e271b9b99d2e1c2a3948ff689b968ae3fd225a774a124570035af842d20ada3d11110985d2e82cd07dacda42d0f12deaaaae75b9db04a93a57567cd67e700089e8b2d21096ab9669cdfe10528a21f0e6fc8e0aff456977764cde31af1c7df636042a08e71d9fd4caa6f5c0ae5582ff30e1b3ab3478ce738a34f2565633f04deb938450b853ca9fdfefa5d088181f23ac99ffa1aee3c04c496947d6daee00c73e34cbd6cf7355072ed3ff28a4e07c1b98566a9159c9d817ed5c7a96093845a44d136c7f43b0e414aec2aba8389eb88accabffae7e9fc0f202dfcd903a38f7a2335a465fe2f5dd15ad90ffe29167992ebe023f4633b56f1775bb1244ada215ad79f1e777398cbcfa7596138c9310dddd873a3dc5a02567e54f23a16d0b3318bd925fa3f9b4fd0dbcc21e4f296508e5c1c901b2190f0e169c7d4b3b08999b0cf6c2d43bc810813e0d70e83e722bdbf0c167fec3797723b2de781cd9289fc5769345e09ba2a060e77d5107c6d0daed126c9df114f96db2055ebcdb049304f12a96a58c8b904ea6daee8554a04b4bc4250013760235640b6901b48521042a96c9d90f52d30c422bd8a43630506cfd141eb5360bde9b468901e29fea0674752098df8131b0b12fe4f862cecf56b87eaed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbb536462299deb34abf610ecd124fa6b593d39c0498bc35f82bbfd9306f9e202a240aa5b608c4f1b48347e21e0b918140a55953659d6d34aefded07640c69909c8711e2d9b862288938a2f7f7d5d2d762dc357594f6f00431ae5ee7d093a7e5065db990006503ed8c964c90cee2f9df21e3b8158f1ace7d7835d3714449b5e6f21b81eba3c7b2b5f9ce4b4e98339ec0ef4ed55a303b4f839296ba2a007d6ffbaae023f7051ed318f070b66aed5e5e84ec42502688a72683ff03d190ced5ea7a08eda2f959cfed16fbda75c1bd93aae6fcd82ad8ab18a938668aa39d83012ca573888e82d0534c7e29ab3df52ee32a158d5b5484aafc41f1e89b21a42d3965830d85ae9191a4fe12a47b84642b4ace6cdc1dd012ea1e45d5fe97e4405ae94dae22ac316883e2851e1c8d9a5be06f9641bc416ae8706dabd2193d61a80ddc95a5a066a5f1ba9cb1e349da757f787ee5a1d18d8d7262baed0394a76337a1adee5484981fe4804a0b3e85c86dddf832c91d4942567a8eb7f14b53ac1bcf19429fb32a1159990bd21c846fed4d574c26f6b6d1dde43766f28f3a81a1696e89a44673be65274d6b6534e895d939911fa8860a7156e4f464151aa7bffedd25c17d92cb0169b28048ba685e4c2114af6d22912040e951ad3d508ebf4b9a21d1713dd7e9b05706651d3b16e55cce3eb97969103db33d344fc9a78281fd8a2ed1ea8128306d228a44250bfd791e1e2734999f7c5784dc60622dd74d4dea38187d9c7a84b4d361b0422f04bafbeafe3861e77d17df886d95b8a56c632a801e7132f876a93197232665f0140a3aa3c35afaa17ffc0be7b9c305a2c045461517dc56b03657752c55a28ba0c6f6425ba375456ddf271ea8ab5600333bcea71cb8d702ce64534574965e0684ec77f70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb1d9c05b98e9f4c11d70967487e1811e3e76081cb02bf947e1d64f834ccc4c12e09239d530933959701c5dbe25d04ba68a1e74b5e7244ce6b4d36522254f6fc5e91de8eb4605c6c894a465749d45884e9b6cb7f6d549dbbe418750dae844dd4bdd6cfa01756404551e702314285e420ef2aaccbdc02e97f52674e3ebd48743edceeb3d51b7e7586e6e37e75b321dc12c3f30ba6ddcae559da356fbbceb147b6c5e7a2b871910f85688754e4322410045acfe0bfee8ddb547a33fc61a8502e873266e3ecdb558472b4d32797952be949966b1bfc09e8c48bbbcde02b01136431daad79f00dbb412865a224b10aca729eb20e59d363e64583ad4c9480b913549cb5b65a35963f07d9e1da04f2fa0124bdb4fc7fe5fdf34e07186f498f04ea5a6ac847a6d1f1de0219c8152a2a9f4af819099a758114b89a889d93423781794badf14f41a7b9c185f56d72b355f5a1524268ec95d9cf32220805fbf3dd48beb1cd68e222e8c858ed754a49aa6faacbe070693101de10658c10642f4d6155a8d2eff1b1d52bc43bbe9409a2f2961c18f72f6a373568050b4c3f270b3473899844568afcff032824af42a900fd5e417fb93aceab139d2b06fa851b486bc9bc0fbe7ff60eab26f6e5d0f40418b954b5ab7633bc6fc332143689606a3e53bf73fa0a91ea0ee0cba04bb7c14c77a5d0e902a90e924a3b11f5f99e4b591732497d8099e87f3d2c74f5fad6e2cbc0f73d3d4513df05a7e2de1fef751fa7c6ec800b6334b82c57ec7aa09cd5c981a62fef25d1c7b9262034af7ca39aa79e374fa8188c1e4e08d2581adedc6455caf2819fd3e91f23f3e55c58571e0fbf53b962f80c4ce03a0273517d4148bc38713acd47b619be3a8d98b8150bc8514ff2fcdc3daee85d7de1adbbba147f0bdde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9437f14d4a995632363d9b0f49aa242aced237d854eff78eab5d707a158036fdb15b30723793b29f89e19df8cfefa7ff31a5d05ec983d9cc2852433ddebd1d3a8b483e01cc32affd13438578ec9b2c975aee1982b8822492523cab8e458d0771d1518410a0804307c1cb8fb0b8d3e997309711061f30e8230a2fd2ed2b0129e4616f04805840216e2d037d2cf736aaae4b69d08b6ef812d13f5883b6ce5e704bc643b641b8d1555de029368c3c5ce68c4382e897e86d277dc4b19212ca09807be9c3395e3a78df8464e960bb398c34298bc73cf970dfcefeede3dd15af9e754f87a7e187bd6bedea0f25133b0714f1593396d7f8f469591c3e5c7859c63db41e26ef1f54763019d7751509c307e5a68bbc73ac323ed04c82630068fff30e1756618b8560be8791e17758336650906457a7e8775327baf0981c7e1e682be508ce652e74d9a079c5e021d69c361eab5666e905168aab3216582838e1317bb8a8a39ef01840e3aada1141018088f2aafc1fdefb3f752757f29dae7a9bd6566f83610a8d3b0f334e33cb1b6f98f07adce88c45b667dbc3d763fc878ab2d458dc2ec7ce6486ebc55029312f9d261dad1ad0b18eedacb9f3f9c83375b2a54170cfd2e6077ce6ad9c0a23565de7ee462648f0ecf6ad4ed6a53283b9a017c0b951af68ec6c54662a1ff2b3876239ad12cd57c1a7ccc59dbb1d70d3ac31f70f9d3924374239632e96d9b0710aefd8e64dd0ab50c01b6473b412f077bc5f62f9494e41b7b333a52d8501b7885adb9c5f25c86e6a48b24d9a2bb7b237440c3939fe320f805d9672f057705760c6ea374625fbc946e6c6d0f37f848633dad5f1cdd1e9e832b3ae209a55dbcb13819a4017248edf08573e6aab7ebe4768dd8cfa9d336eb7187fae6a3b50ab6206d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7e34062f74f0abe07ca0b8dd9c7137dbb1b0cbf7eef68ee8365b3c1b71ca3315e09b044320e361101844159a1167b73506bebe94aa33bcbe856ad925949bc0de61ebc953b76508e7775222db94779ec3dd40829abb349e3e6c19672094857b03f6ab1b4b418739658904dc8bca30aca825ad9dc9118ea2b9354fec3be195429e4ef290c89a2c1addb498e39a4b2e672e3dcfe51be128efaf43d8e45c9942f4ffb17405b21fa549d4a39b0a43e467f76e1f208056b040b7cc4876450d773a46dc26ca5f9034f65a7418e412cac1aed93e9270b92737adafec1134a2572ba5abcd63685fd0b6adba72ffe88ab81f06fb5bd40a4c6ced0604927d52bed45a4a127177f5eb53447f137caa05be50f85f6749e5f3d7bf21da984750a915413c554180c5af4615f82a8284cd5f7704e5bf46340825e70a9f92c6d4bf6daf4a9b004f273955bfce0e4c08b541614a0287f7e1d93aaa4ec139349b38d532a776027e892900aec99cc952c074f354db9f785af528eb8968658816be47c1d6e4ad54dd817a587f1aa6b990ee83034083c128ccb72636d89efb36d2068015d0055cde15312b653fb399584f1ae12ebe0b459057ab55fce808d09f6b6049c04238710cc02aeb321a08762052fbb2b15132e0533e2e338d006f493b50bb0fa361aaf3dfaa0b9a22dc62088b9c4ba7908fcaa8755e134bc42ad715bc4ba03277fbed2393babdcb74360f7c4286dceba92b870437fcbccfbd1467de3de1c6af1e7d2ed0cfa0e2443d420a36fb59c32b63e851f75902814b70187d8c9bfad0f89e668623b4ea5e0d7a14c9614c17daabb7de35940cf87cc5e56fe3a8d8f1b983c98bfeab8a1adb4828d90b24b9f5bfbd53f8ba75434310c67d43193587f24f9252e23564e9cc11ba067cc1b7641ae16d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h92c6e1fa4f48082721e382d2e59b4674fd4af9ee2dd27bf1d6b7bb8aab4e82d90c4667d0b105fa668b82349715426d2c8c2d566f715032ea5e0cbe285d42dd105cf58f33f03e8cf5310a988e3c601733abed03d303451030ea89c251cabd44507eccb389c0b36d9230d8725f427c1269bee2da2eebe5e6b1a4e530eb90a6673509fdbee0a23b7babc1e4e5a57ef70ed9e8aa46102ea1a5251281b75a7d1d6be535800682c720a84cea7de488fad0c5f3be2c8b9fe2b6078f00c6357b20b76a89914272495b633c9c54f9e3633c5e95716b29cafef948d0cec2c347b2523f9fe9666fa7313bc7031756a3743a0ef85ca061bb6c6c63df22adcc20286b1ddbcaa23339521158a4333e5484574e2ac492bbde52129621519c329a1b3c6487e32b14cefda57c4bde336ce1d82d19ae01677d11c629e1529009ca83f4c82a801f7366b7e0b4600ed316cf0fa21095a805cec5541daf0cb4d299eec9d3b834c4088115e7223017100871a5d2c592e2d895336bfc07209e7d1c4d9de0ee3a04bfe10ee2a40ba3e41ef3db2722d1aa7faa45187126ada3ecb03e708b591b303eb11541d572085d78ac7ec1ff477e0f6539c1dd25a0db452b53eded8d977e0cb8e5c41704b896b74c711bb21ee1ba081f4cf991c99c5e936524a0739b6cbcf29b6d91d44b6ce6ba9aa132000572f2f67c619e1847ea813999e24ca006d9ce691f5282ac215344d55139c839cc96b1adf8befeceee6b53b9cbf6a22366aaee31ee689bf18f73f2be026187adff925570c81bd1cc9d6864c358c5a74ded0f693a3b8c21c63fa4285ab9923373f7db81426fa4d4939d0166b8e39293a7392b04fa5d9557f1bf0df741727b7ff3fe09165a09baa168e2e17ba5d9a59a9d3c349a11b291edbf5684f66e1446d188dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4e881d6bb92fe26dee41ecb1312709ac30cd07290356ebd8ff651ab2f456236bae1a45f0f8be24c1a968b8ce47504291c0c77a2a54619f46407430d716ddb9b253f01322f14b70b4130b4383b15e2ec87be2d2fe6ab20c37f0ed9e8f93e4ddd956fa459a00817d34eeb7e3e99ae7644fb0f5a136f6740b16db8b5ab3f1b413cddec5f1bded77d0cb64179424a25e16b85504043c47e8ea0ce3f8e21221c0f9acf48d292602dfd90a9483fc03850466a2738d2a4b80b0598e8e1600b45e2992f129edee34fce3bb056b6c6e139f31c7e1b8d1e89ecb5dc3549e6bcee5aa59aa5c36423f68de2b285bd47e6d7b651e649a27aa7e27830f71a5ec08ba8c0ec9f16d5562b76ae295e22fcc3c89e9c05a8392ccb425ec4d7b40a7703b8d05e1f74bc633b1a1a063d55e6dd8fd8fc5a4e159909ab043adae85a1fd3f926de1f1a01aaff0584e4fb9457b3775b94c6b622af5af7f953ecd3ae83b6b4e5e7ca7645c1295cfb22b2e9d3e7a10f1ecfa5768986cacba217cf706216705cf7d96baddeb727f970693c721fa76b679c8842db9411949145383159fd76ca0ee1d0d5fce61c11f67a239f723cb3f29f0d357fb104a206740ad732a69a76ef4e92d7c99532052e24db9fb5b06ff1462da6baaf9cb38183adbc7dd5fc5137e1e31cb6eaa56303b619310e90e768fed273afe11ba01d390ad5b91f725f67997b4ded3aa08384c9898b4c325087d6a3222539a3b8b441136f0f89b7df85eeff0dc5f040987445d8344f708ef12c400a231063b8e5c3e5e7d03f1b09577b61b7ff3bcba2d39b48175f27c902c3a06141c92a32744530bab5bca214f131b13fc9084b8e14ef7877da1a26ddc24a422f2e7bc9721b64a8cc6ef14d19c516d8c516a1ea58f961ac4ef73ce45e6c7991f70910b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h70a29d84bd114a42489b4e3b6530c8313de2bf189b907be1d89b8cbc8b4551ba9504b484af1c1f7da6475b1c1d4ee595260a12e09b3198df9109a3b06f06d0d170a78109ce3fcf527d9f1808835a1cf9b50101348344e11bdc9d8dc3f30760c6b9d6807f3029020dbe1ffedb6c65de0e9ae585974edea339aa3dfcdef2562272b8390d8abd3d76a1e7a993750be2e91dc6e738af0dda8560ca31b8e0fbc6d6fb76b6b03ca2ce78beacd11f3b201352fa49f703c426997593e13f86686a5080a70ae2e77a97719753d945ec0d7de63b07c2c14a7d67caec30ad782b6584a88d3024ba09090139f0cf610ad2f7985b8331f10e4d1ad2db994117b1b80900ad80d7b7b63b69d0d2ae574fc44cd1c539666a415d5b76bc0a74b804b15e76f22b6b6f0f70baa19f67d39dcb6afa905c38fd3ec7924fc17eb694de07d977fb1a55c10f9ac47ece8d2f02e39a917edf95175307298b61843fc7b0fe91198eacbb622e557314c0db8314c5a31bca09f71afa2c6e2c342b167199d7fd3713c0cb4fc3ea96125b2d16922068423e7391aa3aebb86f3e7d3059fbb2608378d4c7eeb058eba3ce64178806ac0ee74005687eb076eae27a459190cf04042467a35123fb9b02722660c363dae2a064dcdd56aab49c8bf9718539eaa2087e29c923b85a65e4acac11a0447b87d8c7b7a4d80e6b9e565350881584dbe322f69311a75cb2c779961b0632e4775f9dc6ec42073b673ef7c032d1862d6b01009abc7bdfb837acab8b7788fedc2418f0d9bb450d67d3eb925b3cc7b94422cdd662d6a786b02a733ef1ec52d45644516700bfafc01f79b4887dccbcdd022d8e088bb3664dc1a52f26ec5cc6424b4c2ce0900ff5dff006e983bc9bbc3b2ae7ddd3aaa3777ef0b4031236616e4df0217bcdde8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he8e8e754ed805cea04dbd6377b92b951fb96c6ad3c8048d0521f7b90cf3c2519ef6f7324cc415fbd1867925cfb6dbfa059e7fa91f66e8731aaf481144fdfa290ad5207c5d0a4e8ff0e1110d62dd44ab76ad40d5b45983472038fd80c9910c2cc446d6ef940419c0564b9455b6798b8d4c72ce8d39412fcfa399893d3237fc925e5df3eb77b001c548cb4515017435dd67030774f52bebda98ba0eca905db2571805a2d3937a3e1168e4db47a98a5298ad95ecc76321df6e571ffe5008010b2bf969d1ec0361647cdeec81f56ba11bdaa90a6a71d82002cb64b955ba8011d67af7be36210e064c113de10eefd1ac55f54f6dbffe6ec932ef048ac5f6b9f8e9fc83e57ee95cd8905bd77c335593e7cb024def7692f60baffa36f5490d7e16d87846c623c29cac3ba3d660bed4a23a6f65d66dc216080fb7ed11bbc1b065a6f35d6121812c434cefccf75fcaef181a65ecfc3be548f887aa8b3ebcac8fe900cc2962761190b40ed318d97fe6123e2c1cb3ab5c66e3bb4a7df188aee6dd24986e97ae84d9d2456b3529c7be4d516eaa6c8ccec79f77ce499ba86d5b9fad78eeeb2238b929ad23b06b054a87c57c2576915346463d48903ff6c731afaf094fb04a1ff195ef4b0903245ea2e79c90b94ed308716518c2aca4a065467f41476ef0c190e1d1f7b2c4e5ccaaa262e093f74529d041175938e3669afc748ec9f9e858dae7c5ecd34f56b622d9cceb2de4427bc5fd41ed6aa35659ed2a99ab09276af714b641c9b47a3631739f96e517077698b18e6fb67797b5a01f2d8e758cd551be3fd953ed2178f6a78bf522c1e8e7f021dc665cfebd9f1cfd5dd9b2e72e27ad8dc624b71ad64c78b3433e2b8478f97a62b28864957de9fcfc6525a10dcc4ee5f30b6a65c264ea77a1815e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h36f6f53920d32da5472053a3fbe4fb54a3bc4600b949a17a6fb22843faded9a13f09429bc9d5d9212c6e9a65bf14cc845900a7741a3668e22519c73c74422843987a9bd6fef6e9840971c5bc3d85ddf2bf0f30695810bdc188b05a6b4489e46e95c1dada8856ea09f824ad77961e8da02afba64037563d89fc1d4ab41e8e7f680f7f7f5a3f9389d9697b103ea74431c14995ccb81adc7ae5f615c6cb5c47eac38633c158623cf29e5c23ba7a772b3dc10da9e4f0c1722abf0523bdd8b29eb530bf830cc1a8382c6b8ac4efa96386f107b39991c89931e6d1e03c1b47b87b24b8c981d2f059c3bc41e9ebf402cc11317c939dcce427ad9cf9fa0ff624d1341582aeaeeb73556a82a92296307ff6d4eab1fb339ea2a05e9dd22e481ed610d2e0ddf16907eeba7e69be03633f6afd8b957705902df20896259a489409f83a75ff94d4fc211be150564d0a77eaad15509f8011971e8bd348ffc0405ef710bc704e521a02c0cbfd5044dd4219403399e1d37aa3f9ddd2c70cd8b8a2d425a9eb7dff4654927448c762219c5815c08a13d0f854cd8176320fff0d0d02f6568c8a55e7c190c0e961175438c629b77c61ecd36ffa87a517f09d6758b8d622f1341648027b978f842240cb4f54aec97b43bd1ec9ff60f454e845bc2ae136026ac033599ffdc4ff3e792457f2473d26e1482f590e2ebc5de2d2fe75b442d2a52b93c6e93f32ef6a7498f4ac083aada5302d279450447acb6a96a53a63574374e15c8a7dcfae93628db46ff8951b07a856ee75d3f245d8064d991522e81df75e6dce41af226a143a51418988d55bc8908e73c3ab5044d4d55cc5bc87e31831bf241a51bad5285438e9a924a0a9b367f66872d7db434623c866bfabe568509060cb83b85031bb3a7998dab88692e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h50d9378eb81d89d3d79883b88df7da7aac0ec16c4ca4374956221e633d5e5ee623f7fa257b0347b04da2c4ab18c91fd4e7cfda286324fbc8ebbcf33fb647a4c0a3addd54dd5e6fc4476e24cc4ac07d76ff416a8ffa4d2a3c63e3254b7f56e5b07ac003c7e070518775e601dc94a4f95e3687fb47ef0d1472f7a4c252c3dc368352281a910a8d2f196b3f42697235a9a7b92b5c09ce947cb594f9df9b733d24163e3e77352a11a893615b2d3cff15d8936a6966bf15a2ea8e9cf83e1c4c9e31d7596d2cd698fb52ca79f79d63e6f6d5b1d56b9987c8834e09aaf7d63f886137e4da59170d96971a873537fa9e1b38766c650158194c44158d8602511ebb35bdb8955eb1edcdd6c472a8feb3c5e252eb610db2f36dc3cedf7c3263f058e880964712d1e52b52f2df3ec525eba0de4ccebc4fea65ff793ed086a978882075092611c0db3771a8665f03d1409d59c23d7d35967ecc60f2c427d535c2c704f848b7212fc30d94af70b9839cdba99a8c14b7a9775447df7cc73f16b7aa105ceb6050cfd3d703ccddab5daec3d209ae133159b2c53888901c0052b24d5076fcb8a3e5e3c9d1ec3460c7be14a1943034174c10d6c8d0c99f8cf681620c419d7facb2b959bc6fc3ea4ac82a9f4834a39dd5d50f9e0fdc2bbd9d2326bad5587a11415ef219248b83aa7c9da07e99fc277dd58f1dcb2c72fbe025d8fb0b0ba22eb607b12a43172d6e93b2992840ef12fc55c82c93ae2e8b24ac1477f231886b4c9b49feac04f8abeb0f742ac5ce95f3c7764e1f21396c802e8cfc61d4bdf2369da93868e9a4417766e8734878d9f87558e7ad173a76ec6ea67e76d568a1df43300e989b22cfae69007c22cfd96277be0eb625883d289d74f92e7c09670d0c4a24946f5438003086d23fb80f5913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc57a9b7df6aab7d67c9f46c2e377ce35ed5f0a5ec6ed4fc79c201903f9f93828df6e7e4d5b32b3d472f3a342b7042b391176ee8a1f7ba284e88b8b79d210e1480b9e07de523fed81a480e761a5e3401bab5e9c38298f14b5feb7135c6c4bdef5ecd3988c2a1004e7429687acd1dac92fd2c1933a94fb950d627119ae4e69dc1f61473a47d2d2e250f080fc3827a70d42750b21c36478167d316248885b79f7f6b53eb24b90161ac5270177334f9cd96c22a5c5c3c9d375b49bb9b3d96542e5b028e79f968d2c5335e00431d6f42f4dc8e766bca231d8676802fecf1c54bd2a7433ec4f0604566513c64aa1e56dffb5416537e81f39734f4b02464f5008edbd695e4b912eb09527dd02b7aedb56b106643301c2ed1f3c81f9ea906aa469690385600ad5fe19000f9ebb07a159e000ed0e53020006ba581e2aebc984fad630d9a349973b37e87f5810de3a535ebea2cdaf5b69d4e1790b51e7790a88c145ceda4f0e6dc8dfc5b201e3676f6a3392e80a2722d481ba872aa446d881e7fb712e842f3b752ed58a9b2dcdd467562e9319027fefec1600dd35fecb68152604a014dd4717f073c627230b88a3d0cff2eb944bc0e0a581bf48e6de5b722b00923568d6c6af1cde155bf3f51cf2f1f9fba16670a9d84d188a622d647c85cbb3efa8136835346d80f12f47920e0036fa796ca28ce279556e837ab5bc530b693135302ec6dab16096d248e213327f1f652a607568d32f6e0aad1f8edb9789ae1802da222f65ac59ddf1d55e6d7ad7fe4f29422cceed4e6366d9c0b2b0bc6f7260b093d769937fe917c249187772294203434ffd6f77f95c4a8560b21dc71e603f03eb566e1bde99dacef59e8b858268d1089a2c0882b526b0249387c658e297d7ece4d27699f141e858db6ca5cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h45cc20cf7b0ba38e36d4f558212f46e10a9fe8465e51f0341b76f042ec4a9e5ff2b0e8c27e71081dfa96d26e92ece370bf5cb4ecf1983dca99d27ac7fad0f85849cbcd4fbd9ad75d52e249526ece9055f4b557b3aa876fa1034910e1e7896f19e2b181ab6fa2ba841444c93ff573ec491cabf6dff84d33945cd3c52e776149004a09cc55e0a9ccbf3ce1e39b192970e405e9cfc3febf24c5aac8b6193059392243cdb260e1862fbbf900d7b199f979afee50ec6bdede00788bf479b98fd06398b08a3479b78e2956916530f53675588e8b30a7f32e18356dc257c3067a644897f399ccdfc27297f5718f3e70fbd85f258d77aa6761b90592ab8a221ad91161a532c4be33dba81887702f4c4fd6933c048f147d936485d576249662042b424c4d62838bcbc0592a3f3ead60cc592332665b7cbfdc0f7cafd6c9e8a62df583528aece93e7140283760e6cfd5ae19e33b541e050ac9f4e139d255a001e2d1159bb7f5954d3122326aaff2da432dd967208a29ddd63d36cb6e2e5a713ba5a4674e59d78d1e20611c42e7e90063b9267fa86ae624edaf8b163fae83e3654399301d6c6c5771dbe58f3d392e1a1fd2a448eaa2f6253f70f5edc45d48500ed87ec48f10b2c741e36fc80df75942e2bd1170c96273743fde48c3a8c319f3825cc2b5cd0b5a4fa339f66e929c8f240fdb6343fc5f9cbdce808afb80f36123c97432365bbd27e556584def2be72e3c8466620ae854bde5b22764c0a80968c11183aa90e8094403c6f70d6cef62b1af6d5f44bc159b7e0cb7239d3d447794b5ac2b02bd6eb4840c5a90b813bd261b9ec7ebb21f4148450cd648696a6d8cdb5d416762a5e860e0ba90a5ea2264aeb491e2eb815f3bc06ac89ab8aa2d256f4ef79ab55bfcf95b34056b2e373492bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcf5f4423a79e609b9beb21253706c40bfa44677761e258b3a87d1d53622a70f9df7ce78fdec2bb77aa7eb5538c4f607ef4efc9b90676bb6d2690077999c9369d8e8c8762ebc1d5330d2ecdadf3ec30208acd739e38c04429880969ac9fb01c354489c685279b20b4a5de7f6f51dbf2906cb423ff719b8226c9f56ce748ce3bdc4102738962f00eeb485a41dfcd1b1acfb3a8491d8e69f39d7f637f929139244f35df47835c2b63345837c6d07d98cc3e6d2f7c134c6e5d22b409194762a6f743d85bc86efd25f6231c92a517cb672dfe72ebae82746301d953b5e0c078ede48f4e7af5cf5673ad217c133dc78d50218f98c904eee3b9b96e1f132ca58542f3b33297c1117b2d7affc5f70855b76d291fedcafb493631ac68892308795362c1098cfc52e309c4ac5358bd5968798a5ec731685ccb78a0e116086d0c67f23403d0fecc33261229548623555f8dc33956892a013a7553bd627dc24b457a5dea489a99d14b675d3148cfd48edca2b524fe58a6f0c805e456502cc7fda2b41cc20da0452e969711da160d4e920a86f1568d5fc591d4ebf03d05ac055b27b67c480e663837b06ff754199c346ba921e620e9e842e85ccbac47668c757cb0e3ff7b34841d0b6845146b9d7ed379b5a058c06b33e7fa3de0177f84e5ef262e459b3fab3fc5039989024701e509f97e4acaf9e25dae70e07d91e944aff8ac471083e6cf5edda3a12df6ba15f35c924bb1fccf47f1d8c680b91f5a38eec87dcce66dd71f9cdecf531229507b910bf7873a15f2b9c63265936a2fa89f218e7c090bc13414a6e25bfae30b15935769b0cfbcd79f236215e5c0e924dbe5a5295fd178264f19a0c6a5e6e347429b0d837c5bface6da680c37a5d8682558407525dd413f02aead0a06c709e815f6cd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf5d2d5b41000e0cb7b15101720dedcecae45360877c31fee4c9af3f71f38631e5bd6039f6af44bacb14feb08631b27f96888ffb3f8e38a0be3a7387cf9855b0979920a7c3d6344b386b40d0854b1c5d3957109e055b154ba31634e461cbda5d35930fcbb9de3166dd581e3acefefc4a1f3845a5142f7ab8b3c0d086cb87904f2bb4143b0a02878e91317f1a55562fbda1181f40aa82701410273c622a659d21c64115a4210ce98663830764f1f04ba589cbeade5dab769cebb1364c74b72b26950233b94628e8199d18035a6ced05e5b7e453078c2c35703ca1fa7f740ebf1be5a1ac524603e8a6089371c2515d73f8cef9a21a2bdd6d5e7f305f764c8d59797b3bee4335c250bc1e7561201c0fc86e33e131e07d9581bb661349593a0ea391fccc1854bce2f1d7bcc697ad79cea1ecd568e24358cbc8913c65ee8e522c5f4a9ee1647b5875fa3c125f71f1f3a1f8dc0012a4763f65787273121daedc8dd0f266990dc2a26e114cb6504741f027bd418cf3af1e2ae165462cfda48c4163f98f5b8fe1657347bf9dd55434ceb4e7bc0019bd574673b9e2067186b9d319353a29dabc916242ae0a4f0a53a5ca88c554cc76c2e320b5818496584462b8c9e868e17de8f0431141ddca4acfb1ddccd70b34728cbc2544cb58bddc87400c13cc2e456d9ce99226bac60fa894da3634f6c718ade6250df9efa54d607cc722b902c78ea1af6d84ac68460eab8ffc1c0416997a75a1e7fb7958ba43dea6fd6c20324cdcea2243dac291b04a1a41f46d7d71cc53ab2257bf740f36aaaa9ed01a7eca2a3f0961ac25ea71e3b71c51d51717320c50aae5c843b86f3b6ab8803eb321e5e822c6d6955ceb0a555a4bb373c7846e65b282163214370c0c67cf489fffdf5395b23933cb3675b7fd950;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h2ee5bce7dde06207c54e1bcd1b7a2ba0b2a86e2d6b90e7e483a270e8e3d1d9a649b952840b566dfb07de61bd8e63d87749d21d9274b8bbe4c6d8b91dd3e3dacba426376e6aa292ba2c8ca03f6fabbd17f276f9c74ae582143c454245abf82c77fa5e6bdebe8470a10146faad6c2b81bc4b1cddf3d2a37564724c7d5f44630db1acbe1fff6b9e2347f366286787fed5cdfcd18c81a14047c66676bff1525f5d51af22a66875dd30854151f1e6e9ad17a6cdd0ba12ac39f63534928e538ecd872c5a7ac0de397d5d901eb3ce1873315755902154e87e00d8871aa41a43c68bceece387ed3c7847000b4f66198c5097476bcdac042ece3f0f38c605d718ea602080de5971540987fdda281da6d7e83ca1131b343868a05c99ca60aa0aa757af6aa78bff8dcb858c1b144ea1f2761f326edffc617ade00f1332c6e834e12f4bd6a42469254e54b734f8392a16f4cc1ccbf0c82cb4e074b1edadde382951c915c439cb07a6f934927e392e79e091bdd4bfc01f8ddd15b465ce2194bb1ab0dbbe4c4781d11e3f368bc56de0488a6595913a354ac8b3cae99334ca2e8779edb4150c3bed093adad65c918abbd2be897255763d432d792d138633b26e24f4c99ecd7d8a34c9170817f381cb6488dcdbe3aade53fe1b7d8ff6d639ad7e1ff241856e24209ca7939a8ecff8784ba7d58adf289f9c010df03cbf2bafa0ad943cc5a53add7ae4cdaf0f3de66536514285993f5db6b427b25cef38a40865e2f6173f70c09ec42c80f1493e14d63d136dc432eb095854c10330d00838dba89f8f1a9e7df190b73f67849e27ff924bce8dd5b3bb4ed1dfeab97248c127fb70c318b82878d0ecb6a10244574978dd8cd9227256b1d3e71738ab9d759eaffe347c200667e3f19df7ff0895e12949075ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd05f65f0b876d6e5268113ebdbcde6152d9df62a8bc7f61287edc54994a617e784a9bbb96f4359cb5ab725d663d7807445bae933d2231bf96a21a4a5c731c8ea09f23a6d1807800a4fad0f0cc83a95be48f5f8923ed3e6a6f372b424230f132e0763b6fa982588ed6687dfc0872f4c9fa2967a73145e3063197e13492163e1bf2f50fb06976ae911531e565087bb8b118e583ce38726e246caddc1d2c763099dfa357ff2027edb874619626a52afb94d4bcdc86928257d17a6f5fa966683a4c538097f0a5c5fd5b9ac7420859ec20073e0d64442697639c16963135ffc0692f53255cd50cadba6e43585713af982a586555b5f9d778bbae2706ed8fa30a763812a62e89021cf03b4137d918535252e918f3e86fc709ff5da9ca9e89a6c8f094dcdf72841a74695ffadf2bbf01017d34786aa27d3af165293438eee44a33bbceb1d874007e1bf0378dd46c87dff890938b1712726f1e6c882943d7af423ef6173e777b8441edc5ef7ab745eb6752d8687ae577a9ad73367ee2483e0c4e0683c376406c853219914311217e9406bb7a27025c6964edbd9e6f729736c04074c2ba96ed8e557323704422cd000dbc7564dda0a32d55fa5c7cff63c061ee12ad130410195cf9daf0aa18678b8e6dd6c117218dfdddf7c28c69a9fd33f7e1ab7e4e877013eaa773d49a5ee40ca5e44a0cfd39c7ac33c59fb4dffb458213103f1e611df971a3ff58b26678b40b7acf45bd8469ac6fabd4a1144ed2ca58be75c0432eea1f171f6ee4ebb513893fe360ef9de060373f7033350b2e4edf0edffffb8fe81e6386161e6369abdb39220830a6a9e8e824ae5e61c6a5f87f3da23e111554b0054d6f335687e0c2f1e67f07c742c022ba950b4e36a41334a8e8b4d78bc5f24284f5f117cc610d75edb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc17a530b2d194c9ff7d9f2ab90a7de789bc0909bd2c5ce9d18b38449c9197896d6327ead3d2e30f1e0a6ad21673cb820c0203efdd832844c947eba8cb373e8f766a29dca938f6c911476cf4e89c48c81df2448fb1f0836271fab3636eebcf3896f16411e998acb7a28c196e18a2a8c0fedba216086cfe2b8e9d3b135c794862194225fbe1395d23e44a4ad2a8d66ffecd0e97824b4657a64f90514d1370fb0d43782015eea6704de0e5dfea16520e04dc4e00c5f988acea9dc45dbc44937e2e3e49803615312f0970692f97589e23aa2b909fffe3f9622b9e5538e4b68b2d08d95372458f3385c63db56e8b82807de90185b5dc0c1f71faa0645162b4dd59c635efe8f04d69e90504bb9beda4b2c8c78930be03adf152e9bc9cc526e4f68f096796a1b2ddf3e00bc066fc41bf59580d0205c9f8ac614338a5adb0026d2d03f47a9722a956e926405f522b09ae2353a1014116063db0d7fbf5a5a64b1eec57cca5fbe96073addf7415b4affda890c7b319b866bf795632ef43e6deb9070a7960c797a1b327d3e8da07f7acf1661209c79bb041a6c305ac175aedbadb02eafbc8a4402ad3ba987d263903f480a02687049570280e250dc932ca2bec282f87e770138d9cdd6095214625881dc83f8a7c25c0e4da4004135c9f6f912bf89493461715b194da88a6107da669fac54f06d184ba6ea31ce8ab3dc649c51824a93430bf9f8dc06bdeacad6b783160b2ce8ee7ef7bf8fe5279f624dc486ac92bdf23a1901eb934352447c36bac5192ff1eaaeb705c249243baf75e26f7f6e434e9d550dc2ddfd8e892d047585b6817947be7dd5b104ef7ec7fc7d000a98e174e9193c2f7ed8baf44151544adc14f14e8f16459da040f4ed5e1cca7fdc7702c3a2220495fb3b1179846b035188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf25d64c212aeff80452cddecec2a0e6e751b73e04677966b242ddeeac44128fa9f055a48327bdfcb83dd57c20230f2bfa0e04c0d22a8e285993f45b95f9633bc9595a97f202cb56647438f6af24dde8d3a8ed71fbda32784de7dfd39688d35ab28a8a62ccb6a7fd6e319c4aab087720c8b7fa85317901b8ac8620c4530c5e6210f0e533a653847e03cb62254f83c8b852fff8a67270440c6265356f3d45ae36f91f342196e9003ccc77d98360423af6f639a40b9a608d62226b190e9e171a8a1d92a81ad3185d57f4902d3a6ac4c29bac77dce3e84ab18ee5782f94f90bda513ab4369f620c75ef9f0e67eab40be814f7f002aeba9f805dd1fb230bd5e6fd32aed677b2cf0142f782aac119f678f004404c8beb7df30da344eb0e770dd5bd85963f855f0b0f2cc1a462b50c4c7f0d3dbf13b31b0a330d5eccb5e5eb9b2b5da88f8c5d01895fe1e98badefe990fd66b02bed452cdca4566b0b745ec769c701e9d7fb8bcf0f3d6c0b17a94d89fec5468fc68a1e0fad723ba03699d15aba7abc61d172169e9fb5726e26ce38b3e12c0574da5b16ec599e928d1bf3ffee3cc3bbdbcd7963b6e2d97918262904776c34adc1b3ab14997f7cbf036652b9195c7acb42f31f328bce07448c49e0cd7c48b5c0f11257d2b27140251a00b6b1eb9899f68cdce82f0244ab90ef527e2aaa77a86d10dc56007e4b6e545806120275dc7289b08e8d16c7dd4b129de6afa9aa5899b99cbd7c7a1a63d068f80e98532b0912936cc8532f9f965b6139c3ed8acdb1af0facd61afb912a772068c2196f6ab3d3a1f2cae00a5a88ecd51cb74e697a7b06962de9b7cc504af94d80fe345650e77cc6ca38e41dfd98a9af92bb02be72540a08cf8fe4b067c75ca9f270543480abb803771d70c97fa5fceee14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7e2ce138402967e69d19520d63b1623445643af1e6267349ba21b5bdf2b3cac234a305711a3e72e0bbddaa6672f3c2945f0579b81e9d5eb06fe357faeef6b871e525efe0d3fea752c5ba5b25cc4140874269d5a4a458c8d1d2220960332669bbed6eb3db9727934a41bfbc3a4c75ed3d9e03ade19713eee5d625cde98eff8bef8bd487bce7c7423308ba663eaebf55698c13f5c5c5727227985e8466dec8b384944922aeae377e198c2135faefbbdc2ea0e0a5d64e7284e9ccadd604fdee3e1f0f9899170b27d440a7a1981d89a33709bccfb59194e89d7e8187dbc750f184be6a835a6f8638e41b026d22814d42bc55ab24e3def713452624b6c9956f00cfc33cfd3a6cb89a915b1ecd5156ef27312ce2b717b17230b79274f26e477a78bf030c89c6558c0a9bc902d8021762c507eab362893f106d07a8206c6575817a8d5dd89855aacdd3119bb23d30f67b3dee4492287f08780ddd6a97e04131ad5bd939dbd624b403c7d65e723f158b25f672f0eece80561f73c51459c15011abec3d39184b32fb6758eb04769a0b958767042f002ff3cfc8fe52b5aaf182d16f2496c3c0efbb36ea04d3867cb194cc5971e6bbde8a708543f49bea33c72e2cacf37456d0447263542ab6d94397b23a38f8eaeb15acec96d4a7b7c64468cdde331b474f7f244d8b09a4dd33e79b0354995faa831cf1af4fe5f5b8e5e4fd1d1b0462bd98f75cc2b6845763d6b1e5ec9e4754e2a3387d987b62eaf3da4d7b4eadf304a220b0e6089aae7ef17228a677ddcf0147f5deb61f80db1fd878dc390d2bf08bbfe52fe8c3bdcd4cfaf7fdcf86a8d7692a9a6bf3d4420ef068cb33b66e8b97b09bb33ee3f01f986b298bfdf519fea17154625c36426b98041b0f46064556016d1c10e8e87d97e5c77572;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h6f4441638cff985325da13edb59024191f20d27d560606ef1b31a1b112cc1bb5cd55a83eefa65f3b092859c296976c5d211ec7d0de505050ea2c5c248a72277ab6c54f974e97e4b55842edd62d54d22792b4b972a12e6423dc96d5a66dba1d4206d2728b03eb5595579813a091591ac192952031b71daa5d87afc9859f89fa7abeab01979f785bf6aaf48edb78efb724610a765e3843789afdece78672be82d78f4ce0dded3edf61a74494030eabdebf78ac34151f53659a5eb5f9ca2728f81b47b7f73e6bc4fd848b51b2739c7fb90df897b27621cf6b7a47abee12590e73c2e7334138f615268bf2deffcb5949967444a8a9b4dfe322841eb495fc60515e65e0f51bca2be7b66b0e5366ae40d50daf641591bb64b57be0c2df0d25525d2c69435d17afd4628cf52e3eef8583ab5fa87321e448021bb22ab8dbc15d4bf6366c38704e3f7889aab3606e106fbd1b0ffe6f073c184e4745c113c1526c49fac9ae44398fd40ab733462f04caa8b19e5bfa6e1f1510024036e013155be89202c13b9905c48aa0becf3119c857794eb1be8eff35de414eff9cb7037d02ab95d332745cdd704bd97991b3159eca37a05774c5370b36da2873b06c0fed8064849c714757c64922c377158fee0421cbcdb868ed1a9290e6fb9566481effe0104b50353ffaf790ceb8f4f8b88e31c60feffc3c2ca0eaf313445aaf32796a35c848c169cf179c1954f3427b658a099d2d54ea5b3fc6814de4328927b832769952b94842b2870db7bc27554db5c0505c4324a33c16f6a37164c9f29ab04cb515a133eb6e0ee52bacb808f411e4adea9d5f50fe3c203a615deebcec095c96326f3130a0b29f8bf0c96ce05afd6854516e140a223bb6385e66efb85a7ec3e72254de4a698207c78429eb6efcb088;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc42e9a215965a257f26f091de151b48bceb28bd6aba87fe5eba3ae7ff323d3daa7eaf325ffffe010ac570f9af58b887db291c3d665144f702815e275c5afbb7bd5a864924495aee70f6324588a3e6cf8c8aee737a7c39fe22aeb4ebf5f12b0bc1ea9c40d4bf91e0f32267bf3b68ce72553f64e49040376b10dfaa4dd630bff3a0a160ff22bb5f61d5c16dffd0da16327de862d7422bac55ebcce5c2a21913fb782548c3ca7d7fe8bf9f80bea1f0a159f0ea05087f67d8f1e8f62fbccb40053ac2d8e6c5eee8645e4b4b25ef0fd0247c8c3c2f55940494ed2865f4c465fe206d0bfa3306de93bec543c55c6850c98b786daafdc9e36d0b7463b2c5ce6505b3a402c63a3963edef76dd8623968cc16d1d6a925276ac753a9a04051a2725fd74030a0be6e28abd3022391cbce5bff21b63e368f83dddb58ad151331cbb8b9811d4e90c7d3ec82b2a6260c4168fa0b4713e984c9a3534eb6e726547416683b7ee6271a8288f449dbda9b0f86af8496f4be969dacc60ce0948e54149515044ee1a8904c950efdc8e158454ebac0b9e93b19a5e7333813377496863867461e3193707562dfc36f2fc491ac27a76aefa5300fe4c1ef7a2ff879c5c661d14abde412c67e0e550a9713d856b8bc5a930650f2585d4ba8df6da980005949fffcd626fab2fbde41672ea5644b493d9371ba0aa6f72e2440de5b81331e4dc9422d17cbfd23db776b25c42dc977680fe7707646dc732dfbeafdcd2082bbcb5e2f53c3cd92c9af0b3d0a63d0f076942626d036b678da870d4605c822e8046d76fa42f36f7cfe356e72680c59d58714cc6f58e5cfc149ba23de43ae861c603cef91abc6b02cb60f3638f84846fd94b9d0d91c2b01ba5ecf6f62ad26e69e65ece9e4f1a14370e2693eb09fa4b9f5e7aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5e372a0ce4683d0d48585437a409a7253d3846d309e35e00fbcae2b6ca7c9d1ab06a34f6654693aa093839d75c6b393ca097b9eaae4da2ff67b991d27378edff93ddc7002d159c26929c55ee3308f9e6a3c31b82897e2047dd5968a718523968c915294d81d7bfdb351b5b4390610384f38d6f36fbcf5c1225419dc79eea951ffe425bb6256c44bccd70b07cff09679e5e165859d633ceeb76c78616512d259e003a032a2503645ff8a61fcd5c5f0b28ee2f0aac16dd93b5ff26d288456f370b3281359b195a9a7e0fc8549ff369013abcfce8ae012c7e2d63c3252ec777983bdd82fd5585843172ecd637ef621dd5fe09825fe7d4f1b163c8e41b6af371b302c87c6e073f4c948e082eea41e1352be9b1846923fbc27855f44902cd44f114d77bc79d97d976b92356c1b9e10f493a38b8c6040086e7cac7e23d6938d002c53076a3a5b12b6069503600b7ba089afb9060e921e37622dd49494f9b3f9d6954a9706af506bef6d3743e3a25647d4be9d2934e0d558916677cce56d7cd131add270533ae401aa026a004fba3808977750a63ae30c951cef090eff0d5075a61aff616302f556555019d3ff4a3b38da4724328612555bfb5a31f3b1a8199dcbc583a9c3252cf32a7870f38bd9ecc780e0342317ae9337bed578aab6b53a4050221391939bb5d482bca327059e5164421dd8ba5c056644cb20cf39fc98f3b7fa426d37e38aac6081563df35d0d3493fb598f033d0e663e1d6da20e251927f85ec5afecf5689f3729c7776a330f4c5228b59dc76a723b58a46c4944796198e27c3373bce905644203885eb8c219671dbfc837df191fed6fa22a8751b26cab7106c35210ddd8620d256fc6c63219634a46365e9b462ad40ef66d28f7c5eded7b1620b7e205dc370218be713;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h494f0379be5c06790fedca66108d3bfa8d719cb70595097da8c0c0a42d05edf3115a8908f84dcf2709f85f1d956d43389b6efac729b45b6694f03c92fb9ca44131efee9493194b19b4eba166df42c3350cb75ef76b31d6921cd928edb0bfa299b8279ef3538c32c3f35f34ac63f8b4235c7f01f1e027beb2fea47f7da253e181e3f827c7523fa1ea1ac8a3f214340cc0bd4c6f5ac89737c956dfafab896f11dea75bbc1d701cb685a8e43f74f1a003050c120816b25fe9aa4c62c6ffc8d1a0cdda678768e19fd2cff1a4e3df50b5c7f49e7df9afbf394c04bcee08d05396086b961e4d0a95d36196bf7191674ffa56ac46bbdad6a892c4a0c0c4f94c4de60738755be05b89390cc9a4b67cbbcc11f30917f6213d6d6f37b1a3a613d45f9e63f83a47d5cc2e3801bdc022d0382e2589bc7ae189404f5235a1569d904f397a0818d181aa6a2407910383f3253778820f307193d9b71bf3a4fcdbeea9bec8f0f8ff7a30550afe8c7cf4fa92092c09c5559f3ecf507f8a83420816f2324abb6ce89af1c71122181f5c77bdcdcf7b3c622d5d84bcc7a27e0671ec210c134b15ebea4da59c9cc718dcb8689743f6f9ec48f84a945ef0690db74275d0c09d37947e49ea0b47f94573b03553a22d9a1aebeed06e74654acd62b1585331ae5e0e53c6a87f715a1d63f034a6164de89492bc73f4bbd6b6b02dc8bffebbad97d5e531b3e43d6718e42524bb64a172e7f1ed2915074d76c9dc77d12894e61922333cdac45099a6f09c592c7bef4fa1f8b6d25ddd7acebc5bb87817995c36ab8c877f4fdd26853505561e3aa8244803aab4b1e67c19d37d4045548d7aee11046adc6ffb5259c1ad05af52d41b9b269bf060b5eb7a3dfd8f27858ed7a17c15575acd024202afccc6c68b44d06546af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcce969af89c3f1869c6c859f6e63d4fb67ba74b742e7c9367492e901a4fb0f4b32173d994c00ff6e27d58e3403a45d897da185e9ddc959c40a007d22bbee28d1461ab0f5f33c6f6d1e8c6ac889d6ba7e165f701a7923544e6917cfa63ede22035b99ce95e131370a3320c3c4d5c5e2ee03e8359ffc648853f8f46735b7c9eee5e0de493e4ed122d3b40fc4e2e1b0c297f56fc89b40670c7fd9cfe2e9165ce4db498c9329462b352e3abda7a0d8c0b7ac8ca4f52202cbb0404668dd9cce20950edc1956d128a29cd49f2ad4097ff1ffd185fc7aed450f76e27588d5a5274ba746b6dcc8efd6bf8a211f21dfdc00255d1e51f54d45764f5620aafa09658251a1f14a9341e19f48cfde58bfb0f5fba39c11e94a8e55c5bfd18c13fb91553af4d50435ae250cffcb85a6b4dd2868b900470286a197051b09630700eb34aebe39a9552032c53d3c14ac519111ef99eb3aae75f0855c7502f468587a1d5496bf735aa53ff4402e71881ce1bf2bae5e1f501cbc8e7b7dc027dd8fd5c5fc9cdf3da8545a973d9e65f7f16d46c3be7dde039904361099022336ec13ac868b9fd0b3a19b1e4752a0b746fff4ddade3d0eb5f6af57749c433524f913560ff7bef3151bbd04ee40479df8aa4c2775217f4a6a6c0b7a523b7fa074892191be334311e09c730d96fa627ab5df9e49fbd5613d20de2c69bccde8083282bf89d3918ffac7750d238615257da32d0994fba000bb1019f4fd453783bf3eeb6d248a4768df71746b5dbbfa8c41b7ab7149b79ca71527214e523ca7c6e691f8cd6af0b82d0634d99427c6f3b15ca707a3bb3d4079ea4e70a7727fdce2c70c9e16811f78c0e7b445345cbd5bb6da745ae2de55895b5ebf3f3ff5b39bb5e575e0b30b6d748ca0d0526e77f5390efad5fdcd2d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbd61b7d65f81eb45f9562fb7d4d739b064bebaa3f9258f1a97bd1ef742a77fb1ffa9027639c872e0f1e50d22c5e2e03aae16cda140987bb7dabbcdf47029eff18b8528923453f404b500b1fab1ad2484627d2034f053a19526cde5d8c5072d2582602ee64623e2416b90d44d130d60b82969538091db3c12cd8499275eb5e1f9695bca6158b4261fc2f38fd6ad672b5c8163b3df7cccb9a64d99a0d38e45471e8dc8aa996d547532fd046dc697d12003d0ee64364ee16bf2c00b64657c85c21546c53d41e98c29effef90323912724490872d9fee2e3e363ba2d1ce5ac7eca8a31ddc440128fefe48832a2225ab3eac9ef276cb7cd3ab998df09b7b8c65bb5694fbf71617cde3f5e8b278744ee3874c14c4329e086e25ea1005efcfaef948488c945cf9d7e1c812fce7f435eb6f11162c6a61ad7c23fe39d498853f191ddfe2218fc2c2c3f282bc5d8ab6a4579a863911d9a7fc9614f8103aabc81aa377189a4df91d7d9213c59d82a670c8e439332e8278ebcfa7ba6f76b6deca091d6ec88fb8b5da2358901e184a174fb8b32a526e2465e08e7d277dbbefa21d8329f1f3686ea5fda0b26f64a64d3c73cfe9fd6795434eb26be33e091f52dd24fdc2f279624010c227d5c15de8e5420176ba9c160a8ce16158646ff3897314215796a31c18c01a09819b54cf31fcaa05201361db38ff3af60cdc382c8ccbbcb9d1ce9a12a40b2ccbb9bb0b307229b49ebb36bc5f33551546a20e74e37ab443e54529f6653cde5e8c5f9c182068ce61b3c46620879c29aab29343d0eebcf67e8143006be0aacefa3fb10017712b1b20d37ba61d0bc98b40d1171951abb5f469d98474a1072e22aedc90911d43b3b879b4c38aa9d10bf5dc86894b560063446146edc0e31f91e7d50472a51105374;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h61b1e56c1dd7913480d3ee0b5c5116c0e8a86b19195ef8308ebccc63f44a739ae52b86b6498caa8d10e76eec3794bd93b97eef6f119918880dcc09777714721a5ce430575d6a62e04ba036f55ddb6b016d5af649d992f8e6b44f5dcd3367babe69f5e40698a2707f469cd98faf7226bdeb2f9bcaabcd2b2ca089de1a785ddc9d83280020d3b0f26d38b887ee2782ba182fe576614a4feb16a9c1f34dc6ac9299710732e3d7793a142a8de30512217adceb4a7b9e383fd0cd5e8f084d119a1b82621a427b985558b4aa0ecdd93983f7464d80e1cbb62c5fe09afb4f2f8848e36dffafa98ea3ef5d4013a998632cab133880a05700d6fd18bf06562e4d2c645394872e4ebe03f1d4326d4fe59145d220ddda3a04d779caea911fd522a3263e395339b2465b45f84bea269ed858dff5d443aeb3c25d8f3d5948578c042c0606dda794339dd3e326b538873eb494d1cbe48d870ffd0ad1a5175afe0b3c1e998f2ab4c1bb031d1c688319a09cdf16d26afabd508dd00137f7822008133bdf5cae3eac3e0d36d5361603aad477b12b37757734eb2ec83f12793fd81acf0a38a231ad1867d508d5c3130810b8250943b5d376b2d1033e13e35b9d8b518414d607432fd38423b1c03fa5fee7c3b4da150d76b58ee8bfd1bb87a00df9cc8f5634274dd34b5bba1d2e4ac616eeb471682b42de1ad0521864e709995a7c5549f3479618cebb89fbd262853b9553ef6fa9ef8c3b567ab4791d0a4d4ec0525ea1bae25a67763691aa5d0455d498ca6753e5b3cea95f9ddf138377b0418d3bfceff985f137a7d96d3da51900ee15e2e00c09e048678e353d490d63259b63ecc25f7f8364cee2f3f1d1e0e75a1e23128c1e08206d1a5f7c6d547bff4962f04d7f5eb133c2694f40817d75a4059f1dd2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8a834d509fbf6888502333c54d57bee4a85feacbd0c9e69957e02a9d2676fcd8c6cc1625baa8db2e8002609b25507fe74c5bb3c41a5819cc40272cf66016b432c5246f87899ce85f07cf9ec6b88e5c94d7b015aba8dba042d168ef21cb4cf668d7bd93d33ed8f34339e8346d90caf3bb2a11084c518ba331545f0e97c9fd6b8990cd9a678047cbb17306e1d76d3a6d62cb7ce6ee939ae46e23d2cbffaa9f435e154bf91a8fa9612c4bc8917914e7229b8c4b8c7c2acf1617a21390bb8b956e3bfb09e6f481f145e7d81f527fe5ed9414b82887e55ad7201b880eeeb0ea005a45fae76ecd9e8b2ed9e717e9c05ee88c37a877b45679d183b5765fef1b07836de8cad163ea19dcef20269318d312f2e55291bd72b523e0c7cc94df53c7e79471c9ccb840323d228bb18671715ecefa19332df9c91e2d82d57ac2874b90006c0081a42e175d4782c401a9aba2a457300957ac7cc9ed018d767b7dfbd4092736bb9a8d2b38ab5750d67ef354671989f2bafbbb2344941ac3a12b95a9a3faff73d3804c2210945a977e21e9a3a2fedf7c1a17c37bd7356f284c0714e6dbbec30f87aaebb66ac4ec797ad02e689a9eb5e2d71bb9c771a6e6c45f81eea3c41d7a2c4c7a48675cbedc2bcbc4176b2e5ca852648def655c0056a1ef620cb58246310bdd81408ba0665adde378222c50fee7301e9989d53dd092aecd87d720f2febdd3a3052742acc3c62a55e3e4347247fb737b4f0d458aa3d7570ff760aeaf1bde9f78d937b40caf65f607bcec1b450d482faed43f4f6b63941c17a93a03cc2d6e32788f2b7cac78e7a2db30824c8732ebd35e947a4a4b3b35e83da2090d9b5cd3aa8135113b936796085a97902f9f799e19e8f0d3cdd33187d0df890a8223b020b640d09080c07b3323b6fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf97678b49f1a2f1f0dc1322bd6644885fc065c5021c6748f6ca5476b2f5e22ab85a8ec9e6c4b21285cda015997c5bbd18a9f97fb0ccbede010f09a619b76a8bd5323d9ebeda461b18c76ec0bcc6281d96e7b672a7e1007d96605abc3955683dbcb3d52e6bac65fe51c54f253fc5abe6a092d825c52a45e867d305307f55da0b54d129cd6a91938720e3bebf4f8e33b1f7819ff01963f09242811e491698cdc4f1bff6f16761ce45b68b9af5ec24b6a18eaaae5001dc650c36d245bc8bc5e72ae593874f78f954ce268f896742f513c45f5ec1a1a7462865b2b17dd28ab38f77dba2eb02d9bc7a502984fa229d43b8970aa6510e58aebd8f5bacc80efd709a6bc2197fe6014d370ecf00c3189fcb17f971dfe4f5a1d4aeb02ab0b1ea449cf02dadee3c5d062b6ab18730dc36c3232b4d8b4bca75cafb4d70a599c5abaa96fe832a2aca20e45f83ac3c5cd734aab0512f49e1c8ee02af0bc2030491b1d8bf5613498de164747e1454cd5751de2f668bf1812c2cd2b55160a68e08d761bd68a890d8513146856402ca0f693439542b63ef73af287237245f743573fa22b080b4def53fb23c5f8d5af67ad362064d47e817898951c1665393ba6eaa6151931f43d399333594a234cf582528216199c79f0862bd1f21aac5bed5ab507fe899728fecd3c68fdffa233252140784f07bc61fcff250b76d49d3f8038cbe4410395491da619cb6b83ebb9e493baf0b19151949b550c1f48b937ec52028914da77636748190c8b71b6812a2804e9e4ad5b1260f21ea72feca15f60a14f69a0f96292f4708d64d9f839e7c5e3b32b2ba3e990def0d8967bc2871bc28f00dbe911874fefab36d8a203e7c202ae1fd464da350ac9ee2e7c71950309150fa50fcfd810dfe8675d92eb4960d479b3f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd03a91671d861e673095b1d1f31c7763d1236ed7e1594fdd5a4ef46c6a9fb25b325930212aba11d1bd63ef15a6761a2cf3d2f6b61e243c781524e4cc35405afce71c51e87d8aec76287ba2aebda748d6b4c8f8064fa18be91c8308faa5e93ef919758d16aa2c601bd3203f03de97e3745e7771cf558ac7f903729e63c1d807a11ca83a2fffea368336f8b041e496806aea240c501206b8e60741f707ceaa911f9f4e25fc2e7db9cee9c51971d82a5d2c175efaba7f68b4df622dfd24739714c6482601bfee31e8102abc5dfee634a4f95acb900f496d92aa42c5fff20db2508c087ab4f5aa416bb0d12c56a984007ccf2fe5f50fd4a4d41d517e81482f089d80f10eda513697b0208755ec183f969ab993298c36e308e9f76ba5c03c2c0535d030f2aa517a129dd7b5a1bec2688c2fc4307419ad47d1c594da5d1b2d34c084198c220892b7eae19dc0575bcd536bc25bf1966ae3f1de62479111101b9fd9236bfc248f6910d84a0b200f8157b8c0e16599c3e63e9b27887375a2f80ae60f9cfb3be400968cc76f5e3439a198db71ca64250da3a7ce842e04a79bf6091ffedb9a8a8ef00831ea1a690a66a8107beaea9670d76f3893894c36c2cbc845a7aa59d3a176ef6630153bc20b62ab055b02c0fc7468be0a28e1df4fce34b63c51568d195d0f654270d5bfd0c8cef0f15ea5dfd9dac457a9f381604ff43e9e09b50bc431a03fd97c151849539b559022acde7ef4ca796b8ff166ed9284bf6204ef2f852727773dbe5065ef4d695c2eafb52d43f7cd6660be27ab5de7a2033c1aa7e9f9b0feff8a46df0c3c43f51e97d9645989def89a77a92057707e4140f2146e814b5805079cdcddb6491b0c16f67755f1499223d7488faa4ab67531775d7f83094fe21620bfa3e514aa49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha8fddbb5d898a4d575cf809f03c78a8db9e61940aa47e542ebae7e6642edcbf4ea6274e3cf5c348cd7c92982a6468c53e2cde3da0e3fa896ee5fa1f06d08be076fdb9923adf2e83415e5183ce768b591e3f83a08ff320e8ecbbf85d1a081bb8ad7e1d110b7ab8fa041bc0a9feeaf052736f99276ae52eee764f1073ed81e8ce9bbf1d5797648c0ed04e23e143f24f597f715452c088ebd781406bf1945326d03d221a3983476e2df1cd91a48af0fdbad12bdc0c47525eae3d1929acef7f0afc2f0cbadbb54c8e4f32669e78657c04e2378225feb21eacbb9a437671e5db5377c0fbbda56d06df2770fd2c15097d51a99b4aa8df7ddf2966fd9fef679d64de8007efd1e79c15b73c642e11bcda08e297746435598971f4bdd3be66ffed22a173505e74a7974ce42883989e57be599a1ad3e102a912486b85b3213af0e061af6e16152cdf7f4944730c2df4e951492656453db4006aea674f952dcd5a7c9c079c52e03cbdd60fe15dd5d6234aa4ffbf9b5e6d654c9df52e1c9efc6b1341bf3737423fe3709310a676b9d06d7fcff4e6b58a427d9f744df29b79d2087570794578b3271ec3da0f5098e9a24663f960fb150852ca9abbc9325ada44778c09d6379208364eefd2472bc2c6467bf692304f46587133dfeb2e8d39c5026c4093d8eb146e859b9d1db336e1fe1220c68c14d4d1e50ede525db82dfc4e48a96894c6c89dedc24d81273bdc19789227389c79f38f0b08b4c95724ee13048d5be78804b02304daa36eb8b467dad2d946aa7a6584de416f89eea0faf9bb6e7e0da750e7e9549a426e45b35fcdd34b49042d53c2d6fb0f1a24f6a7a9fe70d54ef1545cb91dade33417e296a8418750335a0ba9caf6fc7eee4a0946998b61be784af98b6e006973c6312edc46ad705;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha2f790f73700e5d12f6a5ff74fbc15946f809b1a7e9e6001019179082fb69e2908a493b538207b4aa136c0905c2b0a13b427760d28cf06210b7c095cb51c31d076c9d78c15f39412d1da69ed776130c72e41afcf0668644ca7f273098575c630f173bbcdff853f10cd56427eb406a11008b098ddfeb69bb02558dd023b1395e1c7f703c6e707643b643956b9bedce4782698277635d2377e7093f2bd8eb4b6ac0a6ed1facf9d7b326850e7509287bd3f38ca92cb46c6894d2ae5cb6fa31b53e2a78ccdbf05ec44bc158f322872198779e6a4c044b9ce826bc78d3bba2b4811d7a481878ba670cc4fc688a9538958fa7484ac9addcdfb85dac575f2fc2d0d04ece7e8070afe712fbda415a0383002bbdc9db98df44fbdf34940bf4e79b1693dae1a1173768089f85c6211f97dc683667f1a03d978d7d246db8a9a54eebe956c73abb79478bad18bf701debc5701c08f7c3ed9768dadb1e6f7c34a4c07d7e63627aff0272b667f9a75dd2f51f2076fb255ba8dc75d51fa4beba5718e8559cff2979cef4757a395c9c20fb37d505dc49e04d3f3b16d7b5636d5f92d1fd1e851dc580341773a2f87b60b1e078885f080693116f250cb586b1d09b080c3f02b6d873a0b1d2b0a9137cf81a08b11ec08f143c722b6edd9665d6ca22b3f2a5e94ed0bbe40828ed4bf8bff9ae73d77575b1f499a72476b156250c7fc652fb742055b4bbbb69437555a47ae55ebb51f18aa52ec8486631de41f32a2389513edbd980c881b0a1ffa3384089750cc8ac0abf080dfeaf6ca39fd9d193380b00f24059aeed42eaf5659a5f1af112e2eb1b53c84c8d515a66475a5223d3accbcbd4a44f1d9ca795ae81af3e7b42b120796209c3ac563b840ffa4b80ee81c8aaecc6d3d469bf77850c39856dc19cdb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5f97950143cfa41277a042337600c46b9fa0c549690ce052b324c96b303a4aba9af8c42538a900a731cbdc86106968e0269f90751075e8f7dc9f39f13a58ebf0970dae5b03666af0bbb68aad7e7f05729fd13bd9bee0125bd180dbfd8039540ca9b68e0a8984aa4618bac1e4db8e50be004ee98d3dccc8a39579d73e36248bd244a3a97a81fab685e046f5842eaaa1d92571c5e37c36f9b9a6d77f429abb52daf5b268e74f54ee8230a632e1e3c34c5bb8d08de85d9c1d17b5562668a1138f0edc4cbd72eab6ed9ab9d25f9b05cbd696f931af245aa5a9e8770afcf6ec0d24fe2a662a2b3272b6495cf047ddba25fe550d9b101544b372c64cfb7b01fba1229306eea6ad5e68de23cc0c3d9b93606e8d76312e17520e3eff41750a8cae2f56ac8b613bdb6fa1a206e0cf8da6c693adbb60c88dabbe63669310ecf1d445ed11e079c8152b234e5da77e0b457ac41546eb793d2372456ea3c4262d439f24b9b773e409f3fdac6c7cca979b30d6eb5ce314198f18ed1eefe9e83ec58cf7a46be2776d09c28e8437acf3a3b5d7c2cd1aa314a5d3083d59fa95c37402dee5a895c0d7b9f1ae4915a0eb76b0148059c805f35992e00f255f5da0a30257e8b210b8cbcb3c2e7bc0f39bda194ac1d50775ffeeb9b4100c9eeeaab86c64e29a993b2917aa2562c293c020ca41e5ced4bfc4a22e2def82e385d822ca384fa5d6110a72084912669133b667ba119615abfc7f8cd06950cc1a9ea4e562f21ae74610d500453510c400184466e96cc9bb92aa02478dedd9d0c460f88a50a8114e85ca60e962c9d0d6f299290345f9eb1f117a7ac00eec14279934bc77bbb9260b88deaf1001a5d3e8cb011fbab9a1f3f776d70394d7ccf85b280b56be5ff26187d03b1360b6feea5c42d9bd465743;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h550301f4f73d70f783e9b5bf5193eaaba26345f2eff61d352f2f92592902c54c13ee042eb79054151a46ffe7a633918ed310400330074f5658f23e7ca5bf46ba51c535b3f3282d862b3e91186adc54bd33558332f535f0694f6f1eab0e80acc16b3f544888fd85698302f7869bd87659c12ce95c162f50b6cacc4d152091352334e9e702abd2f06ac213676b7fdfec8f858cb0b525dda0c22283f6fec8ba2e76546b0f7070d63aaf9284391b62f626e64245343f18be4f2080c6af21d484fcc07669e921b442c656c1c9c62f6b2079169acca4a5a63b7194a051f6bfff4df3eaeceee936f68e22d809ac91be3184a1ea5af233e69a0273a39d0a5b352b60656021babb8c806afb452352d6cb933c4c2bf20b9b4a5f4e8e6e3c1357e7de2c2d0ccb98f95a25e51e2c65bab631c56b8f5df3d8b36956567192a8e3e673ab1fef3ba9f575b26746588192beefba9bd8fc3359bacd26210f8eb8bcd3f9a07b11ad637370525b3f782e9295df20a29d9b1c4e16a986697377234ff3ae77e80784a8e20f63d00af2457e2374f100eca8ca76d9b361a20c4bce9c463df8e134e4693a84d8c5714fb56820ea5e6823fd2044a95843c1640e1fcecddf0ae8b387464c7cf29738cdd1828c4e19b4c95bd7902630b5e06f7a7a021216cb95ebe08447e703c0048201939ded08ffd727a559b65c52cdb1fa1cb5554cb37da8fd8f8a65c46b76160b50e959160273e2d8db606b936e71702d2efb2b75ede2e8ae785c9be8e84ffd166e7200737a779267078d99e74f91d788d8ee5153976c0f954df84f4f388b67806f0e37b5fd295fbdf412b8a485e05f704b9246ee2854e45ab46e6f2d92ff87a41b77fca856d568f91b01ff167cd108c284157bd0c0bb0b0d2236ef2a6b4bcebf23a003bc28ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h428c4448deef9990c01e48b4c707c255c1aa2b4b50a3045b1f80ac54a345e1bd0d6f964947a63961d5759801f43c9c06aaa1b7085d2a0b0243dbf6d1da414f3187945b03c1c9be43371bb574a555d18694b943faca9594c74b523010bbd5babd3b063ce3508fad0d84b30a824a59c856e5c2520c98ae56b384ad8c2550d8e9674aa0c80dfe111f69233121ba08a4522c2288acb9eeb93bedfa17bbb06913bbc877dd105dce5e86bc8114f3be16abfe208d9af90eeed603093519a6db197570585d8f3aa7680d77ae45a76b33b3aff79e203e27a2aa4f38873e9aee441a824e0727718416a1b455a4f8a0a8e8de191da40d8848af34a12cf06fe3b58fe0807025a062ea47fb6a9d35d08a4ec6021ffa307f2a12d2589f96d9a6f5a322a416bdc6319360d5f0720bb12accf891021ea7f22b772b4240e1f8291e186b5a54e744c8e52a937eb1d0adaf60da0e57e17106692e588a59b295bd55e0be352c05ee0958385ecb13e10423cc14ff5e84474c1639592ab6e1f315dd27a861fdc6332e846f3e5d963b4f338b0933187cfa6bdb2c95ab8e2a1b52ec591928ed6c0b1c216d195720ffcecedc6bcf46bedf20cf704e8221d295ae04184411f26558109fc73497070afe3cfa716adffcb910660e329369bb57f05d121dabdb1b5fe930211feb1ef61647d62e9e96da0af4b9a8bd9059f582e7c8192d1a771fc5e7175de3362ed8d938e432d5b86e333af06da06c2f349592d5aac3482a66f5e49a46fe4c3070f79d91aa7895368f0b481f393df8f11e1cbe73cb7b95d7c1687d6f321e7087e32c7fc9a5403be407e8fb39fe87b910000fba1174577f1d521cf5b345c1c6d3a45fcb03bb089f72f0b3e0eaed8faf7f5c5f4f629890e5dccefe51afd3361f6f0f52c3e539033136ccec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h26f58ae6b771790cd568e3dc798b43e85631390227ac0b74622719c52d4035a1f30cc9ff8d6d384648bcf80a8960811a227d4dc40e9bdbef3b7dc0305fce5d7e45501e080146111b47e67cf8cace6be32ec7b8753d8b827728850811054553ada8d981b47846d2a89926b16183bc6219ce24fff6ea5ee2a3b4e6c9fb21f9c46accc77b408e01cf5f9692acbc04d39eb3a80cf71b0c60bd61421cf9572ddcfbfe1d9abb1f0f4d50e27f6662809eea439ad98bbb3f1336341edc4d52f33f4b966a1c3687bdba8fdc3a4174c672aa296e92522f988e0e24711fff56f30853c7ebe9229a652a0f5b56b9c3898ae303e144d4e273ff061c239ecf425fc3e2df3ea79632b34be97f75eaea63c105dd479401b9564b9cdf6850520ef57d19625c8e62bc319fe02ac6a07fac1089b7a1c94866e235fa0e79fb0fcc8acfb019bbb7577fb2ed12848be07bf57f82fefc859095a271524e810aaf33eaddf13051a0b80af11cf77dac0f8115d29499140ade164291f0b5701adb9bfeebbf044171d93fb0a247bb628018ed9441a1d3aa8df1a7bf744c29f211f407eafc4f343ac858d39c4a899c4d6dd81fff6a42041295c203bae81957e2a59b7f05d38f1ba8e453cfbf41b5cef75c038ac1eb609869523bc46b67af99a89524f9e4aa56d6434ae42c1b26bb4b4baf1592e542a7b25f767c1abda6b254200fb209b2a43ef1f25c1ee71c1080144982105b992786ec63fa8999c6726e3789f23e741f3d521913e159893f330448b4ae631f6ecb2bfb24b72c13cc5a1494f0c4a4792668594faa88ba278a35f600b4fae559ee81a9ae2a27e6b9c8dd58e679f44ce1831358ee92d01de79d3aa6765a1b71655b760bf7f47bdb31419913af2b6b1e85f8ce061949986f74a3a3f5879b2467a11afac5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h29684736853a5fffeab31e82bcf9309608dea988292758249849aad5e089ac561b85d31330679d5b4b6ff85110fe7cc32a15a0592a007c196ed21f471c22017d5d4ddf6ac94d753676c987e5f51f326ec05f9e56383b3c1e60753a27efa6cfd3d2519438043de5864fb9409aa57f87423d1fbdd87c5d3d5a95057591ebb668f88031f621c8d52407cddf0baafc54270416e321963da1246da8bc7d8fb7e917458280059604c6591303f120d415a11a48009900368c95c9fc3b861a9c7d1f7c32e75fabed0d64d6d44972aff359b686bf94196ccb8d098fcc9872af58b403696c7503fd70a7be6b623d1cb788c8bd64c40f34993d67a03767883e5b318674b217c7b5b3c2d9bc7242e0345360e82661c3a9a6ea6ad3adb688f8acb31941eafa11fda33c6a44230443a5e78d8e4859bc81d1a89bc1b11f4fcd77c6b8a609064e7450170ade4082bc4e9f9916f1a4d2df9f4ee2cb9f7318dd97ce2d847e39cb7829736bcbde581d92e20037741ac40f8d416b21b8f050c8ead3e5b7014de9a7e2740953b8c57d0b55e736887587e7d476692a68e335fc1e18cb3d42b22a59549c6fedb22acab31c0e8bc2252fdc9ac1f5dee65d4f59ed64ecb83eea89a3e710d0d374fd69c171ddff253c46bdff65cdfa8517110e906339c95c188183b4484d98e23e2eeddf1d8375ba0bf3a81b249b8c408622a62513054470c66fa66c477babb6b7e6bd7e25b303a0bf91f6c4e521b700f91de5bc07aee1fb91b147fa96b0a2946f92671c2dc97891cc300d397d4a560a55e3ecfc6db149fe28278405e6d57ac4f369d9c63c3b0a3f60a4b18cfd010e889e1847c13587fa417ba7f8ee2a58588d1c764f6e37bfc73f25d08f7f14ef9f83d1df6b15d812742d3213662ed884bbba2b5a77aeaf9db69c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9756ec16ded01ea43644303b5cc1dd1098f8ea694f4adce80bd3b13c85a41c4ccf18026fc3c3bb7de9caba15592a0d5c898388e66dcd5f1c5927dffee561520998e258bc74b4f63f8682a453c68ad57e749537d1dd0f2dd2913e861e0daa9bfc1d8e93c0540815e3362c54a81f0cd391f0a85358cf3454ec1aee290b03b8a7f3ec8c3bfc9d6a25f8069fef51d8f2d739be0a6dcace8e4efe1389abe9dfe7ffceac48c8fd4d21966aaeacc6b8f0717f1d8c3a9194e38b35e091c26a994c03d64e10848e9bb22449c10831bc2169aa4125741cbf61263fee69cc568a8fd456cc061c3d6b44602453733f392f3e69b9f9e335982e6912c0eb9fa9ac6dd29f77061dac8990266218b8988db3949cdec2a7cb44b1803ab9d141b18f8f17ee6c99ac4c819d573bf7473f0d2d789f320fd92f136836e488843474b287d5479445786ba21d10d5c2395e546fc78bc0fd985e3b1e7c818e7c0e67101f5a680d081f7b8e756e9b2f8768ec49885142abb8294f4e5bad9eed2ccccdd191961f352b73b82fe70f3dc3b0141cedbf52ae28203bd0f882753474ed1e2367ef52a33bdc3a53111d21f2e6769cf7af34b3c2afbb24e24b9e062407449c196f311d95a472e16bbe13caec12bdf41bcf918d06d5dc2a3940b065ffb1c0737e4310c3549d2185e3c54192a1d33145e12b4afe2fecf2aa40dcbfcfb050ccd8cbf4362154cc8637dfc0015f9322f67d46f030926455d4d74d54c0f238c883560606286792692764a1ec5599155a20f9f061a9016189ffa9ab168728e77d7b0329c8f3ed5d4338146b0847f8d05f4162724812f26f350541b23cd5d4d7dfeeaf5e04728cebfde3ff179162c5d00e372355ea86e0aacf19528ce9de400514f787193f5b066531132920b4a4878b7b84b94da158;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha132d0cf34c88000501d3919f56c2211f9b767806e4442e7fefb1f7f09968a073379b763519ad8f96e28c28248fa01b2cd3707b74d37a2ae77303c8d27a07fc1fc5801455b1f68564ed02d51b0e326963ebd6129a8bf83c83bcf5542bfb18dfbc89f31117ca553fda02f5563b91203cdf9d97789e3fbe8e99a051cb121dedeae3ba48715935ba9be0eb45e960d07cded4fadc7fd91ef1f5c68ca010227ce95d4cb4b3955fcb511f42f4a43f44dee8b0ed63ec7d29bb86a2a50d88930e7384f5e8c10ebab04f5a089eb2c07e7cb2158949ca280fa233546933a6fe331fd49273cd410cab457974769c24b2aee39e2ba19ba659218421763da09754fb8fd9feee3325fe58e9be96a1f91ff309a716407d941bf80edf60d1536ba4d6c050a7fc2dffe82de80db10c96c432a7d7ab5bf54456f54f6d5df55180e4af7400d19f177c559a8e7e57151c7058a5a724b80a8d1aba0f23a3d2a234601c19c5553e3c8387c990151db31354ff13751cb42ca1df048e14639e5d8c57c436486f4d506cebb2db4cc52879cc13ffefc53fd9e795593b6c8f9162e455b5a2993f6bc8a2c570472f50a949cdd80bbe135409c2590aef2b75f3fa77c8cca44ebddc58ee940e08994fb302f46a820ea9504eb66fe4fc0bd88a1ff968237c0616ccc21a5ee3bde41ab37ed449e95205fe7cbfb9bfcfb2c00088d31aa97c91311afa7f28f8a398e89e2db60b76464e9a0df0835cb00a5cc950fd9c3b10a41a3897f162c2da688f8b5debe4e6fb92a1cb2037f3fb7721d1d453c08735f4424bb2b7926d18c7526501b695305af2a4b381cbe2ba93e789a231a8157d890de66bfade9634ebbff13c3a0be5bfd85793d148f18b000620032e6a3d26d2fa2c58cb5efdc5866181cc7c60ac6a848f6d25d33b4c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he359b240d70c1878bde7acf6ae5f0c6ea451c51679748cf248159650c9fd0bc103be616f01b3cc9359af7495f30bfddaa6e6f200375d4a9a810d8fb4649671971839539bba3cf4b9ead824e5eedb117d2bff99e742534b6e153dfdc62cf60e310d7b9a6b355282c834903a3c8ad0b7c8e3ddead7c4ca5787e6eb662bdb048f6eb55377becff0b799d75a07c318fed54254075cb523f060550cfc2e6fe20be5e8e33d8722df4fe531316073b6f058f0a0f93d0f350c8f6f7eb736202b9b664d364b4dc2b6af7da6a8044b73029e898c3f237c73d4f6f00bd35c1914d50cd4b3b12941864cf782d0762ae8c233d050ee148e11b19441cb851044a2a77283d3ac2ad1c1b6cb8709e105d3cfb90edf49d8486baac8fd65ad6ce8d27a0fb3ab10111a40a7c02840de3ec6cb96ff6979620def0cd060bd90c31535cbfc5b854d777b39e0a105ee221317cf451012a09581f9edb7680e4e1adb6eec30cde3c539f6f475266135ab6f6440b3a8f74a988c29ff8f113b37a777784e4ac2c62918ce0856cefb9c3cfd890801556ee3443b03b0a33976bc2c517fd4df2f2489d8c80462fce42cab8362662afc97372c0effba9154316f0817da3ea8df43cfdafe1bcb8fc64fef0757520e5eb3b756b36859503d8d5ec9d6f15a1198bc532ef198e5ec46016eaa673a409dd45046b43592fd3c0d51e5894deeb38512c147d1a3155b6eeeb2cbbdbd05b27fea23b470c78338e8cd6df20bf5f2f2a935daa5b5c71f068696957a157427a63b0aae58e150df6ba1ee58ab1f1ec4bd3e57ac9d7980a1dcd96604f633ce01d322fd40dcacd6088bb5697771906176ed6530b62f2ccc934b93e9d232e77a237b895b9cc29146f4ee780d3f1e7075ee094a7d3111da4f13ce60f58f45fcff801409c6c2e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h906d89bf8402b151ce21bbc0333b836bce4ed2f7100199f583e47a44601fb559bd74b8f09e76cffa1e77982b1b5c8829e24624c11225c166b42448e348a4b5f14b935a1c08a21a70c5524be52a5dd88e15097ae81d24eb0dc29d7eab0f81a2a3a06c009af19cee36e22b81c5e136f980a71c26695d4881bbf13e46def1301a3c0d6fef0684741712bb3ce8aade8d6963b27c043c7d3bb23cbf64c012c778bdabcd547a829e2c761e310c2e96ed0ce06da4a11d8f36a30930442ab7ac06433ec8b0a7c7fed6708646abb9e70b357ba2e1495cf6d02fbc59b057e2a93ad01d0acb4190f6160b7d8f9f4b52a588d1e4a5089307ea9a6f8f1e7378dd35d36778ee794e7a0d9083e7b001a8e44b9515333c65471b20d311d2a84016afbc772d080784b947ec510d48ac122b5c87b108d05ff9e397495b6cb684107604198a22e027a260f6d179e3de847d5451dbf328ce0f0712d79faa568450a5fcfa82d2fdeb5234b0d549523460eb816e24681ace4d7f270787408322f0b8541f130c56e681228ecb3258057f9503760dd5ac943c1c39bdc7121d2e4f4c5b87d8ea79ab52ea9f09310fab5ae1fb3300d832b935861c3c9db436ed57515ece28762fa6a5aea6ab3d41c916f5f06b73e0f643da8fcce3c5c4430edf5045a7eb4edbedf971f04aeac0c796de38fbdbcc39277487f0d3bf36928c2a9831f680fa3bee4141501d12ef7cdf4c27c991f2c44657397b1c03f6415067e39159df6ee341c64d37238c46c4a0840ff861a97929a646001770ad32768a1935939a54addfd08ae72a3246188c36f8e030d11049fffc03a6a38971e1bcc35b15d2fbcf79d18426eb2ff4644c37dd65d6ebc63157480a031cc62aaa6bd62470427fc5eaf7757ddb7b7250f19fa713d55c066dade58c88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4c75827c9a97a42f1d4ddc7c308e8b5180422901676a63db587a907912eafa437ecdf4bf30e2d65bb8a934fb99b402cf7653ad7a92ed3c66247797fabf2f99a0e80efcb7467b14ec663fd82d56e11de5ecfee414388d19352db2390be357279a438b775097a1b6f601dc1a0614b4ef5bc4d249aba90818cd07c4cad243327ec6b605d3878595195539766eb9ae3e22e48d2b1de05d96f0e17ad8a89dc163cc99171c3701f61d64deb65abde8178b704ab1e09552182cf623e40a2f710dc34890b37a538f33c4b8f61f18655eaaceb993012e0afe93f4a1831fe31f0c6b73531616b7f78aa9d4628df21d4de7d20e0e4e54c7f7df9fc2ec30d69a520f3d703253070675a609d69e8be6972106fdfa0c39cdf66b4050f5bca61d1cc5713ec2f0373221080f8cff4c5abf2214823cee2a1fe1e8748ce7bab72537c63ebbe22ef7334fda05bd0bf5eb44d1df078c42be39c51039ec300c0b4544d9e81b2c847c69a36fa4421c940a248b3f2acffa31dddee862573b7085dffd644616ef30ab089caf27f3514cf8cc19458a87853a294e5729b1c9a1efde7a629e86aa2a1da6dc8a25b344b41bc522e7934bdd5991e7032a12ae3ebb706a9a9ce0f99320dfb302a3e0ef928d6c14c41311e56f7677577aed52b7fa05a9a94e0daf6d6899c19180171369efa723fa517971a718627bcebd6f3dbafc1fba8eed63b73f4a01d2751846d2f3e04d3fb63598192e0e69dd2b4b7f4a1b69614b3997a451dc7a0eebf55935cc522ba3e5b1f2a2973d4e267513d03a45148c83ee21fa4d66f85a834fa78d98fc83d13d88ded2393c414b407e0d40fcb8f624ba6798b243c7eb428efb3590d03e00d1caf61eccd653d16c82657649321146eea5e6f7946d55d64f26c405fa972beb93642f229d2e2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he04d5c5fa39cfceb252aff5459ce3d548bee6581d9c848884e299f7bf9c75df7bb45a42894c0e60768cca3638c680bf67240c22e7fa4c3efff09630f969d91948001d786981b53a0c2845dec1e684d07a3e3c9fc7a0b35471f6fc70fabd39ab0dd716e50c395abfc101b100a17ca9b7b54742861b6db05332345b19fea588a9f57a3e3580cdfbbe0317e1ad7b8363849ab6fd565e5e9548f5e5ae7475afc9ebcb2205b46c87d7d2e896ca74e5eeb59586e743e343f50ec78fdbf0280e15bdbd7c9064e0f422fc7d0551fc135bb09d2feadd67c8f3520f28b41d27bd406e8e0f71e590875cac3e99f82bf3cac603815302603ea5f36a6af123213c0f4f38c761d484db866361b1ddc9ea0f5445a343d51975cfffa142f34fb451796b78fa128e69415c61fbc323884f3449ee138b95c9a72364a9a1e91800723e8cbbe5dde29373ab9b895bbabeacb64fb4195bfc52bf8f110a4c2c06015394de07bcdf03317d531feafd8ca92127a988afdd108b121a759c4e60c4626f2f9928c161eba9f5690998a87951121a4d4e798eceefb56ed7b5de98b5602d28088c2f54d7ef565df5fc457471ccc871aa5b175ae82b039e310e5a656565a0c52086a77df58a70c257c3cb42f4413836265706d3190d1d057e155428f5d5768cf5242cbcdaa1a26d0e6158e9cf7fe80d6a70240efab6cceae93c480fe30c0397505ecd87d088633415db22e93e5272f65851bb3062422ee66c84b54896e53edd871135d869a59aefd00bd3659813dcc2a2dc70e1871fe8f51deb040b07dc24a9726c3399c86cb5dfda3706a7f8656cec3c4e053c64ab7d9d209edb5d7d11530a0e23551dd440f238be5e1fbb60de1a7bc355661488d213789edbfc956130e80fb0ffadb1d5bd6e89d3f135cd1ab28c563b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h164e95d3330aa2fcbf9e9a32a7e149d9465fed7dcec680ebf30b9f31cf4668c42df17fc82cf89ca5851a3690fce850e7ecaa11e0c149a0cc1b725830abeac82450b1ef58d86bd5b71e3a429910314b0c266c34e039f98930d30cdd2e83c3365c95405c668df480e9a29d69c964958aa364763f9fed2fc8d9ea94313ba76e8515df39d62c994af1645f533fb9f48ae22d4ee8010ed8fe7e16f6016f2f3992f906a8e8c3c928c19b9bf299eef19af853d06138b7f1070cf98f59bcc2764c985e27f73f1591cac95f5536e4c93d100ec4656ac0e7ed1409a53958a4ee08c171a0ea50bb1160bdd697bcc3165278dc547c60bb624e30d1126a5d73a0cdb6f88be9ab118dc8637687ec7ad22d7565094dbad5bf14489801ceb11683d1f670e0d71256bc83cd7422920429c0881dbf52daab1a5169df755236a588e6185a93a2ac88d037447a81cb7e4c15a37e477852a610b26f61a65df72e86af34298a48e6a6a49869434d207cb75d49ef4ca6f66cacd5241dd2c1bb506a8911a28679d496287d90a519a3c487b6f2cc4bf1f1ef4d46cdfa5ea22eae904ad0f78eb6a182bff1d5704b17cee4f40259a921eb3a8660683809a32e9336f5fa76c6e380ad498e3bda5cf567ebc0b071321e38a581aa285e70e41af25e95d76abc74db432506c9ddf4359c94a953c3013fbe8d80e4a81850dec888eb4edd09839f3e9d14aebdedae73793e4dfb1b5be3b7e8b1bcddb2bf6a5af8b8e8095d58016be7a9678fe98de2f5aec989abe90ae1b3e8165fba8c33d043467ae904cabf797a696a86c1a83f28ee11dcb2d02cc906fc028a5dea2c54cc07546c0f3561b1addca43b1872b574d3ed275821927c1b451c48361daef7a4f1f1b3887c838e2eb219865ef7dfe89385a2b8280266e7ba23195d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf3b3c2b75c187d4f0eca7da38d8ecd8fbae7f320a6f42d227fb5754341b349f22c9ccc581d95f453d2bd606e030dbc1c3ed7df61595af425b98fe0d3f0c30fe611f699eddc6aa858662d6cd662200bf154e9295ef66ef13b7582ae6d9da2db1c6b6d527d68982b06d82cf30cbaccf9f08e233e1d0f682e21018a659b817a295a92bab1158e9e4507cf5918ccf9829a3887417beac01f7064a1ba2af9021cb66a622a2b334af297e267b2b23efa98c80680dead76b8effe90c0eeaee22673ad563e9fbd191f7bcbc043ae5163c4c9be7bae1d5880a2dcab09b5feb2a62bb2289fb82e1d8ffd9f0996006ddf54074f0117cb37bce67265aa0d6f47d778e2b479cd408898df078417248c61154e997620aa8fcbeab5b869ae572d677605b5bd7b4fd77babc82e7baedb4079df11f79e90e57d3d0d86fbddf5e1e81d9acd0317211b04ea32e365a90a7ac55d339a2e157dd1dbcb19bc9988d337cc438256bac53e121e1a5a9d67efcb95bae14d61260caa9816000e1f866fe50b6b5c74344abbc52f222e0c0f21c0ebb2811d7e12925229a8a210922750f43995e3ee0b151af856c081185370bb6a76d936abbd89384b1b8d1b2d4177bff38cddde9a6c2615d1263a634fb766c09f39af52e00301e2f0a3314a12f12a967d6f03f8b4c5f286d6fe1f660b6b1e0a3cc35ffda7770e50998baaa6eafc98baa6ef13fa324113b987558cededb301014150927a7f75cd3687f5142af870fe3aa578cc274085c930ed9e8562407fdc513715d2362d2237b310ca8f2b1bc29fc24940f9f506cc2641df0a39695e51411a59946fb0d3b1a921eede547eeed86e1c2fba3665e6c9d6a752b22b06196a275590c88ab4704c3500799ca48408e8593f10bb689bbbf8d46805d4269a8c59216d4b5879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h220f0cda436ffa86891391bcf58f34f1e5763210eea895614330221d7ec3267d611ad87054cf406556708a3d735931134fd03565ea1d36fdc57752714604b8424b919b638e626b9e4afa34e7e41acff834540d72133e7ac3e66b50ade654351f6e9fb88c89493a8e676881dcea34e33e69cf43d3e83bdc6b40f91196558f7386843d5bf9295fa5a4ffe9eecb090b97acf122e5c0300faeb764d540d1076850ca7f7d385e6c61664f427c4413aa24094157f8d5d3bc5546617f3f672f85a4bc5859c6c8ebc8ef2d4a61e21a2269d7e3184da68ce93d65b07c21822621dd8d92db336a67bec01a0a912287857cd943b9dcca8cd8bbb28e7631dcf61172ad97a8ebbb397ad2d53422b4af6a416331e58165c361d2f803f688af1d32a10638cfb02b5ed482f265ba7f5dd930ef8f5b859698e53e9c79380a0a2a03b0494d0024a752760ab571979b943bf78e39cb6ee43310ef487e35faa5e7fc759374c2d242e997639d8ca400c9316f75ffd2c605efbcb1d9d84310d3ea5041b31a73c57b0bc1d09a1db5ae258279d61263049d0b97045d5d4a3d73ac9121b46573cd3e1336f62908343c7abc993acb204d585c13803abfb17603deefc363a14d82b99bc2e90f718d48c790690b57ad244676691fc20ca83b26bf1515da928c65bd1969bc0fe6264488e78744f8f429082d91aea791bb41c326f3558877f0746beee28e3863692e92f203ea98912b522f95154a3167f70a49aef664fa1a4dfcf66707ae17acb482b993c00fc654d9af74b7ee8e2c9f44535de884df8b6f00ee72c885b7b0019205ca9221344d0980108726689ecc8e8a6280a25c6f54b6744ab56e84d4e8086f0a4912b82ca54ffbb7e71a61cb8d24fa679dc00052e6c78d75a0f864696b6ee869c4444f1c66415cd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd886a2cbe05de2945f93d9288407e6432ebeee9cd8703465387c86354aab94521d7df69272ae0e96d82dbfe7166bd9dc49eb44b8b647f9ddcd585be482c2993df0f33484db874240e232678a399855acd0f459012f862cfb89a049923b99be8ffbd385c0169c052a2994eb1e97b8372dbb93e2e6fca000606d8af4c315e7eb621189e82e810c211e1e2ff850a6a32274c416b567c2e15e2831599b0474b74522cbb04011a94d1f7d2a8ca1e8f9d70b7fee59d715d81dbc51c2a443647cb1ffe4f96c1748db290d913e61deff3fe33654b6428a003d0c363e23d4cebc5071b6cccfd293619f07653a40207ef6fb457758f16025361e594e539d4e2a063cc35224e59ea2a35b54480d5072bfc388be41fa4fd11776fa7a72a0767a435d16005be552aaaaa54124b86c863c0d592d10a8e188b826239ed6537b260fba84ff62a8da2e2848df2cfe3e3cccbbfcaccb206256d4ad10fbc1d072d072e2e0a4c3fba3de8251024d1d52ac2dc8ff18bd2b09ba270efc5e13aead9451fb7b6cdc7e8c5d617ebc29998427778230823b5741c94be8faa188371be4cd51df9b48d9676a80ddc3849f93139b2376b368c634572a1f931c5bdc9438d5470109789b0269993bc012ae29f3da466296d202dda0d14a6ba9a9595beecbbd521297193bc2658a270dc928c5a11e27f74dccb7bf3bee8ec7bc5b04f6427a0ab4bc4022847e4ee87ca8f30e25185cf42477c9a175b4427ac0f0bd8cd30bce93c7c7c3f4fa867e511a6a022c4e2efed58a5ef2acfce5346fb21998e8c47c19db73dbad118172790e49cd4f69171a9cd9bbaa0d47880188e4317fd0511369c447ba170c7afa2ebd7f6aeb5203ad251b36b4328bdfe8722648e60400e409437cab038d10ed8cc8f046d8981003efc719642121;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9411c7db87b45392612d7d4c0c7afd53d24fe08c515ca5a38459bab37fe5d2fa7487bcb2b8a9ec96db82b0a19722c34369bbdd2b2079a0ccbe9c0049a8774531b209563fd3bfd8e34fd68129be72d664eae4b51b50a4ac413c9c65153b4819de25331e1d3529b022f75159bd23c29c050405f341c1dac2e3d6f1c4be38bac99e8a87505ed39d8b25b8654c40236c470bb497c268424a6ea71d0485bb6717dd201227507b80c7f4b789050b78377242b038c99bad75e6a290a0cbf9f146269836f894cf8cdc3bc8317d77245c61192587362b7d036a8652962feba214cfe02385391611f0b4a1daa9fc7e3edcd2207f3962b4abc1a425d3aa2cdfe9d108c44bae3cb0ccd02b386ce5d10dc5b67a4cfd535e7a57fd2bf06f0fd4674c8b869de9108d22a62ba57459fd5f29026c8363d22440275817e0f3179443fee03a762a3cd3bf30a40e5f1d31ba25870e3f83289e7b8e69a29fd08917966231562f25b9324b2a6bc60d238dcc049d7c01931bb6b9404861841de76e9fa2dd8e6d34c37e9e56ed1c147f5e8a5acdcbc4c05a4835cf1c25204c61dee685f12c90c24b593b609f58edb9c50dd6ea94c8bbc0a9bd914e5146eaa50e1f52b841849de863e93c2d700ef5d688993eb2e798c8a39572d10262a30b626203b637ebf56a5032c4151f2593e11497ba1a9cb78f2a4cec88247935bdd4c3608d978687aa6055cf1bbb60841da717890bf66d8ab796cc91ce75aa6a924c9e3338ded0ad195d5c07151ed3784cc06333d2d1884da593247ebd97764b2302761246a1c9ad8b9301ef1987e6129f906b18258baf7c12c8d439efd3f4366288262553ca0fbb988b5cf64791d4b5c61812c9d1c3a54fd2232a976586c593e14999ee15096a6dc9ee5d17902fd759fa8aa6e40e95d4aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1d3ce924a670480b5f5bea06314e289bf463ae511b57aa26ab3df7f8695ac3785aca01c3f4afa11b8daa894db9bbbd00390f13aaf3dc126cf562e31347b2af7f4c4b8cc9b2d4dad91d7d4e65c2b6c6d649776a702159a352f85d2336fc8bf3d231b4eb876cecedc88e442be72348d06e4524f671d31eec1f1663b0749ed248baa9a2ef208284690d05681c667b1ffb11bff3e159570df9effae60f556653f56c30e20ae4965a7aea7b76196c1c66d7ff66254f47432e96aec010802706e4bd6fef4e4cbdc8a6ab687d943cfe1f60f9d3d4ea61764b7a4dbc59240ba2fedeb894582fbfa344fe94c57df2061530210bf4ec5fff133dfab1f1f51ac11203badb6223aa928fb3d46f1e7b79e1533bf0cb72878406cc55d898c6e0c6b483322264f8172cc5cab465bf2fe159013f8f0c03a7d6d78a141b6e4bfa35ee9358c0815957c5dab4c168a6b04d156b29a3a6a9d70ec614eab4ef8c5590319902d6b6899d3c26cd52a11193548a12840211129fabee5eceb586ae20911885110e9ce50c6beaa6982e3d2da3798f369c91aa09b9accfa75a084300492b55a37ffeb9becf000d161a9b6fbd78162a1a729028daa22c8771fb07bb0e629dbaffafff7d758430e03a5f0bcc4e0a9f7e385c40d0b188bc959db57e4f933a6860f956c2299aaf71c723e9d6662cee2216eb05b7af9b08149fca1a71d39e2b33338bf973f6664337e84741e0772bd03c21bcb034ea8d493db5497bad82266fd7414df08ccc82497ad82f06f7822614b398055ca2dc6344eeb388ee1a7d41f6d7d38ec4611f22234d4ff75f6e3f0d73fb5a0b8fc5bd2e3fc7736ef73377d429aa9710ed560b853752e9eff53d3b1a58dbdc78633c04fbb41cdcbe05cbb1d37c750eb834e6ccc747bf631d966c39f6f64f57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf78d080deca8f9e92cb0d15c89eb1099f29cc67fabdd117a42b848da5c708aad5599bc04c9837d9840fc676aa0125441a1fc8b2667b48326232244dd78d02729e90fcf7e020d962d6b3f74ff3e752e28da8578492bb42724b4eff38665ef756d8d1327fd9a9b66b6d793f80755b893a110bd528aa9e280f3ceeaac4d8a70a543755180b62a98895f0ce0fd41bddf7ca79c10580af52ace0f8b1fe678c9111b99e132b1e8b634f4834878fc59521649dc31e194a3b1c90a3e498caa3045f56978c226295994f4bdd76ba6f61f4dd13656ad86caded953f0bc878a23c21ba7f585ed97fdeb7864aa06c247ac2a82b3b9af9b2da727de89b51a013dbf96804cd6d842d847a8beb5c686931db41b3d9622d9328d815133c39060cc222a909085352514e38d28f7f002260a9d7be55f0247a76c017aefa681b72c1cf0d95329f47be6483676610da18b2dc31ee93a8684060df9208c3b49a3430c179c5a65d8c2cbc3089df0c4af285607cedbb68eb542f5e75f701d3c3a2725584fbea69ea2ef61be267bfa1f2286b445eace0c807176ff365dfe4a3a8da531817ad42a2dd719909589634ad52266a1688d06d0f2543bbe1450b139b92f68949ceab7d2f48109eb8451d1bcbe846f5e926f5c8cd7c4b6d42e0b1b0078199facd61a290b4245f04b37ab96423e8a54d5f61d88a4ee01bcff6e82d18143ed5bbdf574c69afa42095366472243d80d6429281d9ef4040581d95fa8adccafb4de4f3d8f66eabfd77f03f94b5ff668d50e73f5047df76d32006ab77806f26bdf21b7a3fcf658c6f49fb5b30da6eaae903f197c68fefceab1613582de39e49665359b21b046720b5033eb1a46e8fb0fb77eb6373552f54f16cf3339d8f31873540e6953ef82a32e0621e836708f33978cb17f61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hab6f1d00c0924e465a3629f7185c3ccf407b5cbe90fc570aaf394d9a48dd1223c1cee5a9502a1da1344c5cf47ff0ebccc2ff6a8d9f6c924fc9df42171979ce1b09525bdaff137c57b6f541d28f3ac5bc45dc3774dd46393ee1dff0cf924bbe10c536a4eceb7282033d23868e6836588786a40be5a69554d52c3d2b517f408bcead03bdc5021554becde8d710ef1bd3e86c00f3f8c77a3a1f90773a818bca5f24ef6d50b0e6dc299ae44d6f3b060bc1e13fa6476c41b2d5b4ea570f2c132376b3eafd42aec1384b426cfc39e4a8cdfc25261a2b0f5da0441e9203be912b2c4e9a2973a9cf668bceeb4b5e076c2b581a14b297a8e32abde8ecc56f2d3119b48a4f6fd42a372ab6132c2271a0d93a5fc7838714e1a4a884180dc46719eb918e1e01270f9775fb8ed293cc1f4273913f82d002703c6723829dde7aafe5d982e6fbe9877bf9a82228a1031bbb8d6f11fe04300df3b15f722aa811957418da2a3a3898adf470465894d8d5940c0b1aa860b3b622c79d0d2c41b43be1a3c3509ab2cf527e30a91abf8d6bfcdea50bde0c5aef19e11a0d46ec7553080a49e93721b4c6ceaee9e08c62ddadb69b92f4ceb85b0e23ef4a6894694549a2958e0fb5e1a373f081614caec4eface85fca0d4d87503f6a76ca6bd1b2c991cd843af9fe36a4912ed0aa8538971040c2ecff19f0a47482bcd94f88843759683c76bab163ddeef920f2244670f97bb12ebe053f4b1d58473dd621ec40280525b2f1c86fd39e43dda7c1e08d982f1f2e52e877e5edc382fece1edcb367b2b258e4b83f18ca6aed211ee98a32d62a4292e81d6b8ba4d92c4ad02b0db16cbcacd432c794a5e9f3fb18a8b575c316ddb9ad9ac012356b53389874b679a4cc4dfc2311560ec59d7f4656ce65aa44f8a8168d9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3176a0836802fa30747f2c0c4f79d4fa7af0f9a0941b7b2d75aa95d4079c4ac9820af5e0b45fdc4918bd131baedb79bf3cfc1713afe3e47ebccdd04e0d0d3dfe83051e89a037b9fe5769259e633c5b5ef2ced3d229d92f4c44d56490e9f69afa305e688333349e2a8f17176055b820eae9fa3e800cc6d8217ebd79170a352422c5e451492fa47d4d0e744ddff10b47540e9e6fc190508636b110efd683af73d94d9a4c8ad4cf7c1e465bceb94677c7bbf50e8968466d1fc899bc75e5aca16715248d0e94e6e7d0f6c441bcfbacbc6699cc15fba6b774949711453c97374ede4f578cdb09e3b4859b1e24837a0bc056cbca30cc208e02d70eb03ee2e67da724031bf6a568b51fffd4d7cf913da0e2739829580299f28909960568b5be360231e4f3984c8f9453004fe6f162c4c0874754453662d81c2c02bd970ac94388fc0f59fa12c8e8ebd78b55904d7643b58d75bfb8d2e69b6e962d0620602c843c9ef65474ef45abb222a92a9b42249f376a9d7fb4511594a1b59a5bc40c23ad7fafd27aa85d6f0a7517eb8812d927497b4b61ae9b57157d64c12347f4664a9dd29624a64e092aac44caa3ec230d7b566ae067f8b153448ab0b6bdf2ce2c367c5767eac68705df07ec8bb3cb995d43f531ad908df75ad5e35a7dc9bb07908610e94f39a207cedaaf97ae93f02fba6d3c7ad59a87a43e035868d49036fe15e81f7151cb12e6ef69c974303f3885f958420513580a06958bba00b76a0d0fc3775c88073d84a3a06be1507d34ed2be61733a80515f4fc5991d3809ec6141ffc3a251977c03f6ae5bd52512b3c5d8b884b5e0a90572a16912f49b8d5818630982f6ace2e06df0a187817c1dd5d7555448ca8b53737a879210886d9a57505fae17fba767cce346f1e030aa8f8dfa5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbfc8fd57f3444d6d17b5f34c595390d7cb0f99938bd9213a5dd7b62513f7da555025372b6596169d0ad1fec01189c64ec8ba61df3633eeffb62ed61800aeed3521337d00cea54d9f31b82a3955b48c06995573dff483bc0fb034275539e829e1bec213a3cd5dcfbfc49881669088cbddfafb21c35c9d8059681a1d75215834eb02850133b3c02e1255a4cb43f67e9571252755a01a9563b9c209f81cfe1dfb324f364d9edfe1fc613475adba9fa379e56fe045cd524d38975e5127c51bab9bb4c12d6be0998f10181fe5943507c2d2ae7e17ed9d89171c017269d55d052211e7b5eff223ce587136df3b6660d93d14913fe9d8b41aeddbd5913234c83f7c73ca8008c5944b67b21cccb3732b2f4c0209bf377c28d36d36fe83bc4b0a1e934b333612b14ef33c2ccaac380e7dfa71d16e6e6d661d4dcfd876420d0580a5215433106a4d11dc98c7fe216ad9b7d0c519e268c3cc937cc9fa0258c59577fc7885f42034abcf4914d478632b1c80f3979c828bf9ee701c98f6f6113b9fa19abb8c0fb1fdb3364eda334ba705e61e8be89666d8fdc0ec3a368a8b68e8bac3c0b0cdadca092b9a86b0425bd438d78bd17c600c29f874b15bd029162d4a02da9a519d54633b05f678ad3e96e4ede6689d4b0d8d28839eeba7226c8cde334bfd57dad96898b0da80b155b643d88820b462197908a2ec4a354324b715114bfc117d6ad2ae22a614223cfb4b893d06afd9a957341e2ba4db8e40f74977727fc9f8fa3fa4de99740b2a5d9efc39fa7bf4e2789f8ea68d4484895d4057bd5f12fdd149f2fd50d690f98502d4aa5971f9215b0f48c787481e73b0cdc97ade79657c30eed5af9134008b2ecec0ca53c13ab68e90366ab2895907774cdf802b523aac22e0a1610f1dd934dc07f39ae6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h304b5d5d7136b91ab7ce9e4d416ece0b4f1506911ec0be4b8fce267ed05a52a5bba41801ac69ef8dcb423ef9f5fe82b15098471614b021edd65761c8c45155a3f1813e6d4f37b1f74025d348630ec56a598c6efe470b9e2fba9f3dc8b2584282ddcef93e2fef59c03610438763d75a96d7aa21b8b9e9d00feff484ad99d998696448e4221603377dbac5c139fed3065cbeca5ef2630f2da910ff0875363aaccea4e8879a5defe7ecf07495cbe0c7b21a570427dd3a734a5e008ede166ccfeb6c70e80bb2c916f43dbcb72c0bc7080aecc30649169da71e0b239907222c7986d70a2426a510ea9544029a8cbb9200c1b1e6b26f0bd4597fe57b0121fc701a2cc0849b12af0289d0f9c355813e0824d13b03dd1e70bd7c414d1ccf84ebbe983a288ab9784a444c580cb1e1f52592f43199be993ce323f09b34ec14e9dc248b045893ac40f56e0b373e25016c7ca5a25634b1fbeb879343a6982805dcd7c8b6fb26c5b6928f28147d6e8b1d4e4302ff15bba9d21b679de6717f5f510331348ffa3977c3cdbcc91e3d9eefc7d5ba85507d31070a3916e51005778d0c5a081660978ea57de20e340df47dbc7a9108bfd2d9d576ed5dbfce1d441687ebfc2ab8407718f222693e0ccb859b2c42ef4e44a727789dd8bfb8ad5846b7049aefbf4898cc060689d642da8c381bce19d8fad0d31465e645cab26a4ea9ac79dee6a5f0360338c6bd0be25b53bce4ec72e7af9f04920c405145f6a886d88b351ead5a4440c2b3faf5afbeb8f195724ba9511bd77b89907c4345aa732bdcef52f6c0d0fd267856469115b7285a48d589b8556ead21d6406d7bfe275912adbf1774c33f20fb6c6d0d385ee0dff8b2c2c61c5e6daa8921c0d0e19e9284de2f4b1cc7610583700155da755d515b0e9ed7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9adb86694abed93fdd121222636e6710434ba57921c6719025e04c821fac98f55ca6f2e9f99059831c4c8032b7b68902d5727fc73b4e03150fe0885ed0a7a24a6ce13f802a9169b215a48c142f168298b057fb502becc9c8f57b84261e7d3622a209be281bed85cc9ba682025740eb901beefcdbd42a7968905dc20a04c5605f824c0cfa061e55470ab4b83c46d9ebf948fe7aa8bf330d92af6ccbcc0da035046e26738915ac5d8c1cd986eae63abad60fe543d646c0fe2f9a961e7c9eee240d634322dff175893567ad160b5d593c126fb0bbaabe4b40e3b1ec8b4d2fda60b508ed0157224ad74555dac9fb0680a45eb6174460ea4643acd40f9e45e925ba80d7542746695df81ba065a10aac17e1cf88cce9f384edcbad546994514ae9b7441f8f9b58dd0e7c46fa6bbecef6638203dc893d2c72cc919770ee619931ab9b91ef15041464f74afa1d350476a19e3c279b7600851df8fcc5270e818c1b2ff1cc94ec40748f52754bfebd44ed93f4b92ae4ce0841504c720ec1a1cf9579ec0fd923e5c2bf7d3b1a63a349ed9ca39a87f3c7d690b110e5104308b53bdf989d68cd5b8bc3a11e89a44f65d3c0c3a71b7e940c533544c0933deb440012e10c7a00262015da912827004be2778b0e41e23a37117566e0be939de7f1f0fe6f1a4d6055fe7f4eaec3ca9c74692d5fccce3a6b4860c3eda79d4a3c90e594841c17feb9796ac40f41301f51f463fa60407eb2a2acdbdf8ecd61af6e5aba203ca63d1e323b1c2ddf4de3ea5d0e0b5ce612150e7bfb099e0832db35c8d8d31af0e2c4e26f922905d1d3a7f41a5d0c2fe8630abe097cea019631d954b990f4139d59f01e9bf1b5270e9d9c01246c6be6c02362ae559c17dec1f3db8893399e2e9eed4004aae31d09c2d950209868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8582a0805afc0d9b621f2fa609b83dc27f4e2c2d2d2a29dcf4df9b9005ef48faaba9e61b13447142c209fe864a8d140761f130e9fd4de51d7b1c1e7e59f39918d5af83ce7c235a94445c58bb37ac3d9a5fec978a2a8b0ecfdbb24473b172829c676209c10a41915c9b21acdfa4e33de25ad4a9d975bfcdd46d1498a0b80fc3e81effb22215e9e390bb8e6c78cf98f52c0bd41aefaf100d8f8ef06228f1c6b501496e4e5c93fc8204fd76b5e022c50854a96d5b5c38845983ebdfad2f8d587c05f4b78a314f75c326f7408517e026349dd2d0d2c37b19bbcfb52bbfea4467e4cd120ddb3978c28d49cff85ff105d713a6bfb840ee083bf09dc1f84a1c1c9e8c00d7090d70dd1c904ecf25c7affae953baabd477d6e9c11ab70b53086586474ff3c078df822d0ac92acaa3b0cd8727c37d0bc983f9ba1e1e89ff15abcf0880c2bf193c9686393b0436e0f7df703af87dc74323b0b7bbd8fec699395061a640d0dff78318e97512487ed9b9623a8dbcc4253250d8ecc76155c007755532693a434b424545938ae7bb7ebcce8aec34e63f04912b5366a3954e66789b261bd27bd0763391a6acc0e0493f57aec94ac124a5e89c5cacb3e3f256e3e985357fe935011c81599df9d8e50ff32afa7d98aa8c1fe0e19e9a2456638bd876503f258dfc6b0520a0139e51126e222defb1f4d72e0e184e393674023b8943dbc59eb4073c0ceba0d334ffcee77d3d8679ea33e5d29e86c20ffff64915fd93db6363dfc471bcd6316d5791e42e61e712acb8c47893efbfa12497d871bd7b5ab497ae73e6c2d1fd78fead0e0e1351a2e7c26f3d71a2e053e88af4ab14e73eb1fcbcae85eaa091df0f36217f7551327bb6f610fcaff555d5f8acc03f86a6cc442415f02e0851a52d169c673a7b3cc13c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7bac865e31f35f2d012f5c6c50f2f51b2034a896d297dbc5190b586795e45700a1aa94801fcb569c5120e5adb3652a85f70dc748e82361cbee04217768580efd0dc6c849698a96f38400811a58bebf81014fef59fd49e71a058c5fd03ba8ed9bcaea7ce02315d8323f374a36da034589b665c74d740bcc4140fa110f2bf0a0e994b366e67159d170921371bd133e6713b3c549c0a0c797a373ee5f3a102c03d9aa6c68c508090ebd86cca5220a727b7ddb635b3a00f28585aa1742494f23db3bc6f1b8662227fb0689dd294f6707a867aa910aa36a436b5039633fd4ef983bbcb02cc8cbae6f764a6bcc364333609d3b16b233484e9aab6b485d83a30203bf78a0a08c5d6b59372f3526316ac49157197a143eeaf240c8af0685f52aef95baf52837df81ae46a46ea589020f83af7d183881ffd78cc674580613f066832170636875404a6dacb441df553a7377cd54ebbffae0e061ae984f0bb89a149c4b987b094a51467d435f1154f39f4a4b4a90f1938a14f550783bf13eb8e2eec456c2a652d3d30dcd1e1c062cebfbf705a1184cb897937714c14eb3e576ba9d4d9c1dfc932f031a50225bf8e57ff7caa267f2515d4eb2c9082c1426246134d200c9ae56b54ae2bdd1c6890fbe68d228437d710da868f9b08a715fc9a12e3a010a0247602f41f459dc539ce288a2ca342ec8dc66b5ada60584fdef794d1f35705dac8a2d1ac3359c95e0f985183f24e20babb7f677c3a2f97729ba9e21fc9e0becf323a958c12a87afe3e548fba5babd60aec1a64509310c335d9ade40490e542d6a0555088a6d12d517d739f1e64c6ddbd48e8230c02fde23f6504bd594d6aaab1e71035eb17cd3faf3894d02c298547f3505091def161f69fc1d3e3497d2098897eac55fa00479022b6ff6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he498c762b8b522dd6fcf2d03c19f28d8c07f9237cb8292a5cc57b897b59da5fd3da1a832d308487b32197a987dc195a2b4d3d8e0069628a3cc26437b42f973896e74e31b24a5cc97ca6a5146660f9d08f3ca09621215feed6bb65a3efce005635a64ee722cf2b51d8d6d14312b31b1918cae09e721b7392559594f9a0692f066ce8f6e30e5e0b737ed0bba4c3f0013eeff4c1507a86066ac1f32a8041d9c3e94cc88ce8a44f3953c997a9b4a52337764af8a1feb8a68656d3542870d52f0c6635fed79308ef09fd9d2248b75235bf8416b1d93bdb94e865b9dc4f90b315170f193ed69b3b65cb2717abd1ce05e7507feb690fdbc476e245539fb7248dc4c0b459c1ce6ca7dc35c11a8392aff5700658c4ca1ad45c4887ba93fe933477ddfb9421d83b0e423e71dc0e376371362f04cc894b025b96318e6277f44c5bc684c6b3ae50fa18baff3fb8873955a476fb0d8050476775a99f7e5dce251577232ec2aece94c01c67b8f62b6a1f49dfec44f0b0a719b12ef498b2847584c908bdc50ebf1e196a732c61c1188e7dc3c73cabf9d6045b02db0acb549fed97fc0a2018d790435240adeec4583296f6d7d0f59fb511ee094c4e49e9da33641ef1809a38fda7bcb4b80029ea3d9f691130517c405259b19f1cdc796227e1b7a43d1125e0bf5944c9ab68cbdc0310f1668a997898634e4457e08a24ea5207998d7278dbc1b924cef00809f27f17c9624cc725a39f0bc664d10546dcf81b33d02e7767c730a5057ffb2d6c03f6825ccea1f4078c9cd9b78f71aa8627186e7b927e81e32fd971709a4127e18ba22639597334006f6b06f18a71a7a7475aca73874aa2d91ddfb7b8022e321716c9ff7899ef38a6014a69c78f0d906eaabee475060f6b8ec5c4b7fd14bcc6990d83c92b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h27d6a3cc995368a3d44596e2f5c13abd4a6b90693ec70b04eb68ef1807d8b184cfa43040ab15a7bcdd613fe876efd3a15b342107d02210ae26af18716d9131831fca97adc6b99e4d76a32ac346df3d92848aa313ab3b0ff68de827068ba54b6b8de26a8bab45ed1b3037a121473a84b12ce00f329305a9e68fbbeea7b04fb0f3e318aeebd28fda830e6c73434f4401c30df058324070f90849a10371e4a09ad7096c77265c4f4f10af77dc71dec211cc836d0def82b9735a6f359746e224d4590d93bb7f8b6169514e04937157b7a139f66d1c0bd19fd06e1aa3aa9eb13f7ca6dddf535fdf1ff86c2ce06988b49b5fdb2bc0028b1f4e6b769b086d7c9ebe767cac0bf1ff670622a592bbee9e402207746ae2b3b4f164e3bb264da7d2078ee4e72b27f5044b7d330ac02094d5bb03378489fc289d798cb8b3b63680465f5a9fb95643c0bcf4860d8a28f25ada05766440c1847ead00b2c01566a607f94ca86bb3cba87d2067c6329dd3f8141c5dc3853716c573acc899b14aa7e739810f31b1b9a22e3f23f0b41bdaf589f95b05a8f1d2af1cd568a47f748f856de1bf32f6b7892fd567b5ebc81884fc5dfe5072037ac2069b5aa8be18a08ea411abb118218966c1bce851f95fc1de642acf032fd53517772b827279ce89ad1e42db142f2d31153280b6d11386919044e4a408d2e762f04a332e0baa7ef4816247b8ca2a7636da0a9a6561e2fd9d8cecc2f1f6d1aa7258629cad30ac1e8861d0d803ffc99f4951558d72fd4b5eada94cbe1c1b8b6a36740efbd843eb7e483972a846065ce579f18152e8526289d05d2538b8f1c7ddecdae3e4da2f58137781ca215141bd81785bbf4103d710bbfc8016a19a6f1f6874920859cea16cd5317a2cf6663e5f2ea1281929784c1958195;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfbf5e1f376287025dfbe1bab34b1277b3b3e8ef24ce38cbc00a048a5434d8a2160e5389ede8c652f5e67ead4994dea0309de64208d7bfe49ceedec7120a5e25aafdaa6859e1922e785df24aa8429545be92f6264db3b110bb5e8d4be70556fc015e5dcc778b3e9bd590551834f486aeb95d367fbd4198bd3b03eb72c5d99a874fbfbe63c4c1e111425e781843338968dc835faee9cffa08f6160978dd3ab9b8efddc3d2352a8ca00249e8a519b5679c75e65e22fdcf4b8f3c8ccae16c444b70f51fa54753954d3b2492e1cfcac7a9f1e11abf3f66094e44a1ba123d10de50d7737a7e542c7c43ede223f2c878ac53344de18aa8ec969bd52fbc9a6b2206f2fa6a0b9f388429202148fd938dc61478fb780ad21d67fc540c9666d0040c35e4a43f15643842bc35881745b97f5ae91780325cbd0c4b68bc53796f2daa7e2bf2afc33788a72e3877539b0806e07160c1c0049c6fdbdfbafc3b17cf8c40a12200139f382419422dd3eff32df995f8c64eb7eb340be1b62a47993079d0953bc8f877ed6e8439b6a38477e270b3ac5bcc1481f099d3d2b0980f77f74239fe5e84089b14f1591caaf0d6b1716b3ac29a9a461f7ef4fc0be36ad23a845106593630fbce63c69f1f25a63bdc10b04ba6f2213408a76d2e2022358be372a3a993444fc8d0f7a02468f9210192114e17f9e181b32dfcd261edc8c2326cea28c7dc067f1a6cc12ae77a16aa83d5259f249b2a5d44da047ecd67df33dfb1c0daa930ca6abf22856049229cd1b11c1ac06c977e16c8243a17ca2e596b7c4ff63c61c9ab5df63aa8a1217c81def15dcde1b8d617579d256615db1e83928925b7b4ac2d0e2064f397b56dae506ab4ac99423e03caef8a29a1caefe9b5b02cf43ca5619faeda057d1bb451c8da6fe2660;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he55541177add719417a8b7c3627bccee2c93136fe5a61e60ef723f9d7e31cf185100d62f253270108a79e423b8f97aaf841b514879147fa04b8428bf92ae8ac5cc8b342a2861f0ddeca3b7382ada34844c20c193cfc877e173c5b4acf104d344d2e40ef3f4867953015bfb83182bcde4dd970185bfe0f353393e9d4ca060869a9849410dc39002c326bd204d4caabae249474c1750b610e68293ceabf8d448589230d0b31841b87a946f567286a1beb1275a506c51620999136d4fba8ce00c6f0882e6601637d605d3ab67adf018dca20621fd723ad8b9d86575afd92b0edc533d532179be60d554b68a9ea4e8f3e98fea72c127bd5bb0a10ccfd2e8a4be47901449ed81aae731d21c5ddfd1b79ae0b2e0890032b391f35c39d55d9a040e39bc0dabae316ed45c9bbae47590e1bd0a13dddc87eb7bf1302e862b1dbd017b9c0d9abb084d9af06b5798a765ee9b44f8789ab0fd5d8dbc58df58f616c21db943038d8b45053f0186692b0c4f5bb2f1324cdff641839c29f19ef89e825aa2684dfba29b6b81db1f0050c258f416eed83acf4be7ba756c6906b4728b427292c0dbe3725d09a65bf5ac7c0df204052eca200c6d9e762edd241de047a8dc872a0c81209341d3e8e560b9f1400082d59ff450b27ad0ea7d2bfdcc7c1e4ca11e9c9fe192cd6670ff12fa7e155d06a9c6c6acfbf3c4f1dbf4477e9cd294e15dcaec10c18a7e1716f72b43b59b45ffefb3656b43b185d5ba5e99432f3c6244d16cb2ccd5f57862d0e7ccfc822b66af1cd285ececb657f62ae0d9d041985e01adcbaaa4f0b566b3fe12e92228d2359a4dda654781fb2c03516c21e8ace9fc310552ffa2d19961632208cbc9f8f27e90e791b6932b8d3984e8b4b64f6887ffeb9f7749cc1b7056186cb6205f96da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb41d3303d00dc84ea0257cfb8c96374d35ea7cb180bcf2a957c8759f7b92be9b71e77da2c56596078bc6c90c908caff5786eda81f70620dedbf99d59837289c687dcdfa9fbc589d8e468867ced0b645c1e073a2e46579ba3d36d9c6f86bd2ea9f9c43cff58404d2430313c5a306f9a78fc22b0e634f5c68204ff34f8a509a45463477741b620e52ca12c4e32f4f681bb7a762ccfb9d03bd6ca5539f4c16e2ce05a962439e3850121b70860846d122fd576c830c50f29fe44feeec4416a7748225c7d49645f803eacc30c7feacc5570bb0ba3a8a635bb8263cbe787f685d8f9586d25b0ffffc71fad727f7cfd84088e678e5dd0e183d12175f35d155bd00263cb0c0d9077f258bbdb59923ee3c924f018ca8abfd960979961359a47841b3b3b9a2d54e7e84279c68f6d6562b2615294df5bd5a0da719db1394f037ff7c4649f1d2afd88944f06948f6df21deaeab80bc6c9fed1ad33ff0503657028daa7869c00e26b8ae1374e49b33674e7a082d5409514ed1a164900a92dec8a4bbb25f8538141a4894f540b2da0f98be90b067348d29a606047a93d0de242c8bab700ef06f547eb28132e871a82d15378593158ddad610f402fbd275c2692e6b9c2f09dbe5d00701e041d3259bf414bd5713650b7a97e9ac5f9033993c5768f322fe0e94245c008d26384363d365fe97081011ed2139d7e28ef84987a140cc1aeb7a23f99d2588b96004ffba094f883898b96fd91953c90df94af0eb2ab42078a4418507cad612e04b5f077ebde8e9e3a46d26803327300b558a7b533da2fa6c486e2dcf692eea2a2e1c6e8aeecb4194873bfaee8bab5f9c7a55d3dc0fa92357aac530d66b5a761bc9251a02f4bf77e7698be5018b87f9f0eb6d4d3010bfd8e3cb1b9a05d7c685c65769262fb8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h92104ea2cbfee5d959032c729e1f6425a429de2bb939fe0c7f74c02537975755bd550e55846cc964e51a6cb88dae247908edca389691a20588464651111302055983565c01ec00749dedc21e93b2f4ab3d95c0af42608dc576811170a5b3f428b5870d9ff3245b2564ea280ce4cbe2a16edd27225659c37646cd6d0043791474a3c938aaf3cb8a1d948c477fa4f27931188a5d67db7eb778f4eeb45da4a37b43d0f3f73611cd3630dfd009f059e75659c817d03b424104ebafb6ac49c78941b172fb9b149b8bc32731f08edfb28e9af0673de3ea108c8363acecba36694c6a9d1bc76333a3214b2742dd2e7fa4ce34a7c24ddfce87e3b5e2187b050b5af64167f6d57828c71d7b264bf9e27ecc6191fd89c06925986299859736127bcd9020265c9871269871fb896edc7943e2eea456a2e170e6c2463d42624e798f726c1208ad83cb374922a6ad8d004c576dfcd3372ced4408fc8eb913ef44d0a79199d234500cc0b71aceb9dd992a180b0c69d4f20d92f4778e222d4a1fcd0f0c2897f831afcdad74864ae27f2b3ad5a72c4dcd3a9192152aa830155693fba5eec60d9df9f3850e74ce7d07e013d780c928efa5e40571cea2136385730ee15a820cf01a3cb2f5a8eab0065409b3ccfa8d1c97d9e1c6f1c80d14a10cbd52fa15cde9f8b52574991faabb120a9c4fbb60f5a83581d907b8bbb4154d26556c5ddf8cfde19d9c45dc009f9fad09c366335e9c06d7b613509f185a38405de710caf897723b6e170e655674e4ce63ed90628f627863032f612c0f90c5a96e11c80272342a1952267064915900d73cdd8344e41782238ee7e9d851226cce59ddc2e9f1cf2627e25d6a1a1ba7a94c199fc1a7ce6dfdb413e3b7199e0207f818997cff0aefa2d850ee3c91fcc667e23237;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcd793e191c198fe41eb49fd35e8e3c828779f4b82e4c8a494ba58fd0428fbdc34c35c83052aa8e6f3d7cd4f99fb2706d545084c743d8c2d0ea0cefdef5a690a6cbaf5c0dba3691ea483cf5228064f0232fb74319543018077295378842a67f49e84ff56ff2cb2230c3f0b6b10efa4c7190c23c23531913c0da9c811ec8447ec6c5d2d613a321e256adcb4f066c70c1e9458ef66505bbeda3c10c06e493fbdb10f28778e3392715b1f05ff240407c705e21b72a4af0abe00040546f6f1fd51cc5dee21f036a90b371bddc48798d3f2a94408f89dc21eb9be6b3c3096dc04078a1040eb3368ad82014e41a8e48cd3f0774ba063c906fd27fb92685f88052670b7aa7c9c2763475b1a2bb486a3638df71cf5eba1978b49a25d6fe11d07879a498a51d1fccfcdcf1e73e415869aa2da24c69e435e92f6712e493928194fbc51bf9de4e483528b9f70a1db6d40c7f25b9f42d46675a41dbfb61c3c06cc4d6cdccab71a4fbcbe6ca7e6f3c67a452cc61e1dec332337ff27ad46d8bf88b544beabd54d89394a5305e51c7a87f1749218d2d60ed2bdab8a095ab705229b2d4602cd63d298f3b8f62c1b5331e94330743c1233930dd30b6a6a7ceebcd7b5cef5ad07d6add73daf127c493ef1ee16e0c3f189dca3acbe704ee4f4dc99b95dc18b50505079f60b657cc37b350d4dd6fe72cb8390337f142ec02aa88236468f909c226514148621e6176bcec9c96e10295666d794daa2d5acf40e0615aa683b369dcc4ca5d095d1cd07bf0c4cdedaf092f7daae3a6b8219f89127bd66d8cf51c2d8a30a6f44d2d94d71d3c6dab337a995ba0dccf19c27259e935d1101c444b901c873e785f34197f640f372844706b424dfca6538bfe6c3b1fa306378ecc96b619a10af252b381773acf75e447d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h383bb240c0338ddffd30df01d9d80c0baf0873fe7b345ceb62b2a866384c07124513e8de2688011e320a218135c65515e8800ca48e803f41e771b83784df972b3234c1f08a35c8413862dfae8ca879ee45429d470a0ae9d682f35c9cdbdce199e26853ff8c8e50a41b4475973c94819c2d6c1af680419d9c682645971c0f2042569ea63df987a20b6119cd8f483d0e941ddc28ad1ebc536cbd15a6c75d445f0c5d1c49083da46165de0bfbbd68ce8a1a86ea815ddbd9f3c22476b076c906c07ee0cc3a6752be89d9281b6755b60095361bc0d161eb2b2a81facf4ecaa9d3c6d6b1d45f61e5bc79edf0f285ba1778e51ddc3cec19583cb0b22f8be79a6b9ac28125883af776ffcbf4b438e05a2f271e06872d9242c2f4d6a07379ef026328b6ffea6e68fbf56e33ce8c08fa232b3d4d0a6b41acc568205316228f86a5355e45e179ac2fa2c6b84bb66fd9d0e8999032b967037692b2fdd702596f0948f79e534396b89910b5e309621fef8f7aa76a7b70d36e927ce13f6c8874873ce1a18b1ff72dcdd9116c5bb332963fd023dbd9617b55c7c18265295150f63abf91e584c21017a8e2190dd5cf4c1166e7477c59864b1e6871992a6020c19ff2ac70afa2e5852102e4085a46701a45f310abb7887430fa7038a7c4c4589aa4dfeb0b74002f3a879bf365a9fd5f1b41f4287ed2cb58d06f81618f27f93fa7141394fca169569a7f764ac172521b37e2c0730eaaeccd29bf8e37923c0fe99b959dbd976dc094accc84aa69fd4019235edb15dead58afcbba418627e6e043e4a1f8a9d4522df61a24536cc4ac3de1acca421f05fce3d4ca2beee350a3ac9d45764c75debc3240f29e169e6b8ba204aec0c76da8af7a945f17f50b928b880d67dfd09ac1ad19b5d31f13731cf3d961ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hdf63c0839fde30aa7d1b745b4e34e21e05c3c86f5c96283f8613f8540136110a241d81b9b26a48e6ab3598f959dda810592313a4f03108679f35daba66a70ec04bed6de33d3d39dba35a42bb49598d6d883ec5db0ae74b2b8b2107137666115322c5b1760959ba2027ac9fd26d564090fbc0792a65bea338370ec8e725978eb890d5c9bb2068189b5752547d6a6ae54d87e14b676b2da1dd4936ebacd841d3bae9bc50222479e5ad3f8a1da962481d08f2a6505c6febdb6e58b62882869406f61a79a8f8ecd17b5d63922fb8d68fb2fa6c6c1fe4e42b515b7798df796b0a67a0581b6e65b18e0fca69407d7424c7302fc1a58052ba28fa4736d61a496badcdf104db5b882f93db50cff44d3610aa9872695c9e620cfe4a03a121d106f90a3ce89b45b500084aa22adce8ee04cef0d5dbee6e9442ccb10ee5efa11d68f8c80c8dce5c5b4ab10ed9b3ca53a9f2c5b53776445a1845446d25c92601df41cf284320a9b4032a4b600c4060c668b089989e5159f5854e609e44e99b7b5fb8c3c38eef20e6190853669e1d3b17120c899b61d5259d2196e5788eb3debaac4699b1428f8f97a62e28a6d265b68ef08e9020b29575d1169be0199e40ec7a349c643690669fcc6b4d91a7b67553048dec73ff69b832fdbf3a65ce5cc3ce688421aca4de9c3c2e3eb2c882a7efc9e012863a00fd312c1681ea9f8f15cba312d61c2f74e7a1252289c89518a4b8a618315bb18b0cd7935c242fcebe3745d15f36c1d2cdb3d2c610ec93d9166faf3b491bee25d63b831bcff4334ad7fbb2db8f9b795e3cee4667c8e05982c5fd70344da5c39f4a997b30824cecebe5496a81c5b32c8323799c42815427060cb56ca0a4d32f291905762bb67cf986ee80acbd4e0eab2c5b66c07f7a976236309c08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'heb8feb9188e7349de1fefbfb6f121fd311da7331e903030eb50c855365e084273629ec343db66e4440ee83d014f5bfe013931a3651a074ebedea4874cf184cd3a656c90f32006e40535008363e0fb97148c98d61574175ed07f3393efb4013424912dac8c8fb400cd1d30b1697085d059603ea733068caf32e836b0a3f2a9f36169e40d264d269de30eb16aa85e47a9ac879d8f5c384199699ee6b37552a2f344d1472403af405f3a8fa31cb771dc768b33e307919f630218218e389d849040fc45ad2146747158f8ba8be30d24e40066b2da78affb39c74b84a4577e63c13283b0fa9e28e2375680abdd187f1c8d7ecd0b39b24472a99f12430f625d16dfb6363e63a8c4e40c2bb658330aa588c0b1652d28f362b4c9b4de620578e8a3e95bbfbc07b1d38b362d6031cb761ac6c92df7b98eee8a8f7aac9d1925a4042b8116de69202020814e2edc479426a8dc19059200ae1977f3156ccdaf78ff03520e5305958501c8fed168b7fe662176b9cad128d361f158b94b9e7601394c6403365bd49a247fd322cac9bb0bd9fc883cc88e6f293f8c5c7012222670e700d36d0677f2d287c3b656c3a2e4eafbc364048c19b8ae714b6667cb520e6f87b58130a29870c58972e91e99a78770032f3c4ca21aa08baf8de41749b7ae0bfdb29bae17d21b5f198676f8aa3e2bc913bdb8381514d611e7da76ae3fc43c0de2dd5fb6e7f8dc6a43ef53334750409eab8cbd2458b57898f60a566f66a0360e4f1f74847bd190a58f27b04aaf8ab854b2706818bb02ccbbebcbd4f8f66e68065f76f94901d7599642ae78ad2e78f1824b868630ac8060ee407730de0cb61560c89846b5fca329c30f3ed7be533060efd9b34840fc13604690a733c1b35a7af73704787991aaa913bf4c58af9cd31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he565df0df7ddbd05b0e21c912dbe004b8a0ce532601b4eda6ea21348d4bc3d92ad684f769dc6e7962d44fcd0b994bc4f51d8e67281721be2ce148c16c7787cdaf6cee0f7d28b44d1a356682d3d32e392b19e25c99c2eba62778eb5f3b0e95707ed35020f8428c3f8d8410459280cff3083f06436c3ad5d2a522e1c01643285f1b9705ea9e31f2855cb02bd26ac2d5b89c256fc0768db100d4fa6b82adcc663813816bf544f27a7e2c18ab8e410ecf308275eebd8e490d4f1faf574473c3ad65a83ee3fb2f3f31c0a1ac1a60901e16eb7ec97ece1cc3951c5f136f5bb92f8a9ad5223c3685661e7bed7f8a4f7bc6f3d8efb706205012e5ddb9d7209f5f4b70cd1a68330223bd2daef6c2efd81c03ee956c3ef1aeaed881f918f312cf9d53b65757eea789dffead717c1d09c1be58b6f9c027b49639f126c9b8e82442c296d9db7bafa7f6bd55e64f857e621b5e7a9e56d31d1695f9505577a7d1cf78ea37836a76745fe005db60698ab0727f39faca40cc22a26571edc6f3380bbd74592caa1569471e973045389ac0b6880c7d646eb1e9bbee79b23f131372d354cfef773d4bf9aaff3729731d779d1a20509b5e24fa5c5094a92bda29bb0e4603acf3a619c1ff77aab2aa1da2b3dccffb966eddba1c2b1a821a90801465f33ac1c4e73ea024402409d6fe13788d3e21796cd7d0c3578a8f33def074f46b3e30649e5c0465e44a0c08da73f2b9a5ab22c77a604e9abe8418808626c7082448db4208796507c56b783853f77868d2e2ed5c3a5cfa7b59b2d7fe8b70efc232dc8f97dbe448a7fdaf76a25553753e00d42b093f55581939acbaafc55bbe8a6471417961187f46b8b3542fb1792c5316e722541233775e32bc98128d698313a55adc69fffa63d8c8638b8b6d057327a93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha0f707576a6aa8603dfd2ebd64602a208fc7d3fe790fc2eb87c8bc2031b53c0c41494244a1f024166e3654bbb841819796a6fe4cba48a3882633cb2eb27f2c0137bff4cd63847327ca892cb0c8cc621c110cea866c418e31689694c90cc3863cb84d88abcf771fc78708097d1256f57fcd10e354151f7889698cd166890635fe600a845860327b6b98b0b2513e3d63f166889871b9880a96f2c9272955511d8629a0c5171ebc41a514cd47e9512c306d9501616a12ce25e7e8d4ae5c07d101513a9963cb17ff9afa41ec4c2f13fd5eee65631ed129a29aa1cd3d75a8a6e1f3a1bcecf4ef30a1e4890d28d399e4ce3329702e07269aaf8a70464cea31fd034269e1c70b3a8164475af455dbaabd75c494bc5371b80099bea48d646d98292eef986f46d06ca7e46ca23207f369b4b672d469ec33047c2ad357270df06377c541c991ecc49d586d16059cd7af35d92ad9979ddb3d12934a81c8c6f6c53ababcccd92042f5785e1945d86da6c5f466c2bfcc46afb32bdc55dbe1e9b320d643fd355ae04f374bc5acf5179c9c7e80c6dbb608a6f00a0e6857a4ab6cd0f5f925a3d847038578be52e1cbf47b90c540899562e7de5ece2c708dc1695a6dd654930888fe99ea9d1459cd5a054fb12e631e0f93ea5290e1f76c6f8ced8017437b285f50b3d51d0239a522abf68c5d729a7b1757fec631a6a150dd9c18c80f5e0516b69f3776b9e9c132fc7b8509954608d5e6124bf2a27faa862ddf491ec336f1e2ce41c995d53302b12901fc92404cb69a1ac84f121689ad9a996e7977f7fa382190749e36a05836edf1e9c9eefb744f371e9a8ced677ea16f5d2a885a065c066e2c03089d0f03160ec42613cb2f07a32ee5a98b7ff7cbdfb46debe7ac0993d2347adcfd9de8d61cf9b54079;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1a1dce4ee37523e67395e1a171b3d041e75d59e9df355254a5bfefffd3a313d78771032022978725071be3a3dc662deb966c23baa6b97ec1aba407e37a8fb3e97dbefbfe6f9992a78a4b7065671441074a5a028092e8229e5126b344f3df6325db8a1ee141982b895922e5c4c0cf281a4956267ae73b1835e871efeae5ba689727369fd5aa43bcda11423c0e30a27f40f13530dc2bcc6f49b2dcc970164a8070c835a925f01f849741e05238b5d5514c2ea475b9e2646eb5fc55572b7437acc74e054e658f1aec39b9356910838c2e624f98721435c60356a4f288642aeb67db13c71e793c53c5f65bfa31d36299eed8e094b19ce85502399efb74942dc911f2a31f0cae16ff9fd07106af8e92b035dc4c537fb05850cc74c104e11881a5a6e33ff4754bd07af67371b1d84c99511ce7e3b3628388a1940e28382789d7dc8fd684f586d59a1ac900c235c9d952ab9bd47ded2faf966446a4916f8dc760da145c33ee279ea7ef09771410d37e1bdeae18ffaa86534ef3237464bbc34dfc1fe50ddd89339d1fdc4940fb699b2e4670d42c2face8852a4971038b067ccf43cb5a433cb0903238426a7c80f340329136f1d49f5f994b3361eb0d1e801c79554310dab6589a46d1932c935c2e5701b4bc6560d0b9b9dd34a061dbddba32fb1edef6225ed69aa7162e9549e3197dc17567edddaa833d4839cc2c726e76d762dd9983382def1832dbe6c0463e9cd43d97ec56b886fe1be03f73250d3bb8968a5456217f4a5bc705f76befa9e48b8ad50f624dc5ff5a641627ed3d5bfa116bc7945f45189f23338fb5f53a7ca6036b83346e616490624c8bae8b64c9812452de6b550f31187aaf0a4f375f4ab641d97030f6a67b6c9a24a48d9a31f7b7585c4d5a334977631a80bd9d1505ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hdee6fb30464eebc120b10d18f55bd77d0e2052bf69507259d13a3eca7a09fceecb013f9d06dcc1277513436283232b286f70ba0bc141685a2627faf2d22f63c5d39a62c487f117b2f7b0b69b7ab1eb83bef2dddce6e5525491fbba3a24e9db2e32fccfb2bd95ea91020a2282c18cf7cff4a55a476c77cf49345d448970c0017c10543e7361fb0a74069a9d65f42f3f4980324d8580c3c78c81080c7e1e72c1122f18d98611a2afe8fbfb6fa5f324e140880d1ba8641db760ba3e7cc009ffc521973212ff97ba73b9663f9e6da6db505868c641f1099af5135557bd27e444b5f3d7eeaf599040c98ace8c1d47c475dbc9011bac3448f94f4e8707e743995873944455ca37fe7ab951a5e5a4b634196761898222b4106a0ec337eaab55fb80af71512147da5bc06f393062ccd1f0b9a86b7ceafb9991db00676ad4f56c3bae4e2e79c5a3a2eec89ed08dd792d203f031fdd095b9b356466fa496085816bb98e06076e8298ea2ace9f7003efe32e43de43ca593fc757c5ebcf67869b11e4120d9d3495cc8acde3a5fd13b5c8ef009d9dfe5f2fe7c8d6d0ef51dadb12695b72d4b295c35120476a433abcb8dd81c939fd3505d43d6d354e225b1ba6b520d1578f585522b4c87997a1d25bf767d6fb7d371dd4bedde1928a96613522e0b6da561fe4efe1cc15bc6954c6c61348b8b3bfb9fe1a1345b45b5a7d62af6e5edd6495b2d8c3b385ab3043e7d834b4edb34dc3a88175425ab39e63c73c6875c461bed2ea8bbccf6f083ad0ff2950e5d4d78692cc4608e75c8b07d45b1f600fe834746a5d3b85bf1201628a8752d6034e4c9818e76b4fecdb74007e9bdeee331bebab85254e7d98a8d1e63d229bb2a405f5ba8c7f1e1ce983f62ca2b4a40fc9dd576f42c523b2801eed25b2a23f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8fae489a116b1493ffcca9506e4e6e1a28318ba8926af68fd235cf980690e8eaf0561b09d00ba7272ce2e8be21baa8e76aa0594b2dcb6424963c86446c1e000a067b65a12daca12c00b18825f08b96b65c0403ca15a62c100028bf82e39a4d2aefe680ba900091df939fa235e1e67304a4cb32ed900c7c80ff818f3f7c1f74181dd66a6b4aae1680fc509181dcf59103d19f7ea3b417486cdc49e86ac2ec2151bac33562fdea02dcd296fa98de24fae478bb36ef0d87c2c647a551798f265e5e5efa2c618b2058cbe65d1d099928bd95817c3f25496389653e39c26d154ced30f019e252a2ea25375fa271c4b6a459d1e097ea3fcaa188852e33bfeca6f582806b844c8d81dee74b92b67b0e32d8dc2dd1ec141c4e72ead5f563cc366ca434e2dd9427f93420273ca17d4cc9d1ac77ba0435ecfa35b2f149d5f5ab9f757d57c7395292d380bee022215a1bbc34580f3437968349566ae2b950ba7df24b4c5dee6f5abac82cb588edf63220de3b291de1b02c372192cd19daa25ce9836522ae70e68214e45bfb92198b4596ca629ab54a660dfd6d626f3ff199d4a0f834a9bb06188c87a0e0b9a579727ed11840729cfa47b14c86a0e23262b06d574b1fc22f883c388e2b50a24071c2995f7f51dacfc87b0e4b8a621b7540e02bc85409af1a990d5766a31bc63bb7da6f3e7d8942750b0491a23e37dd46bc6846d562fd72341848db703a6f27f907d2bce4dd1638a46e256311d884f9b80bbad3e278a29479605d6fae4bdda40b221f4cad8020af17c424a22494dbf7f1e7f5609285784e5ada0e4d47a5c24f4717e85c6bfc2a7c14cf231d6814e0ebca51b453a2e33fe083df9fa16dcffc3594db01e32af8ed1bbe509d88f90c6437bc4870a72a22af5a178c9f651a1f649da9d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfd1311177a3b426af67ab7210119dadca993ef850bf6dc9230614e4eaf37f842af1fcba2d140ce4a03166daa8dad2c368b8d5b7272b170653a18be563000fbb8f650a9685bf3b34d477d41ce4d9bbe0d36f86aa5dfaa1c269bc07ef68f1888d7fbe49fc12938e26e836fbc4e328733d6292a2b0f9041a154e583ec97f3365fcf662c624c4302d758a151615b6283b8a45a46db8cc4205641e7750a22e1891731bc113286bbd67f405d76e4b1037ba656cf269b576d7bc09d69fd993db4dcb863c5dbd944eaa2dc8e317aa5aee8e40e8deb4d663226fc0815eeea80137019510cb3ebf6ba75c11bfc5858ecd495bfeca7b7d189c2a6b017a28202d6dc3218df1a6bde68daad9c86986dcd7d2718ae8013823ed6273ad024f88eb63ee264b85be9265e4db56432ab7f4bcab9492f4c15d00d948229875656e7f9f4eb0735fb6417eef4b0715a91e843afc2b1d39deff57ff07bae708fe4fd5806cb9d4ce95c484a200ed27e9fea0a49c2b50a90ba047fd73a1594e353bbebb1709e51d349b4f4bf3098206b6c9ffca96c082680e0e5f2f9708c9754786c967d43f46d6370bb9d4f5bb46ff7bda9a1f025e2c6e014e1eddec4324408f028a1cef840b98022aadf3de98abb93b9fd0b9cc365d227774fb4cef4d71fbaf9ee42bcf64b50d1750b59221fc54a2c589317da635ae85dc564464b4ba45e55eb0be4a621031a134159e2c1c8f34ab3e96ce4b1f73d45b224245cce3a342f5597d5f1d9e76d4b4ec4c26f68cb22e6b0b1ae176e1bef018e576f87209240b4504dc53e06388574bdde277fc04b7d9bd3ad6ce4ef38ff39868b5c399ae0ebf0dc2602548ffa32d1c546750054dc5ef696ac647836919077ea7ddeecfec22b1018736ff81cf87702f186f4bbd0b5f6373c2983097e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha152d766db4ada58aacf142fa5aceccae59f2e90241b6d9baa649098f13ebd91e7bf0aaa2a3bd5bedf552219dace6cb325177ed7d15617c12cbfac813b56768a7eb240d2141af8f2d75eefc7382ee9a6fa960486c1801828a4902364d3752be2985f95e07d3715f99bf7a40be84142b1867be6c419baa0e04eead2132a799ed55ba43f955241a8b8e88abbd38e1a15560b5e195d69db83947777bb681e44af92b9c4756884452a948b1f8042c337de43d6cdfd45cd82c89e065cd03132910216e662e7bf85e794c7df0af980a787d860b6d53adfc8768393349f189537be82f696887b9bb99b6aca88f9c547f6bfab8e3a1346558e5daef8073fcdb74f0d46b5b4662b9140b877c59de1698e0a38908c1fbeb658a1c79d9d6c80b0a70fc26fa5ff8c55152954f0fa5f576ae7ac232d02d01ce6201b4a31acf3d196b21f2a8388ff52b17efa2129bc791714495ccfdad8fc5716db5b170a6a47b6455427b1e6fe9bfd1567717ae4c7a982195738594e3e971ac5fadb31fd38dbe0e19704d16dba168f31dde69b33fa44a0a112f3697223355b3d5eac498fabe3684b37121671a5daea26ca10cd3470d4d7521dc33533740294bc685d2f58a01d44f5212ff478de3d7c03b2eb2cd133103128a469c393743fa55793796deabd01c5aed607959c7e374d0cb1a8be613b82fcf6cf217012a8f4cc59f5c0dde1d0802ef3e36336cc206c4f479deb7d6f4f0eaf415a845369ee89bfb50bf4fdcaa91af851adf761003b448e1355eb9b0e41cea94dc40ef3d548008894d7e220471f4257cae146e3cbad20a2a972b7bf08d83c339d2de399f9756454f43db74cab2d1ad5f6ecdd4f1056047c14d9265db9615f3fea38a8a9e455d1ea0da3cf7e41a21c3714caea9877049147d52407cda588;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h627a77552a4f565467c4213b7a74f05d69d455387c2baa12afb0f80be3e86a9d6ae1e8001fc5693a0dc2fbc4360dd41a5a50c666d960a88960f0bac07ae0d5bd32e185f6c9a428b05e37e848eab4b711ed618f9863f7e89fc4c00409b348f52ad8e2779f95ac7ccd9374ffc30f5d87f098dcae170a5babde83ab0ad12a37ea967471673428175eac7e2ed50ac31083b1f6e2497e344ffa32a4a32c0dfc142644cb7bb150a7b7314cf03a7f5c767972a6a59f6ec7978cfc180bf5746d02917ed546e395848ff283686c48cfef6a8e7769e1112e606e505dc34d85321c049173aa0db746bd848e71998f266064ceae31c8d7c6c25975d027971bd5ba018e78ae9af6d64464f1f885ba76b49e079b22ea03c9cbd9c38e122d05d8dcb88592ce067733c70fefb05e18d639097b248c3381e4034f27d8bf09fa85f252401076d86f24176f71e7001bd6d9ac50a269c2b8100e67afbed4419b4b607b592206fc97bd4322df4a682cdd33fcf0736534cbc70ead45ac8a3c2b59349cfaaa3005380e0357fbac084cd433461241a311d558391fb1e57a7358f7edbbaa2e49188491c8e916dc87caa48d02f2eb699af289adc23e2746b5f341ff8c1f57689a0e87e4091b6d9dde6f9d43f07beca1681e4334f44d0a4b1287db4de094f74996c9ffc7e4023b9881aaf34462a564c0fd85caf33d8348995661f44e69929f9f53a18249efb789298bc27b41a9dce4d03867ab4fe1859835c578c3e80eec7a79130d60c09f63a2d8faad2936a5c0161645aa51e451bb15debc22e7431a6d827d574c33267866ece7b108bf84ba4330330504fcbbd5a76a5576584f13ce0793bbda087f69fff2c224b79a55e8d6044233f6f446cd292688c652eae18c1ee7474ce531f2aab4c33d156e13582cabd86d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h49b98fca255c8682884b09a01ed23ba7c1d5e892186a4d7142653b2ace7ab03968131a7a774e9283386668f9d004cc0fc62e21748f9476b2984664b775047eee25640475b6f926a724726d19cfd2c809eaaa067954986fd8129ff187ef2cfca2bf65451e099489414e103b8cd75f46b709e8bff2160e98208c1cbadac1fc75b4bd6ed031ae6ae234f324beca70c3746d5438f70f8b5cb8bd4e97793ee788bbf1f34633badc6dcb71ea67a11b984d8a650b2622b00fb9542453704bac40bbbe099fe9c16531c0302d7c064dfe7a477325e1a89cbd76a153f2fea74d6a80dcd8ffa315466dccf933e90e6bf0842b210274991510e5e79b0189e7c96d21039bb51ad46b2c01b1ba3667f9bffb67e0a9bf3ce45fafcc057439652ddaa881daad65d812df6ce48ae99eca9d2235a95150d23d0160dff3ae09ae5f56ff3c4a67cc8b3098f62034eb26eee7c0035068e22aa48121bf76314781efa08403a5cfae065b94c5ea36e695cc11d6507a276bdd954c8902cc02417370c8ca97fbd94323d892055b954ffa59a3433247f2427189d2a221276fd5f2c6aff0efabd65fe4eabc3445dd78a94b048faa84a3de0b79cfaee3da6adbdc3b7fabeb89c8425bead993f16e248f17fcf5f49f2d68b60562cb9f4b2feeb1da169afeacd19c3d9abb94d3af49a1df7d144b6e19618c4fb6430eb7eba0603e801b85a884faca500d3b4d0daa588b5584729cd3dee68e24ea713da6a8133c33de9d86910d110490d439d1b6f9620e7f82c7ebffe7c81f43903163f8642ff7c5187f415eae6a8436d0fba73a2dc7b505b2388e41b7f8da9517b4801aed09a3f227726bdf271b0ca4da9e243fb3a9b907358f946a3bf6a31f84a5b04a1a8bbdfd4211b2737662a7d43d68108acd8db336da81568e687e;
        #1
        $finish();
    end
endmodule
