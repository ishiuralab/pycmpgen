module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    compressor_CLA54_32 compressor_CLA54_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA54_32(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [0:0] comp_out37;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [0:0] dst37);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [15:0] stage1_0;
   wire [16:0] stage1_1;
   wire [21:0] stage1_2;
   wire [21:0] stage1_3;
   wire [32:0] stage1_4;
   wire [26:0] stage1_5;
   wire [32:0] stage1_6;
   wire [20:0] stage1_7;
   wire [25:0] stage1_8;
   wire [35:0] stage1_9;
   wire [17:0] stage1_10;
   wire [28:0] stage1_11;
   wire [23:0] stage1_12;
   wire [31:0] stage1_13;
   wire [30:0] stage1_14;
   wire [27:0] stage1_15;
   wire [24:0] stage1_16;
   wire [19:0] stage1_17;
   wire [29:0] stage1_18;
   wire [31:0] stage1_19;
   wire [22:0] stage1_20;
   wire [29:0] stage1_21;
   wire [21:0] stage1_22;
   wire [28:0] stage1_23;
   wire [23:0] stage1_24;
   wire [22:0] stage1_25;
   wire [17:0] stage1_26;
   wire [24:0] stage1_27;
   wire [25:0] stage1_28;
   wire [24:0] stage1_29;
   wire [17:0] stage1_30;
   wire [23:0] stage1_31;
   wire [16:0] stage1_32;
   wire [7:0] stage1_33;
   wire [9:0] stage2_0;
   wire [11:0] stage2_1;
   wire [16:0] stage2_2;
   wire [10:0] stage2_3;
   wire [9:0] stage2_4;
   wire [11:0] stage2_5;
   wire [11:0] stage2_6;
   wire [15:0] stage2_7;
   wire [16:0] stage2_8;
   wire [9:0] stage2_9;
   wire [8:0] stage2_10;
   wire [9:0] stage2_11;
   wire [15:0] stage2_12;
   wire [18:0] stage2_13;
   wire [9:0] stage2_14;
   wire [11:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [13:0] stage2_18;
   wire [9:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [16:0] stage2_22;
   wire [16:0] stage2_23;
   wire [17:0] stage2_24;
   wire [11:0] stage2_25;
   wire [8:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [10:0] stage2_30;
   wire [9:0] stage2_31;
   wire [6:0] stage2_32;
   wire [6:0] stage2_33;
   wire [3:0] stage2_34;
   wire [1:0] stage2_35;
   wire [1:0] stage3_0;
   wire [11:0] stage3_1;
   wire [2:0] stage3_2;
   wire [12:0] stage3_3;
   wire [4:0] stage3_4;
   wire [2:0] stage3_5;
   wire [4:0] stage3_6;
   wire [8:0] stage3_7;
   wire [8:0] stage3_8;
   wire [7:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [5:0] stage3_12;
   wire [6:0] stage3_13;
   wire [5:0] stage3_14;
   wire [5:0] stage3_15;
   wire [8:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [6:0] stage3_19;
   wire [7:0] stage3_20;
   wire [6:0] stage3_21;
   wire [7:0] stage3_22;
   wire [6:0] stage3_23;
   wire [4:0] stage3_24;
   wire [5:0] stage3_25;
   wire [9:0] stage3_26;
   wire [2:0] stage3_27;
   wire [3:0] stage3_28;
   wire [18:0] stage3_29;
   wire [2:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [4:0] stage3_34;
   wire [3:0] stage3_35;
   wire [1:0] stage4_0;
   wire [3:0] stage4_1;
   wire [2:0] stage4_2;
   wire [2:0] stage4_3;
   wire [2:0] stage4_4;
   wire [2:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [4:0] stage4_8;
   wire [3:0] stage4_9;
   wire [4:0] stage4_10;
   wire [2:0] stage4_11;
   wire [1:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [3:0] stage4_15;
   wire [5:0] stage4_16;
   wire [1:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [2:0] stage4_21;
   wire [5:0] stage4_22;
   wire [2:0] stage4_23;
   wire [1:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [0:0] stage4_27;
   wire [1:0] stage4_28;
   wire [5:0] stage4_29;
   wire [4:0] stage4_30;
   wire [5:0] stage4_31;
   wire [3:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [0:0] stage4_37;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [0:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [0:0] stage5_37;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[15]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_1[16]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7]},
      {stage1_6[0],stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15]}
   );
   gpc606_5 gpc16 (
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13]},
      {stage1_6[1],stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc606_5 gpc17 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage1_6[2],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc606_5 gpc18 (
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage0_4[20]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[2],stage1_6[5],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[3],stage1_6[6],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[4],stage1_6[7],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[5],stage1_6[8],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[4],stage1_7[6],stage1_6[9],stage1_5[15]}
   );
   gpc606_5 gpc25 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[5],stage1_7[7],stage1_6[10],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[6],stage1_7[8],stage1_6[11],stage1_5[17]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[7],stage1_7[9],stage1_6[12],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[8],stage1_7[10],stage1_6[13],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[9],stage1_7[11],stage1_6[14],stage1_5[20]}
   );
   gpc615_5 gpc30 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28]},
      {stage0_7[36]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[6],stage1_8[10],stage1_7[12],stage1_6[15]}
   );
   gpc615_5 gpc31 (
      {stage0_6[29], stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33]},
      {stage0_7[37]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[7],stage1_8[11],stage1_7[13],stage1_6[16]}
   );
   gpc615_5 gpc32 (
      {stage0_6[34], stage0_6[35], stage0_6[36], stage0_6[37], stage0_6[38]},
      {stage0_7[38]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[8],stage1_8[12],stage1_7[14],stage1_6[17]}
   );
   gpc606_5 gpc33 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43], stage0_7[44]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[9],stage1_8[13],stage1_7[15]}
   );
   gpc615_5 gpc34 (
      {stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49]},
      {stage0_8[18]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[10],stage1_8[14],stage1_7[16]}
   );
   gpc1163_5 gpc35 (
      {stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_10[0]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[11],stage1_8[15]}
   );
   gpc606_5 gpc36 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[12],stage1_8[16]}
   );
   gpc606_5 gpc37 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[13],stage1_8[17]}
   );
   gpc615_5 gpc38 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[18]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[14],stage1_8[18]}
   );
   gpc615_5 gpc39 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[19]},
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[15],stage1_8[19]}
   );
   gpc615_5 gpc40 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[20]},
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[16],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[17]}
   );
   gpc606_5 gpc42 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[18]}
   );
   gpc615_5 gpc43 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_10[31]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[19]}
   );
   gpc606_5 gpc44 (
      {stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[9],stage1_11[11],stage1_10[14]}
   );
   gpc606_5 gpc45 (
      {stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[10],stage1_11[12],stage1_10[15]}
   );
   gpc615_5 gpc46 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[19]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[11],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc47 (
      {stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_11[20]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[12],stage1_11[14],stage1_10[17]}
   );
   gpc606_5 gpc48 (
      {stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[4],stage1_13[7],stage1_12[13],stage1_11[15]}
   );
   gpc606_5 gpc49 (
      {stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[5],stage1_13[8],stage1_12[14],stage1_11[16]}
   );
   gpc606_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[6],stage1_13[9],stage1_12[15],stage1_11[17]}
   );
   gpc615_5 gpc51 (
      {stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43]},
      {stage0_12[24]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[7],stage1_13[10],stage1_12[16],stage1_11[18]}
   );
   gpc1423_5 gpc52 (
      {stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage0_13[24], stage0_13[25]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[4],stage1_14[8],stage1_13[11],stage1_12[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9]},
      {stage1_16[1],stage1_15[5],stage1_14[9],stage1_13[12],stage1_12[18]}
   );
   gpc606_5 gpc54 (
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage1_16[2],stage1_15[6],stage1_14[10],stage1_13[13],stage1_12[19]}
   );
   gpc606_5 gpc55 (
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21]},
      {stage1_16[3],stage1_15[7],stage1_14[11],stage1_13[14],stage1_12[20]}
   );
   gpc606_5 gpc56 (
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage1_16[4],stage1_15[8],stage1_14[12],stage1_13[15],stage1_12[21]}
   );
   gpc615_5 gpc57 (
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30]},
      {stage0_14[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[5],stage1_15[9],stage1_14[13],stage1_13[16]}
   );
   gpc615_5 gpc58 (
      {stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_14[29]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[1],stage1_16[6],stage1_15[10],stage1_14[14],stage1_13[17]}
   );
   gpc615_5 gpc59 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_14[30]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[2],stage1_16[7],stage1_15[11],stage1_14[15],stage1_13[18]}
   );
   gpc615_5 gpc60 (
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_15[19]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[8],stage1_15[12],stage1_14[16]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[20]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[9],stage1_15[13],stage1_14[17]}
   );
   gpc606_5 gpc62 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25], stage0_15[26]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[2],stage1_17[5],stage1_16[10],stage1_15[14]}
   );
   gpc606_5 gpc63 (
      {stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30], stage0_15[31], stage0_15[32]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[3],stage1_17[6],stage1_16[11],stage1_15[15]}
   );
   gpc606_5 gpc64 (
      {stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36], stage0_15[37], stage0_15[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[4],stage1_17[7],stage1_16[12],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[39], stage0_15[40], stage0_15[41], stage0_15[42], stage0_15[43]},
      {stage0_16[12]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[5],stage1_17[8],stage1_16[13],stage1_15[17]}
   );
   gpc606_5 gpc66 (
      {stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[4],stage1_18[6],stage1_17[9],stage1_16[14]}
   );
   gpc606_5 gpc67 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[5],stage1_18[7],stage1_17[10],stage1_16[15]}
   );
   gpc606_5 gpc68 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[6],stage1_18[8],stage1_17[11],stage1_16[16]}
   );
   gpc606_5 gpc69 (
      {stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[7],stage1_18[9],stage1_17[12],stage1_16[17]}
   );
   gpc606_5 gpc70 (
      {stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[8],stage1_18[10],stage1_17[13],stage1_16[18]}
   );
   gpc606_5 gpc71 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[9],stage1_18[11],stage1_17[14],stage1_16[19]}
   );
   gpc606_5 gpc72 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[6],stage1_19[10],stage1_18[12],stage1_17[15]}
   );
   gpc606_5 gpc73 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[7],stage1_19[11],stage1_18[13],stage1_17[16]}
   );
   gpc606_5 gpc74 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[8],stage1_19[12],stage1_18[14],stage1_17[17]}
   );
   gpc606_5 gpc75 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[9],stage1_19[13],stage1_18[15],stage1_17[18]}
   );
   gpc606_5 gpc76 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[10],stage1_19[14],stage1_18[16],stage1_17[19]}
   );
   gpc606_5 gpc77 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[5],stage1_20[11],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc78 (
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34]},
      {stage0_20[6]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[1],stage1_21[6],stage1_20[12],stage1_19[16]}
   );
   gpc615_5 gpc79 (
      {stage0_19[35], stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39]},
      {stage0_20[7]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[2],stage1_21[7],stage1_20[13],stage1_19[17]}
   );
   gpc606_5 gpc80 (
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[3],stage1_21[8],stage1_20[14]}
   );
   gpc606_5 gpc81 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[4],stage1_21[9],stage1_20[15]}
   );
   gpc606_5 gpc82 (
      {stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[5],stage1_21[10],stage1_20[16]}
   );
   gpc606_5 gpc83 (
      {stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[6],stage1_21[11],stage1_20[17]}
   );
   gpc606_5 gpc84 (
      {stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[7],stage1_21[12],stage1_20[18]}
   );
   gpc615_5 gpc85 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[12]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[8],stage1_21[13],stage1_20[19]}
   );
   gpc615_5 gpc86 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[13]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[9],stage1_21[14],stage1_20[20]}
   );
   gpc615_5 gpc87 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[14]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[10],stage1_21[15],stage1_20[21]}
   );
   gpc606_5 gpc88 (
      {stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[8],stage1_23[10],stage1_22[11],stage1_21[16]}
   );
   gpc606_5 gpc89 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[9],stage1_23[11],stage1_22[12],stage1_21[17]}
   );
   gpc606_5 gpc90 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[10],stage1_23[12],stage1_22[13],stage1_21[18]}
   );
   gpc606_5 gpc91 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[11],stage1_23[13],stage1_22[14],stage1_21[19]}
   );
   gpc606_5 gpc92 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[12],stage1_23[14],stage1_22[15],stage1_21[20]}
   );
   gpc606_5 gpc93 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[5],stage1_24[13],stage1_23[15]}
   );
   gpc606_5 gpc94 (
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[6],stage1_24[14],stage1_23[16]}
   );
   gpc606_5 gpc95 (
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[2],stage1_25[7],stage1_24[15]}
   );
   gpc606_5 gpc96 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[3],stage1_25[8],stage1_24[16]}
   );
   gpc606_5 gpc97 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[4],stage1_25[9],stage1_24[17]}
   );
   gpc606_5 gpc98 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[5],stage1_25[10],stage1_24[18]}
   );
   gpc606_5 gpc99 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[6],stage1_25[11],stage1_24[19]}
   );
   gpc606_5 gpc100 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[7],stage1_25[12],stage1_24[20]}
   );
   gpc606_5 gpc101 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[8],stage1_25[13],stage1_24[21]}
   );
   gpc606_5 gpc102 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[9],stage1_25[14],stage1_24[22]}
   );
   gpc606_5 gpc103 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[10],stage1_26[10],stage1_25[15],stage1_24[23]}
   );
   gpc606_5 gpc104 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[9],stage1_27[11],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc105 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[10],stage1_27[12],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc106 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[11],stage1_27[13],stage1_26[13],stage1_25[18]}
   );
   gpc606_5 gpc107 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[12],stage1_27[14],stage1_26[14],stage1_25[19]}
   );
   gpc606_5 gpc108 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[13],stage1_27[15],stage1_26[15],stage1_25[20]}
   );
   gpc606_5 gpc109 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[14],stage1_27[16],stage1_26[16],stage1_25[21]}
   );
   gpc606_5 gpc110 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[15],stage1_27[17],stage1_26[17],stage1_25[22]}
   );
   gpc606_5 gpc111 (
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[7],stage1_28[16],stage1_27[18]}
   );
   gpc606_5 gpc112 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[1],stage1_30[1],stage1_29[8],stage1_28[17]}
   );
   gpc606_5 gpc113 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[2],stage1_30[2],stage1_29[9],stage1_28[18]}
   );
   gpc606_5 gpc114 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[3],stage1_30[3],stage1_29[10],stage1_28[19]}
   );
   gpc606_5 gpc115 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[4],stage1_30[4],stage1_29[11],stage1_28[20]}
   );
   gpc606_5 gpc116 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[5],stage1_30[5],stage1_29[12],stage1_28[21]}
   );
   gpc606_5 gpc117 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[6],stage1_30[6],stage1_29[13],stage1_28[22]}
   );
   gpc606_5 gpc118 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[7],stage1_30[7],stage1_29[14],stage1_28[23]}
   );
   gpc606_5 gpc119 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[8],stage1_30[8],stage1_29[15],stage1_28[24]}
   );
   gpc606_5 gpc120 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[9],stage1_30[9],stage1_29[16],stage1_28[25]}
   );
   gpc606_5 gpc121 (
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[10],stage1_30[10],stage1_29[17]}
   );
   gpc606_5 gpc122 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[11],stage1_30[11],stage1_29[18]}
   );
   gpc606_5 gpc123 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[12],stage1_30[12],stage1_29[19]}
   );
   gpc606_5 gpc124 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[13],stage1_30[13],stage1_29[20]}
   );
   gpc606_5 gpc125 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[14],stage1_30[14],stage1_29[21]}
   );
   gpc606_5 gpc126 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[15],stage1_30[15],stage1_29[22]}
   );
   gpc606_5 gpc127 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[16],stage1_30[16],stage1_29[23]}
   );
   gpc606_5 gpc128 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[17],stage1_30[17],stage1_29[24]}
   );
   gpc1_1 gpc129 (
      {stage0_0[47]},
      {stage1_0[9]}
   );
   gpc1_1 gpc130 (
      {stage0_0[48]},
      {stage1_0[10]}
   );
   gpc1_1 gpc131 (
      {stage0_0[49]},
      {stage1_0[11]}
   );
   gpc1_1 gpc132 (
      {stage0_0[50]},
      {stage1_0[12]}
   );
   gpc1_1 gpc133 (
      {stage0_0[51]},
      {stage1_0[13]}
   );
   gpc1_1 gpc134 (
      {stage0_0[52]},
      {stage1_0[14]}
   );
   gpc1_1 gpc135 (
      {stage0_0[53]},
      {stage1_0[15]}
   );
   gpc1_1 gpc136 (
      {stage0_1[52]},
      {stage1_1[15]}
   );
   gpc1_1 gpc137 (
      {stage0_1[53]},
      {stage1_1[16]}
   );
   gpc1_1 gpc138 (
      {stage0_2[50]},
      {stage1_2[18]}
   );
   gpc1_1 gpc139 (
      {stage0_2[51]},
      {stage1_2[19]}
   );
   gpc1_1 gpc140 (
      {stage0_2[52]},
      {stage1_2[20]}
   );
   gpc1_1 gpc141 (
      {stage0_2[53]},
      {stage1_2[21]}
   );
   gpc1_1 gpc142 (
      {stage0_3[52]},
      {stage1_3[20]}
   );
   gpc1_1 gpc143 (
      {stage0_3[53]},
      {stage1_3[21]}
   );
   gpc1_1 gpc144 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc145 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc146 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc147 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc148 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc149 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc150 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc151 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc152 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc153 (
      {stage0_5[48]},
      {stage1_5[21]}
   );
   gpc1_1 gpc154 (
      {stage0_5[49]},
      {stage1_5[22]}
   );
   gpc1_1 gpc155 (
      {stage0_5[50]},
      {stage1_5[23]}
   );
   gpc1_1 gpc156 (
      {stage0_5[51]},
      {stage1_5[24]}
   );
   gpc1_1 gpc157 (
      {stage0_5[52]},
      {stage1_5[25]}
   );
   gpc1_1 gpc158 (
      {stage0_5[53]},
      {stage1_5[26]}
   );
   gpc1_1 gpc159 (
      {stage0_6[39]},
      {stage1_6[18]}
   );
   gpc1_1 gpc160 (
      {stage0_6[40]},
      {stage1_6[19]}
   );
   gpc1_1 gpc161 (
      {stage0_6[41]},
      {stage1_6[20]}
   );
   gpc1_1 gpc162 (
      {stage0_6[42]},
      {stage1_6[21]}
   );
   gpc1_1 gpc163 (
      {stage0_6[43]},
      {stage1_6[22]}
   );
   gpc1_1 gpc164 (
      {stage0_6[44]},
      {stage1_6[23]}
   );
   gpc1_1 gpc165 (
      {stage0_6[45]},
      {stage1_6[24]}
   );
   gpc1_1 gpc166 (
      {stage0_6[46]},
      {stage1_6[25]}
   );
   gpc1_1 gpc167 (
      {stage0_6[47]},
      {stage1_6[26]}
   );
   gpc1_1 gpc168 (
      {stage0_6[48]},
      {stage1_6[27]}
   );
   gpc1_1 gpc169 (
      {stage0_6[49]},
      {stage1_6[28]}
   );
   gpc1_1 gpc170 (
      {stage0_6[50]},
      {stage1_6[29]}
   );
   gpc1_1 gpc171 (
      {stage0_6[51]},
      {stage1_6[30]}
   );
   gpc1_1 gpc172 (
      {stage0_6[52]},
      {stage1_6[31]}
   );
   gpc1_1 gpc173 (
      {stage0_6[53]},
      {stage1_6[32]}
   );
   gpc1_1 gpc174 (
      {stage0_7[50]},
      {stage1_7[17]}
   );
   gpc1_1 gpc175 (
      {stage0_7[51]},
      {stage1_7[18]}
   );
   gpc1_1 gpc176 (
      {stage0_7[52]},
      {stage1_7[19]}
   );
   gpc1_1 gpc177 (
      {stage0_7[53]},
      {stage1_7[20]}
   );
   gpc1_1 gpc178 (
      {stage0_8[49]},
      {stage1_8[21]}
   );
   gpc1_1 gpc179 (
      {stage0_8[50]},
      {stage1_8[22]}
   );
   gpc1_1 gpc180 (
      {stage0_8[51]},
      {stage1_8[23]}
   );
   gpc1_1 gpc181 (
      {stage0_8[52]},
      {stage1_8[24]}
   );
   gpc1_1 gpc182 (
      {stage0_8[53]},
      {stage1_8[25]}
   );
   gpc1_1 gpc183 (
      {stage0_9[38]},
      {stage1_9[20]}
   );
   gpc1_1 gpc184 (
      {stage0_9[39]},
      {stage1_9[21]}
   );
   gpc1_1 gpc185 (
      {stage0_9[40]},
      {stage1_9[22]}
   );
   gpc1_1 gpc186 (
      {stage0_9[41]},
      {stage1_9[23]}
   );
   gpc1_1 gpc187 (
      {stage0_9[42]},
      {stage1_9[24]}
   );
   gpc1_1 gpc188 (
      {stage0_9[43]},
      {stage1_9[25]}
   );
   gpc1_1 gpc189 (
      {stage0_9[44]},
      {stage1_9[26]}
   );
   gpc1_1 gpc190 (
      {stage0_9[45]},
      {stage1_9[27]}
   );
   gpc1_1 gpc191 (
      {stage0_9[46]},
      {stage1_9[28]}
   );
   gpc1_1 gpc192 (
      {stage0_9[47]},
      {stage1_9[29]}
   );
   gpc1_1 gpc193 (
      {stage0_9[48]},
      {stage1_9[30]}
   );
   gpc1_1 gpc194 (
      {stage0_9[49]},
      {stage1_9[31]}
   );
   gpc1_1 gpc195 (
      {stage0_9[50]},
      {stage1_9[32]}
   );
   gpc1_1 gpc196 (
      {stage0_9[51]},
      {stage1_9[33]}
   );
   gpc1_1 gpc197 (
      {stage0_9[52]},
      {stage1_9[34]}
   );
   gpc1_1 gpc198 (
      {stage0_9[53]},
      {stage1_9[35]}
   );
   gpc1_1 gpc199 (
      {stage0_11[44]},
      {stage1_11[19]}
   );
   gpc1_1 gpc200 (
      {stage0_11[45]},
      {stage1_11[20]}
   );
   gpc1_1 gpc201 (
      {stage0_11[46]},
      {stage1_11[21]}
   );
   gpc1_1 gpc202 (
      {stage0_11[47]},
      {stage1_11[22]}
   );
   gpc1_1 gpc203 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc204 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc205 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc206 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc207 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc208 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc209 (
      {stage0_12[52]},
      {stage1_12[22]}
   );
   gpc1_1 gpc210 (
      {stage0_12[53]},
      {stage1_12[23]}
   );
   gpc1_1 gpc211 (
      {stage0_13[41]},
      {stage1_13[19]}
   );
   gpc1_1 gpc212 (
      {stage0_13[42]},
      {stage1_13[20]}
   );
   gpc1_1 gpc213 (
      {stage0_13[43]},
      {stage1_13[21]}
   );
   gpc1_1 gpc214 (
      {stage0_13[44]},
      {stage1_13[22]}
   );
   gpc1_1 gpc215 (
      {stage0_13[45]},
      {stage1_13[23]}
   );
   gpc1_1 gpc216 (
      {stage0_13[46]},
      {stage1_13[24]}
   );
   gpc1_1 gpc217 (
      {stage0_13[47]},
      {stage1_13[25]}
   );
   gpc1_1 gpc218 (
      {stage0_13[48]},
      {stage1_13[26]}
   );
   gpc1_1 gpc219 (
      {stage0_13[49]},
      {stage1_13[27]}
   );
   gpc1_1 gpc220 (
      {stage0_13[50]},
      {stage1_13[28]}
   );
   gpc1_1 gpc221 (
      {stage0_13[51]},
      {stage1_13[29]}
   );
   gpc1_1 gpc222 (
      {stage0_13[52]},
      {stage1_13[30]}
   );
   gpc1_1 gpc223 (
      {stage0_13[53]},
      {stage1_13[31]}
   );
   gpc1_1 gpc224 (
      {stage0_14[41]},
      {stage1_14[18]}
   );
   gpc1_1 gpc225 (
      {stage0_14[42]},
      {stage1_14[19]}
   );
   gpc1_1 gpc226 (
      {stage0_14[43]},
      {stage1_14[20]}
   );
   gpc1_1 gpc227 (
      {stage0_14[44]},
      {stage1_14[21]}
   );
   gpc1_1 gpc228 (
      {stage0_14[45]},
      {stage1_14[22]}
   );
   gpc1_1 gpc229 (
      {stage0_14[46]},
      {stage1_14[23]}
   );
   gpc1_1 gpc230 (
      {stage0_14[47]},
      {stage1_14[24]}
   );
   gpc1_1 gpc231 (
      {stage0_14[48]},
      {stage1_14[25]}
   );
   gpc1_1 gpc232 (
      {stage0_14[49]},
      {stage1_14[26]}
   );
   gpc1_1 gpc233 (
      {stage0_14[50]},
      {stage1_14[27]}
   );
   gpc1_1 gpc234 (
      {stage0_14[51]},
      {stage1_14[28]}
   );
   gpc1_1 gpc235 (
      {stage0_14[52]},
      {stage1_14[29]}
   );
   gpc1_1 gpc236 (
      {stage0_14[53]},
      {stage1_14[30]}
   );
   gpc1_1 gpc237 (
      {stage0_15[44]},
      {stage1_15[18]}
   );
   gpc1_1 gpc238 (
      {stage0_15[45]},
      {stage1_15[19]}
   );
   gpc1_1 gpc239 (
      {stage0_15[46]},
      {stage1_15[20]}
   );
   gpc1_1 gpc240 (
      {stage0_15[47]},
      {stage1_15[21]}
   );
   gpc1_1 gpc241 (
      {stage0_15[48]},
      {stage1_15[22]}
   );
   gpc1_1 gpc242 (
      {stage0_15[49]},
      {stage1_15[23]}
   );
   gpc1_1 gpc243 (
      {stage0_15[50]},
      {stage1_15[24]}
   );
   gpc1_1 gpc244 (
      {stage0_15[51]},
      {stage1_15[25]}
   );
   gpc1_1 gpc245 (
      {stage0_15[52]},
      {stage1_15[26]}
   );
   gpc1_1 gpc246 (
      {stage0_15[53]},
      {stage1_15[27]}
   );
   gpc1_1 gpc247 (
      {stage0_16[49]},
      {stage1_16[20]}
   );
   gpc1_1 gpc248 (
      {stage0_16[50]},
      {stage1_16[21]}
   );
   gpc1_1 gpc249 (
      {stage0_16[51]},
      {stage1_16[22]}
   );
   gpc1_1 gpc250 (
      {stage0_16[52]},
      {stage1_16[23]}
   );
   gpc1_1 gpc251 (
      {stage0_16[53]},
      {stage1_16[24]}
   );
   gpc1_1 gpc252 (
      {stage0_18[42]},
      {stage1_18[18]}
   );
   gpc1_1 gpc253 (
      {stage0_18[43]},
      {stage1_18[19]}
   );
   gpc1_1 gpc254 (
      {stage0_18[44]},
      {stage1_18[20]}
   );
   gpc1_1 gpc255 (
      {stage0_18[45]},
      {stage1_18[21]}
   );
   gpc1_1 gpc256 (
      {stage0_18[46]},
      {stage1_18[22]}
   );
   gpc1_1 gpc257 (
      {stage0_18[47]},
      {stage1_18[23]}
   );
   gpc1_1 gpc258 (
      {stage0_18[48]},
      {stage1_18[24]}
   );
   gpc1_1 gpc259 (
      {stage0_18[49]},
      {stage1_18[25]}
   );
   gpc1_1 gpc260 (
      {stage0_18[50]},
      {stage1_18[26]}
   );
   gpc1_1 gpc261 (
      {stage0_18[51]},
      {stage1_18[27]}
   );
   gpc1_1 gpc262 (
      {stage0_18[52]},
      {stage1_18[28]}
   );
   gpc1_1 gpc263 (
      {stage0_18[53]},
      {stage1_18[29]}
   );
   gpc1_1 gpc264 (
      {stage0_19[40]},
      {stage1_19[18]}
   );
   gpc1_1 gpc265 (
      {stage0_19[41]},
      {stage1_19[19]}
   );
   gpc1_1 gpc266 (
      {stage0_19[42]},
      {stage1_19[20]}
   );
   gpc1_1 gpc267 (
      {stage0_19[43]},
      {stage1_19[21]}
   );
   gpc1_1 gpc268 (
      {stage0_19[44]},
      {stage1_19[22]}
   );
   gpc1_1 gpc269 (
      {stage0_19[45]},
      {stage1_19[23]}
   );
   gpc1_1 gpc270 (
      {stage0_19[46]},
      {stage1_19[24]}
   );
   gpc1_1 gpc271 (
      {stage0_19[47]},
      {stage1_19[25]}
   );
   gpc1_1 gpc272 (
      {stage0_19[48]},
      {stage1_19[26]}
   );
   gpc1_1 gpc273 (
      {stage0_19[49]},
      {stage1_19[27]}
   );
   gpc1_1 gpc274 (
      {stage0_19[50]},
      {stage1_19[28]}
   );
   gpc1_1 gpc275 (
      {stage0_19[51]},
      {stage1_19[29]}
   );
   gpc1_1 gpc276 (
      {stage0_19[52]},
      {stage1_19[30]}
   );
   gpc1_1 gpc277 (
      {stage0_19[53]},
      {stage1_19[31]}
   );
   gpc1_1 gpc278 (
      {stage0_20[53]},
      {stage1_20[22]}
   );
   gpc1_1 gpc279 (
      {stage0_21[45]},
      {stage1_21[21]}
   );
   gpc1_1 gpc280 (
      {stage0_21[46]},
      {stage1_21[22]}
   );
   gpc1_1 gpc281 (
      {stage0_21[47]},
      {stage1_21[23]}
   );
   gpc1_1 gpc282 (
      {stage0_21[48]},
      {stage1_21[24]}
   );
   gpc1_1 gpc283 (
      {stage0_21[49]},
      {stage1_21[25]}
   );
   gpc1_1 gpc284 (
      {stage0_21[50]},
      {stage1_21[26]}
   );
   gpc1_1 gpc285 (
      {stage0_21[51]},
      {stage1_21[27]}
   );
   gpc1_1 gpc286 (
      {stage0_21[52]},
      {stage1_21[28]}
   );
   gpc1_1 gpc287 (
      {stage0_21[53]},
      {stage1_21[29]}
   );
   gpc1_1 gpc288 (
      {stage0_22[48]},
      {stage1_22[16]}
   );
   gpc1_1 gpc289 (
      {stage0_22[49]},
      {stage1_22[17]}
   );
   gpc1_1 gpc290 (
      {stage0_22[50]},
      {stage1_22[18]}
   );
   gpc1_1 gpc291 (
      {stage0_22[51]},
      {stage1_22[19]}
   );
   gpc1_1 gpc292 (
      {stage0_22[52]},
      {stage1_22[20]}
   );
   gpc1_1 gpc293 (
      {stage0_22[53]},
      {stage1_22[21]}
   );
   gpc1_1 gpc294 (
      {stage0_23[42]},
      {stage1_23[17]}
   );
   gpc1_1 gpc295 (
      {stage0_23[43]},
      {stage1_23[18]}
   );
   gpc1_1 gpc296 (
      {stage0_23[44]},
      {stage1_23[19]}
   );
   gpc1_1 gpc297 (
      {stage0_23[45]},
      {stage1_23[20]}
   );
   gpc1_1 gpc298 (
      {stage0_23[46]},
      {stage1_23[21]}
   );
   gpc1_1 gpc299 (
      {stage0_23[47]},
      {stage1_23[22]}
   );
   gpc1_1 gpc300 (
      {stage0_23[48]},
      {stage1_23[23]}
   );
   gpc1_1 gpc301 (
      {stage0_23[49]},
      {stage1_23[24]}
   );
   gpc1_1 gpc302 (
      {stage0_23[50]},
      {stage1_23[25]}
   );
   gpc1_1 gpc303 (
      {stage0_23[51]},
      {stage1_23[26]}
   );
   gpc1_1 gpc304 (
      {stage0_23[52]},
      {stage1_23[27]}
   );
   gpc1_1 gpc305 (
      {stage0_23[53]},
      {stage1_23[28]}
   );
   gpc1_1 gpc306 (
      {stage0_27[48]},
      {stage1_27[19]}
   );
   gpc1_1 gpc307 (
      {stage0_27[49]},
      {stage1_27[20]}
   );
   gpc1_1 gpc308 (
      {stage0_27[50]},
      {stage1_27[21]}
   );
   gpc1_1 gpc309 (
      {stage0_27[51]},
      {stage1_27[22]}
   );
   gpc1_1 gpc310 (
      {stage0_27[52]},
      {stage1_27[23]}
   );
   gpc1_1 gpc311 (
      {stage0_27[53]},
      {stage1_27[24]}
   );
   gpc1_1 gpc312 (
      {stage0_31[48]},
      {stage1_31[18]}
   );
   gpc1_1 gpc313 (
      {stage0_31[49]},
      {stage1_31[19]}
   );
   gpc1_1 gpc314 (
      {stage0_31[50]},
      {stage1_31[20]}
   );
   gpc1_1 gpc315 (
      {stage0_31[51]},
      {stage1_31[21]}
   );
   gpc1_1 gpc316 (
      {stage0_31[52]},
      {stage1_31[22]}
   );
   gpc1_1 gpc317 (
      {stage0_31[53]},
      {stage1_31[23]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc319 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[6]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc320 (
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc321 (
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc615_5 gpc322 (
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage1_4[2]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4],stage2_3[4]}
   );
   gpc606_5 gpc323 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc324 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc325 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[5],stage2_4[7]}
   );
   gpc606_5 gpc326 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[6],stage2_4[8]}
   );
   gpc606_5 gpc327 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[7],stage2_4[9]}
   );
   gpc606_5 gpc328 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[5],stage2_7[8],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc329 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc330 (
      {stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc331 (
      {stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6], stage1_8[7]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[2],stage2_9[3],stage2_8[8]}
   );
   gpc606_5 gpc332 (
      {stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[3],stage2_9[4],stage2_8[9]}
   );
   gpc606_5 gpc333 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[4],stage2_10[4],stage2_9[5],stage2_8[10]}
   );
   gpc606_5 gpc334 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[3],stage2_11[5],stage2_10[5],stage2_9[6]}
   );
   gpc606_5 gpc335 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[4],stage2_11[6],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc336 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[5],stage2_11[7],stage2_10[7],stage2_9[8]}
   );
   gpc606_5 gpc337 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[6],stage2_11[8],stage2_10[8],stage2_9[9]}
   );
   gpc615_5 gpc338 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[4],stage2_12[7],stage2_11[9]}
   );
   gpc606_5 gpc339 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[5],stage2_12[8]}
   );
   gpc606_5 gpc340 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[6],stage2_12[9]}
   );
   gpc606_5 gpc341 (
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[7],stage2_12[10]}
   );
   gpc606_5 gpc342 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[4],stage2_13[8]}
   );
   gpc606_5 gpc343 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[5],stage2_13[9]}
   );
   gpc606_5 gpc344 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[6],stage2_13[10]}
   );
   gpc1163_5 gpc345 (
      {stage1_14[18], stage1_14[19], stage1_14[20]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[7]}
   );
   gpc615_5 gpc346 (
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage1_15[24]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[1],stage2_17[4],stage2_16[7],stage2_15[8],stage2_14[8]}
   );
   gpc615_5 gpc347 (
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage1_15[25]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[2],stage2_17[5],stage2_16[8],stage2_15[9],stage2_14[9]}
   );
   gpc606_5 gpc348 (
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[3],stage2_17[6],stage2_16[9]}
   );
   gpc606_5 gpc349 (
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[4],stage2_17[7],stage2_16[10]}
   );
   gpc606_5 gpc350 (
      {stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[5],stage2_17[8]}
   );
   gpc606_5 gpc351 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[6],stage2_17[9]}
   );
   gpc606_5 gpc352 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[7],stage2_17[10]}
   );
   gpc615_5 gpc353 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16]},
      {stage1_19[18]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[8]}
   );
   gpc615_5 gpc354 (
      {stage1_18[17], stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21]},
      {stage1_19[19]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[9]}
   );
   gpc615_5 gpc355 (
      {stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26]},
      {stage1_19[20]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[10]}
   );
   gpc606_5 gpc356 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25], stage1_19[26]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[6],stage2_20[8],stage2_19[8]}
   );
   gpc606_5 gpc357 (
      {stage1_19[27], stage1_19[28], stage1_19[29], stage1_19[30], stage1_19[31], 1'b0},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[7],stage2_20[9],stage2_19[9]}
   );
   gpc606_5 gpc358 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], 1'b0},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[2],stage2_22[5],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc359 (
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[3],stage2_22[6],stage2_21[9]}
   );
   gpc606_5 gpc360 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[4],stage2_22[7],stage2_21[10]}
   );
   gpc606_5 gpc361 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[5],stage2_22[8],stage2_21[11]}
   );
   gpc615_5 gpc362 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10]},
      {stage1_23[18]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[3],stage2_24[4],stage2_23[6],stage2_22[9]}
   );
   gpc615_5 gpc363 (
      {stage1_22[11], stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15]},
      {stage1_23[19]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[4],stage2_24[5],stage2_23[7],stage2_22[10]}
   );
   gpc1415_5 gpc364 (
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4]},
      {stage1_26[0]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3]},
      {stage1_28[0]},
      {stage2_29[0],stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[5]}
   );
   gpc615_5 gpc365 (
      {stage1_25[5], stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9]},
      {stage1_26[1]},
      {stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage2_29[1],stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[6]}
   );
   gpc615_5 gpc366 (
      {stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13], stage1_25[14]},
      {stage1_26[2]},
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15]},
      {stage2_29[2],stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[7]}
   );
   gpc615_5 gpc367 (
      {stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18], stage1_25[19]},
      {stage1_26[3]},
      {stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21]},
      {stage2_29[3],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[8]}
   );
   gpc615_5 gpc368 (
      {stage1_26[4], stage1_26[5], stage1_26[6], stage1_26[7], stage1_26[8]},
      {stage1_27[22]},
      {stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5], stage1_28[6]},
      {stage2_30[0],stage2_29[4],stage2_28[4],stage2_27[4],stage2_26[6]}
   );
   gpc615_5 gpc369 (
      {stage1_26[9], stage1_26[10], stage1_26[11], stage1_26[12], stage1_26[13]},
      {stage1_27[23]},
      {stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12]},
      {stage2_30[1],stage2_29[5],stage2_28[5],stage2_27[5],stage2_26[7]}
   );
   gpc615_5 gpc370 (
      {stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17], 1'b0},
      {stage1_27[24]},
      {stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18]},
      {stage2_30[2],stage2_29[6],stage2_28[6],stage2_27[6],stage2_26[8]}
   );
   gpc2135_5 gpc371 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage1_32[0], stage1_32[1]},
      {stage2_33[0],stage2_32[0],stage2_31[0],stage2_30[3],stage2_29[7]}
   );
   gpc1406_5 gpc372 (
      {stage1_29[5], stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10]},
      {stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4]},
      {stage1_32[2]},
      {stage2_33[1],stage2_32[1],stage2_31[1],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc373 (
      {stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10]},
      {stage2_33[2],stage2_32[2],stage2_31[2],stage2_30[5],stage2_29[9]}
   );
   gpc606_5 gpc374 (
      {stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8]},
      {stage2_34[0],stage2_33[3],stage2_32[3],stage2_31[3],stage2_30[6]}
   );
   gpc606_5 gpc375 (
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14]},
      {stage2_34[1],stage2_33[4],stage2_32[4],stage2_31[4],stage2_30[7]}
   );
   gpc615_5 gpc376 (
      {stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_32[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[5],stage2_32[5],stage2_31[5]}
   );
   gpc615_5 gpc377 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20]},
      {stage1_32[16]},
      {stage1_33[6], stage1_33[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_35[1],stage2_34[3],stage2_33[6],stage2_32[6],stage2_31[6]}
   );
   gpc1_1 gpc378 (
      {stage1_0[8]},
      {stage2_0[2]}
   );
   gpc1_1 gpc379 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc380 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc381 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc382 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc383 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc384 (
      {stage1_0[14]},
      {stage2_0[8]}
   );
   gpc1_1 gpc385 (
      {stage1_0[15]},
      {stage2_0[9]}
   );
   gpc1_1 gpc386 (
      {stage1_1[7]},
      {stage2_1[2]}
   );
   gpc1_1 gpc387 (
      {stage1_1[8]},
      {stage2_1[3]}
   );
   gpc1_1 gpc388 (
      {stage1_1[9]},
      {stage2_1[4]}
   );
   gpc1_1 gpc389 (
      {stage1_1[10]},
      {stage2_1[5]}
   );
   gpc1_1 gpc390 (
      {stage1_1[11]},
      {stage2_1[6]}
   );
   gpc1_1 gpc391 (
      {stage1_1[12]},
      {stage2_1[7]}
   );
   gpc1_1 gpc392 (
      {stage1_1[13]},
      {stage2_1[8]}
   );
   gpc1_1 gpc393 (
      {stage1_1[14]},
      {stage2_1[9]}
   );
   gpc1_1 gpc394 (
      {stage1_1[15]},
      {stage2_1[10]}
   );
   gpc1_1 gpc395 (
      {stage1_1[16]},
      {stage2_1[11]}
   );
   gpc1_1 gpc396 (
      {stage1_2[7]},
      {stage2_2[2]}
   );
   gpc1_1 gpc397 (
      {stage1_2[8]},
      {stage2_2[3]}
   );
   gpc1_1 gpc398 (
      {stage1_2[9]},
      {stage2_2[4]}
   );
   gpc1_1 gpc399 (
      {stage1_2[10]},
      {stage2_2[5]}
   );
   gpc1_1 gpc400 (
      {stage1_2[11]},
      {stage2_2[6]}
   );
   gpc1_1 gpc401 (
      {stage1_2[12]},
      {stage2_2[7]}
   );
   gpc1_1 gpc402 (
      {stage1_2[13]},
      {stage2_2[8]}
   );
   gpc1_1 gpc403 (
      {stage1_2[14]},
      {stage2_2[9]}
   );
   gpc1_1 gpc404 (
      {stage1_2[15]},
      {stage2_2[10]}
   );
   gpc1_1 gpc405 (
      {stage1_2[16]},
      {stage2_2[11]}
   );
   gpc1_1 gpc406 (
      {stage1_2[17]},
      {stage2_2[12]}
   );
   gpc1_1 gpc407 (
      {stage1_2[18]},
      {stage2_2[13]}
   );
   gpc1_1 gpc408 (
      {stage1_2[19]},
      {stage2_2[14]}
   );
   gpc1_1 gpc409 (
      {stage1_2[20]},
      {stage2_2[15]}
   );
   gpc1_1 gpc410 (
      {stage1_2[21]},
      {stage2_2[16]}
   );
   gpc1_1 gpc411 (
      {stage1_3[16]},
      {stage2_3[5]}
   );
   gpc1_1 gpc412 (
      {stage1_3[17]},
      {stage2_3[6]}
   );
   gpc1_1 gpc413 (
      {stage1_3[18]},
      {stage2_3[7]}
   );
   gpc1_1 gpc414 (
      {stage1_3[19]},
      {stage2_3[8]}
   );
   gpc1_1 gpc415 (
      {stage1_3[20]},
      {stage2_3[9]}
   );
   gpc1_1 gpc416 (
      {stage1_3[21]},
      {stage2_3[10]}
   );
   gpc1_1 gpc417 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc418 (
      {stage1_5[25]},
      {stage2_5[10]}
   );
   gpc1_1 gpc419 (
      {stage1_5[26]},
      {stage2_5[11]}
   );
   gpc1_1 gpc420 (
      {stage1_6[30]},
      {stage2_6[9]}
   );
   gpc1_1 gpc421 (
      {stage1_6[31]},
      {stage2_6[10]}
   );
   gpc1_1 gpc422 (
      {stage1_6[32]},
      {stage2_6[11]}
   );
   gpc1_1 gpc423 (
      {stage1_7[16]},
      {stage2_7[11]}
   );
   gpc1_1 gpc424 (
      {stage1_7[17]},
      {stage2_7[12]}
   );
   gpc1_1 gpc425 (
      {stage1_7[18]},
      {stage2_7[13]}
   );
   gpc1_1 gpc426 (
      {stage1_7[19]},
      {stage2_7[14]}
   );
   gpc1_1 gpc427 (
      {stage1_7[20]},
      {stage2_7[15]}
   );
   gpc1_1 gpc428 (
      {stage1_8[20]},
      {stage2_8[11]}
   );
   gpc1_1 gpc429 (
      {stage1_8[21]},
      {stage2_8[12]}
   );
   gpc1_1 gpc430 (
      {stage1_8[22]},
      {stage2_8[13]}
   );
   gpc1_1 gpc431 (
      {stage1_8[23]},
      {stage2_8[14]}
   );
   gpc1_1 gpc432 (
      {stage1_8[24]},
      {stage2_8[15]}
   );
   gpc1_1 gpc433 (
      {stage1_8[25]},
      {stage2_8[16]}
   );
   gpc1_1 gpc434 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc435 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc436 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc437 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc438 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc439 (
      {stage1_13[24]},
      {stage2_13[11]}
   );
   gpc1_1 gpc440 (
      {stage1_13[25]},
      {stage2_13[12]}
   );
   gpc1_1 gpc441 (
      {stage1_13[26]},
      {stage2_13[13]}
   );
   gpc1_1 gpc442 (
      {stage1_13[27]},
      {stage2_13[14]}
   );
   gpc1_1 gpc443 (
      {stage1_13[28]},
      {stage2_13[15]}
   );
   gpc1_1 gpc444 (
      {stage1_13[29]},
      {stage2_13[16]}
   );
   gpc1_1 gpc445 (
      {stage1_13[30]},
      {stage2_13[17]}
   );
   gpc1_1 gpc446 (
      {stage1_13[31]},
      {stage2_13[18]}
   );
   gpc1_1 gpc447 (
      {stage1_15[26]},
      {stage2_15[10]}
   );
   gpc1_1 gpc448 (
      {stage1_15[27]},
      {stage2_15[11]}
   );
   gpc1_1 gpc449 (
      {stage1_17[19]},
      {stage2_17[11]}
   );
   gpc1_1 gpc450 (
      {stage1_18[27]},
      {stage2_18[11]}
   );
   gpc1_1 gpc451 (
      {stage1_18[28]},
      {stage2_18[12]}
   );
   gpc1_1 gpc452 (
      {stage1_18[29]},
      {stage2_18[13]}
   );
   gpc1_1 gpc453 (
      {stage1_22[16]},
      {stage2_22[11]}
   );
   gpc1_1 gpc454 (
      {stage1_22[17]},
      {stage2_22[12]}
   );
   gpc1_1 gpc455 (
      {stage1_22[18]},
      {stage2_22[13]}
   );
   gpc1_1 gpc456 (
      {stage1_22[19]},
      {stage2_22[14]}
   );
   gpc1_1 gpc457 (
      {stage1_22[20]},
      {stage2_22[15]}
   );
   gpc1_1 gpc458 (
      {stage1_22[21]},
      {stage2_22[16]}
   );
   gpc1_1 gpc459 (
      {stage1_23[20]},
      {stage2_23[8]}
   );
   gpc1_1 gpc460 (
      {stage1_23[21]},
      {stage2_23[9]}
   );
   gpc1_1 gpc461 (
      {stage1_23[22]},
      {stage2_23[10]}
   );
   gpc1_1 gpc462 (
      {stage1_23[23]},
      {stage2_23[11]}
   );
   gpc1_1 gpc463 (
      {stage1_23[24]},
      {stage2_23[12]}
   );
   gpc1_1 gpc464 (
      {stage1_23[25]},
      {stage2_23[13]}
   );
   gpc1_1 gpc465 (
      {stage1_23[26]},
      {stage2_23[14]}
   );
   gpc1_1 gpc466 (
      {stage1_23[27]},
      {stage2_23[15]}
   );
   gpc1_1 gpc467 (
      {stage1_23[28]},
      {stage2_23[16]}
   );
   gpc1_1 gpc468 (
      {stage1_24[12]},
      {stage2_24[6]}
   );
   gpc1_1 gpc469 (
      {stage1_24[13]},
      {stage2_24[7]}
   );
   gpc1_1 gpc470 (
      {stage1_24[14]},
      {stage2_24[8]}
   );
   gpc1_1 gpc471 (
      {stage1_24[15]},
      {stage2_24[9]}
   );
   gpc1_1 gpc472 (
      {stage1_24[16]},
      {stage2_24[10]}
   );
   gpc1_1 gpc473 (
      {stage1_24[17]},
      {stage2_24[11]}
   );
   gpc1_1 gpc474 (
      {stage1_24[18]},
      {stage2_24[12]}
   );
   gpc1_1 gpc475 (
      {stage1_24[19]},
      {stage2_24[13]}
   );
   gpc1_1 gpc476 (
      {stage1_24[20]},
      {stage2_24[14]}
   );
   gpc1_1 gpc477 (
      {stage1_24[21]},
      {stage2_24[15]}
   );
   gpc1_1 gpc478 (
      {stage1_24[22]},
      {stage2_24[16]}
   );
   gpc1_1 gpc479 (
      {stage1_24[23]},
      {stage2_24[17]}
   );
   gpc1_1 gpc480 (
      {stage1_25[20]},
      {stage2_25[9]}
   );
   gpc1_1 gpc481 (
      {stage1_25[21]},
      {stage2_25[10]}
   );
   gpc1_1 gpc482 (
      {stage1_25[22]},
      {stage2_25[11]}
   );
   gpc1_1 gpc483 (
      {stage1_28[19]},
      {stage2_28[7]}
   );
   gpc1_1 gpc484 (
      {stage1_28[20]},
      {stage2_28[8]}
   );
   gpc1_1 gpc485 (
      {stage1_28[21]},
      {stage2_28[9]}
   );
   gpc1_1 gpc486 (
      {stage1_28[22]},
      {stage2_28[10]}
   );
   gpc1_1 gpc487 (
      {stage1_28[23]},
      {stage2_28[11]}
   );
   gpc1_1 gpc488 (
      {stage1_28[24]},
      {stage2_28[12]}
   );
   gpc1_1 gpc489 (
      {stage1_28[25]},
      {stage2_28[13]}
   );
   gpc1_1 gpc490 (
      {stage1_29[17]},
      {stage2_29[10]}
   );
   gpc1_1 gpc491 (
      {stage1_29[18]},
      {stage2_29[11]}
   );
   gpc1_1 gpc492 (
      {stage1_29[19]},
      {stage2_29[12]}
   );
   gpc1_1 gpc493 (
      {stage1_29[20]},
      {stage2_29[13]}
   );
   gpc1_1 gpc494 (
      {stage1_29[21]},
      {stage2_29[14]}
   );
   gpc1_1 gpc495 (
      {stage1_29[22]},
      {stage2_29[15]}
   );
   gpc1_1 gpc496 (
      {stage1_29[23]},
      {stage2_29[16]}
   );
   gpc1_1 gpc497 (
      {stage1_29[24]},
      {stage2_29[17]}
   );
   gpc1_1 gpc498 (
      {stage1_30[15]},
      {stage2_30[8]}
   );
   gpc1_1 gpc499 (
      {stage1_30[16]},
      {stage2_30[9]}
   );
   gpc1_1 gpc500 (
      {stage1_30[17]},
      {stage2_30[10]}
   );
   gpc1_1 gpc501 (
      {stage1_31[21]},
      {stage2_31[7]}
   );
   gpc1_1 gpc502 (
      {stage1_31[22]},
      {stage2_31[8]}
   );
   gpc1_1 gpc503 (
      {stage1_31[23]},
      {stage2_31[9]}
   );
   gpc615_5 gpc504 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc505 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc506 (
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc507 (
      {stage2_4[6], stage2_4[7], stage2_4[8]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0]},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc606_5 gpc508 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[2]}
   );
   gpc606_5 gpc509 (
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[2],stage3_7[2],stage3_6[3]}
   );
   gpc606_5 gpc510 (
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], 1'b0},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[3],stage3_7[3],stage3_6[4]}
   );
   gpc615_5 gpc511 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[3],stage3_8[4],stage3_7[4]}
   );
   gpc606_5 gpc512 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[3]}
   );
   gpc615_5 gpc513 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[1],stage3_11[2]}
   );
   gpc615_5 gpc514 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage2_12[7]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[2],stage3_11[3]}
   );
   gpc606_5 gpc515 (
      {stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[3],stage3_13[3],stage3_12[3]}
   );
   gpc135_4 gpc516 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16]},
      {stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage2_15[0]},
      {stage3_16[1],stage3_15[3],stage3_14[4],stage3_13[4]}
   );
   gpc606_5 gpc517 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[4]}
   );
   gpc615_5 gpc518 (
      {stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[1],stage3_17[1],stage3_16[3],stage3_15[5]}
   );
   gpc606_5 gpc519 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[2],stage3_17[2],stage3_16[4]}
   );
   gpc1343_5 gpc520 (
      {stage2_18[6], stage2_18[7], stage2_18[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[3]}
   );
   gpc1343_5 gpc521 (
      {stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[4]}
   );
   gpc606_5 gpc522 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[2]}
   );
   gpc615_5 gpc523 (
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4]},
      {stage2_23[6]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3]}
   );
   gpc615_5 gpc524 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9]},
      {stage2_23[7]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4]}
   );
   gpc615_5 gpc525 (
      {stage2_22[10], stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14]},
      {stage2_23[8]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5]}
   );
   gpc606_5 gpc526 (
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[3],stage3_25[4],stage3_24[4],stage3_23[4]}
   );
   gpc606_5 gpc527 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[1],stage3_26[4],stage3_25[5]}
   );
   gpc1415_5 gpc528 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4]},
      {stage2_27[6]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[1],stage3_28[1],stage3_27[2],stage3_26[5]}
   );
   gpc615_5 gpc529 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[1]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[2],stage3_28[2]}
   );
   gpc615_5 gpc530 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[2]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], 1'b0},
      {stage3_32[1],stage3_31[1],stage3_30[2],stage3_29[3],stage3_28[3]}
   );
   gpc606_5 gpc531 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[2],stage3_31[2]}
   );
   gpc117_4 gpc532 (
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5], stage2_32[6]},
      {stage2_33[6]},
      {stage2_34[0]},
      {stage3_35[1],stage3_34[1],stage3_33[1],stage3_32[3]}
   );
   gpc1_1 gpc533 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc534 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc535 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc536 (
      {stage2_1[5]},
      {stage3_1[5]}
   );
   gpc1_1 gpc537 (
      {stage2_1[6]},
      {stage3_1[6]}
   );
   gpc1_1 gpc538 (
      {stage2_1[7]},
      {stage3_1[7]}
   );
   gpc1_1 gpc539 (
      {stage2_1[8]},
      {stage3_1[8]}
   );
   gpc1_1 gpc540 (
      {stage2_1[9]},
      {stage3_1[9]}
   );
   gpc1_1 gpc541 (
      {stage2_1[10]},
      {stage3_1[10]}
   );
   gpc1_1 gpc542 (
      {stage2_1[11]},
      {stage3_1[11]}
   );
   gpc1_1 gpc543 (
      {stage2_3[1]},
      {stage3_3[3]}
   );
   gpc1_1 gpc544 (
      {stage2_3[2]},
      {stage3_3[4]}
   );
   gpc1_1 gpc545 (
      {stage2_3[3]},
      {stage3_3[5]}
   );
   gpc1_1 gpc546 (
      {stage2_3[4]},
      {stage3_3[6]}
   );
   gpc1_1 gpc547 (
      {stage2_3[5]},
      {stage3_3[7]}
   );
   gpc1_1 gpc548 (
      {stage2_3[6]},
      {stage3_3[8]}
   );
   gpc1_1 gpc549 (
      {stage2_3[7]},
      {stage3_3[9]}
   );
   gpc1_1 gpc550 (
      {stage2_3[8]},
      {stage3_3[10]}
   );
   gpc1_1 gpc551 (
      {stage2_3[9]},
      {stage3_3[11]}
   );
   gpc1_1 gpc552 (
      {stage2_3[10]},
      {stage3_3[12]}
   );
   gpc1_1 gpc553 (
      {stage2_4[9]},
      {stage3_4[4]}
   );
   gpc1_1 gpc554 (
      {stage2_7[12]},
      {stage3_7[5]}
   );
   gpc1_1 gpc555 (
      {stage2_7[13]},
      {stage3_7[6]}
   );
   gpc1_1 gpc556 (
      {stage2_7[14]},
      {stage3_7[7]}
   );
   gpc1_1 gpc557 (
      {stage2_7[15]},
      {stage3_7[8]}
   );
   gpc1_1 gpc558 (
      {stage2_8[13]},
      {stage3_8[5]}
   );
   gpc1_1 gpc559 (
      {stage2_8[14]},
      {stage3_8[6]}
   );
   gpc1_1 gpc560 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc561 (
      {stage2_8[16]},
      {stage3_8[8]}
   );
   gpc1_1 gpc562 (
      {stage2_9[6]},
      {stage3_9[4]}
   );
   gpc1_1 gpc563 (
      {stage2_9[7]},
      {stage3_9[5]}
   );
   gpc1_1 gpc564 (
      {stage2_9[8]},
      {stage3_9[6]}
   );
   gpc1_1 gpc565 (
      {stage2_9[9]},
      {stage3_9[7]}
   );
   gpc1_1 gpc566 (
      {stage2_10[6]},
      {stage3_10[4]}
   );
   gpc1_1 gpc567 (
      {stage2_10[7]},
      {stage3_10[5]}
   );
   gpc1_1 gpc568 (
      {stage2_10[8]},
      {stage3_10[6]}
   );
   gpc1_1 gpc569 (
      {stage2_12[14]},
      {stage3_12[4]}
   );
   gpc1_1 gpc570 (
      {stage2_12[15]},
      {stage3_12[5]}
   );
   gpc1_1 gpc571 (
      {stage2_13[17]},
      {stage3_13[5]}
   );
   gpc1_1 gpc572 (
      {stage2_13[18]},
      {stage3_13[6]}
   );
   gpc1_1 gpc573 (
      {stage2_14[9]},
      {stage3_14[5]}
   );
   gpc1_1 gpc574 (
      {stage2_16[7]},
      {stage3_16[5]}
   );
   gpc1_1 gpc575 (
      {stage2_16[8]},
      {stage3_16[6]}
   );
   gpc1_1 gpc576 (
      {stage2_16[9]},
      {stage3_16[7]}
   );
   gpc1_1 gpc577 (
      {stage2_16[10]},
      {stage3_16[8]}
   );
   gpc1_1 gpc578 (
      {stage2_18[12]},
      {stage3_18[5]}
   );
   gpc1_1 gpc579 (
      {stage2_18[13]},
      {stage3_18[6]}
   );
   gpc1_1 gpc580 (
      {stage2_19[8]},
      {stage3_19[5]}
   );
   gpc1_1 gpc581 (
      {stage2_19[9]},
      {stage3_19[6]}
   );
   gpc1_1 gpc582 (
      {stage2_20[6]},
      {stage3_20[3]}
   );
   gpc1_1 gpc583 (
      {stage2_20[7]},
      {stage3_20[4]}
   );
   gpc1_1 gpc584 (
      {stage2_20[8]},
      {stage3_20[5]}
   );
   gpc1_1 gpc585 (
      {stage2_20[9]},
      {stage3_20[6]}
   );
   gpc1_1 gpc586 (
      {stage2_20[10]},
      {stage3_20[7]}
   );
   gpc1_1 gpc587 (
      {stage2_21[8]},
      {stage3_21[3]}
   );
   gpc1_1 gpc588 (
      {stage2_21[9]},
      {stage3_21[4]}
   );
   gpc1_1 gpc589 (
      {stage2_21[10]},
      {stage3_21[5]}
   );
   gpc1_1 gpc590 (
      {stage2_21[11]},
      {stage3_21[6]}
   );
   gpc1_1 gpc591 (
      {stage2_22[15]},
      {stage3_22[6]}
   );
   gpc1_1 gpc592 (
      {stage2_22[16]},
      {stage3_22[7]}
   );
   gpc1_1 gpc593 (
      {stage2_23[15]},
      {stage3_23[5]}
   );
   gpc1_1 gpc594 (
      {stage2_23[16]},
      {stage3_23[6]}
   );
   gpc1_1 gpc595 (
      {stage2_26[5]},
      {stage3_26[6]}
   );
   gpc1_1 gpc596 (
      {stage2_26[6]},
      {stage3_26[7]}
   );
   gpc1_1 gpc597 (
      {stage2_26[7]},
      {stage3_26[8]}
   );
   gpc1_1 gpc598 (
      {stage2_26[8]},
      {stage3_26[9]}
   );
   gpc1_1 gpc599 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc600 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc601 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc602 (
      {stage2_29[6]},
      {stage3_29[7]}
   );
   gpc1_1 gpc603 (
      {stage2_29[7]},
      {stage3_29[8]}
   );
   gpc1_1 gpc604 (
      {stage2_29[8]},
      {stage3_29[9]}
   );
   gpc1_1 gpc605 (
      {stage2_29[9]},
      {stage3_29[10]}
   );
   gpc1_1 gpc606 (
      {stage2_29[10]},
      {stage3_29[11]}
   );
   gpc1_1 gpc607 (
      {stage2_29[11]},
      {stage3_29[12]}
   );
   gpc1_1 gpc608 (
      {stage2_29[12]},
      {stage3_29[13]}
   );
   gpc1_1 gpc609 (
      {stage2_29[13]},
      {stage3_29[14]}
   );
   gpc1_1 gpc610 (
      {stage2_29[14]},
      {stage3_29[15]}
   );
   gpc1_1 gpc611 (
      {stage2_29[15]},
      {stage3_29[16]}
   );
   gpc1_1 gpc612 (
      {stage2_29[16]},
      {stage3_29[17]}
   );
   gpc1_1 gpc613 (
      {stage2_29[17]},
      {stage3_29[18]}
   );
   gpc1_1 gpc614 (
      {stage2_31[6]},
      {stage3_31[3]}
   );
   gpc1_1 gpc615 (
      {stage2_31[7]},
      {stage3_31[4]}
   );
   gpc1_1 gpc616 (
      {stage2_31[8]},
      {stage3_31[5]}
   );
   gpc1_1 gpc617 (
      {stage2_31[9]},
      {stage3_31[6]}
   );
   gpc1_1 gpc618 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1_1 gpc619 (
      {stage2_34[2]},
      {stage3_34[3]}
   );
   gpc1_1 gpc620 (
      {stage2_34[3]},
      {stage3_34[4]}
   );
   gpc1_1 gpc621 (
      {stage2_35[0]},
      {stage3_35[2]}
   );
   gpc1_1 gpc622 (
      {stage2_35[1]},
      {stage3_35[3]}
   );
   gpc615_5 gpc623 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4]},
      {stage3_2[0]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc624 (
      {stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9]},
      {stage3_2[1]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc2135_5 gpc625 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[2]}
   );
   gpc623_5 gpc626 (
      {stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1]}
   );
   gpc615_5 gpc627 (
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[2]}
   );
   gpc615_5 gpc628 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[2]}
   );
   gpc623_5 gpc629 (
      {stage3_11[1], stage3_11[2], stage3_11[3]},
      {1'b0, 1'b0},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1],stage4_11[2]}
   );
   gpc1406_5 gpc630 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[2]}
   );
   gpc215_4 gpc631 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[4]},
      {stage3_17[1], stage3_17[2]},
      {stage4_18[1],stage4_17[1],stage4_16[1],stage4_15[2]}
   );
   gpc606_5 gpc632 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[2]}
   );
   gpc117_4 gpc633 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_20[6]},
      {stage3_21[0]},
      {stage4_22[1],stage4_21[1],stage4_20[1],stage4_19[1]}
   );
   gpc606_5 gpc634 (
      {stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[0],stage4_23[0],stage4_22[2],stage4_21[2]}
   );
   gpc606_5 gpc635 (
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], 1'b0},
      {stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[1],stage4_22[3]}
   );
   gpc1343_5 gpc636 (
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3]},
      {stage3_27[0], stage3_27[1], stage3_27[2]},
      {stage3_28[0]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[1],stage4_25[2]}
   );
   gpc135_4 gpc637 (
      {stage3_28[1], stage3_28[2], stage3_28[3], 1'b0, 1'b0},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[1]}
   );
   gpc207_4 gpc638 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[2]}
   );
   gpc207_4 gpc639 (
      {stage3_29[10], stage3_29[11], stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc623_5 gpc640 (
      {stage3_32[0], stage3_32[1], stage3_32[2]},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], 1'b0},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[2]}
   );
   gpc215_4 gpc641 (
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], 1'b0},
      {1'b0},
      {1'b0, 1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[1]}
   );
   gpc1_1 gpc642 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc643 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc644 (
      {stage3_1[10]},
      {stage4_1[2]}
   );
   gpc1_1 gpc645 (
      {stage3_1[11]},
      {stage4_1[3]}
   );
   gpc1_1 gpc646 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc647 (
      {stage3_3[12]},
      {stage4_3[2]}
   );
   gpc1_1 gpc648 (
      {stage3_6[4]},
      {stage4_6[2]}
   );
   gpc1_1 gpc649 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc650 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc651 (
      {stage3_9[6]},
      {stage4_9[2]}
   );
   gpc1_1 gpc652 (
      {stage3_9[7]},
      {stage4_9[3]}
   );
   gpc1_1 gpc653 (
      {stage3_10[5]},
      {stage4_10[3]}
   );
   gpc1_1 gpc654 (
      {stage3_10[6]},
      {stage4_10[4]}
   );
   gpc1_1 gpc655 (
      {stage3_13[6]},
      {stage4_13[2]}
   );
   gpc1_1 gpc656 (
      {stage3_15[5]},
      {stage4_15[3]}
   );
   gpc1_1 gpc657 (
      {stage3_16[5]},
      {stage4_16[2]}
   );
   gpc1_1 gpc658 (
      {stage3_16[6]},
      {stage4_16[3]}
   );
   gpc1_1 gpc659 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc660 (
      {stage3_16[8]},
      {stage4_16[5]}
   );
   gpc1_1 gpc661 (
      {stage3_18[6]},
      {stage4_18[3]}
   );
   gpc1_1 gpc662 (
      {stage3_20[7]},
      {stage4_20[2]}
   );
   gpc1_1 gpc663 (
      {stage3_22[6]},
      {stage4_22[4]}
   );
   gpc1_1 gpc664 (
      {stage3_22[7]},
      {stage4_22[5]}
   );
   gpc1_1 gpc665 (
      {stage3_23[6]},
      {stage4_23[2]}
   );
   gpc1_1 gpc666 (
      {stage3_25[3]},
      {stage4_25[3]}
   );
   gpc1_1 gpc667 (
      {stage3_25[4]},
      {stage4_25[4]}
   );
   gpc1_1 gpc668 (
      {stage3_25[5]},
      {stage4_25[5]}
   );
   gpc1_1 gpc669 (
      {stage3_26[4]},
      {stage4_26[2]}
   );
   gpc1_1 gpc670 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc671 (
      {stage3_26[6]},
      {stage4_26[4]}
   );
   gpc1_1 gpc672 (
      {stage3_26[7]},
      {stage4_26[5]}
   );
   gpc1_1 gpc673 (
      {stage3_26[8]},
      {stage4_26[6]}
   );
   gpc1_1 gpc674 (
      {stage3_26[9]},
      {stage4_26[7]}
   );
   gpc1_1 gpc675 (
      {stage3_29[17]},
      {stage4_29[4]}
   );
   gpc1_1 gpc676 (
      {stage3_29[18]},
      {stage4_29[5]}
   );
   gpc1_1 gpc677 (
      {stage3_30[1]},
      {stage4_30[3]}
   );
   gpc1_1 gpc678 (
      {stage3_30[2]},
      {stage4_30[4]}
   );
   gpc1_1 gpc679 (
      {stage3_31[4]},
      {stage4_31[3]}
   );
   gpc1_1 gpc680 (
      {stage3_31[5]},
      {stage4_31[4]}
   );
   gpc1_1 gpc681 (
      {stage3_31[6]},
      {stage4_31[5]}
   );
   gpc1_1 gpc682 (
      {stage3_32[3]},
      {stage4_32[3]}
   );
   gpc23_3 gpc683 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc2223_5 gpc684 (
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1]},
      {stage4_5[0], stage4_5[1]},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[1]}
   );
   gpc1343_5 gpc685 (
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1]}
   );
   gpc135_4 gpc686 (
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], 1'b0},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1423_5 gpc687 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc1325_5 gpc688 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0], stage4_17[1]},
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc689 (
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0], stage4_21[1], stage4_21[2], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1]}
   );
   gpc223_4 gpc690 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[1],stage5_23[1],stage5_22[1]}
   );
   gpc2116_5 gpc691 (
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage4_26[0]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1]}
   );
   gpc7_3 gpc692 (
      {stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage5_28[1],stage5_27[1],stage5_26[1]}
   );
   gpc606_5 gpc693 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[0],stage5_29[1]}
   );
   gpc1415_5 gpc694 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4]},
      {1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[1]}
   );
   gpc1_1 gpc695 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc696 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc697 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc698 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc699 (
      {stage4_4[2]},
      {stage5_4[1]}
   );
   gpc1_1 gpc700 (
      {stage4_5[2]},
      {stage5_5[1]}
   );
   gpc1_1 gpc701 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc702 (
      {stage4_8[4]},
      {stage5_8[1]}
   );
   gpc1_1 gpc703 (
      {stage4_9[3]},
      {stage5_9[1]}
   );
   gpc1_1 gpc704 (
      {stage4_12[1]},
      {stage5_12[1]}
   );
   gpc1_1 gpc705 (
      {stage4_14[2]},
      {stage5_14[1]}
   );
   gpc1_1 gpc706 (
      {stage4_18[3]},
      {stage5_18[1]}
   );
   gpc1_1 gpc707 (
      {stage4_19[1]},
      {stage5_19[1]}
   );
   gpc1_1 gpc708 (
      {stage4_34[0]},
      {stage5_34[1]}
   );
   gpc1_1 gpc709 (
      {stage4_35[0]},
      {stage5_35[0]}
   );
   gpc1_1 gpc710 (
      {stage4_35[1]},
      {stage5_35[1]}
   );
   gpc1_1 gpc711 (
      {stage4_36[0]},
      {stage5_36[0]}
   );
   gpc1_1 gpc712 (
      {stage4_36[1]},
      {stage5_36[1]}
   );
   gpc1_1 gpc713 (
      {stage4_37[0]},
      {stage5_37[0]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor_CLA54_32 compressor_CLA54_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hca332cab7e8b10cf819bb5a39cbf55f830b512395dd4160ec3a6f325ac55f1c039014afe23a765cd4d7d2597770c669b0acd59fcf3e45d448745de186f66a0c3d49ec1e821d92a3ebbe60747b776f9e12eec7104f2ced0b081c891ae6ff0708b623733dba617edfdd616d00c3478e23f25d4ec8c87bb4d7190dcb6cd95156d28e4c6f530aeed588db6975987e81eb20a3e74f68d5e740240388e52f4b291241937fce8d0c894ddd07952e0b75d6ad4c4654f37d1e7e460d92ddce5352beaefefc3c47ec5b335589968b95995c36d149fed92547a4ed82f53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha840790010773b726439db71f14c733c286303d1c49b2f14f30f18eb5a36cd03cb1de2fc1c135f90fc4d29f899432c8d8ed5f51295c6a183c112325f57c25a564e38cb03a796d5f11d4a9b688ee96f111d0e7b6c7501de6f03810f037d8fcd5c6f3fc82f43a4f6a34584c8f0ea6d00784caccaad41c7cdadc38879fca8eb7cdc351199306ba2a61731475850103e343dc15cbf2266add4e173d956beaa036bd9fd654bd63764c5f8c075ff8eb3ffaf669303da7a2849d146db073e482b79944e61bfa644e5ef8da6a614f5cede08ec32fa90e014c46a96c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hbadaa94c2f28e0faba52e8a56168caf76f3c06e84623ec0f3a8a5400d8760c815f7067af1da019de3f67ff30acea88a5a89a924fd6f55dc312421e86d012903abc34ab022ae6d2d853870b9609f61b0be7ec21082f66b3a023a6449583c7bbcaf018fb0bcd7066ed566ed2a39cf25849089cd8fa13b1f8b0794a99390df78eb94c8c0973e6336eb0e8a4a9cc9de43e8b48d44aa2f2295bfde96df3bf474a8899342d5a5aa0d72cc2c37ad1f9f284a461b1c5d09b1acd720cc17b18f405a246d0c7c6726583c26759817e291f7be89f5bda91956f78c2eeed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h787675d0ba92c8f89eec3a3bd596ebb4f9616ddb9ce006f9433e39dcbd25f01e8980f1ef271fdf11a8f1eae4ec536d347cd4353ff9d19589fbdbdea91f011bb4ef12cf95a1aad7aee7a5ba8fba2428c8df701b3771c8516afcddcb79c77bea8eb055395a8fbf7efa438311901811d3095a3e2830cbcda9a0cb4475cd6c43261d17b78f59177b5e7e5895484ee79ca97405eaf41e5c95457b0196635effd59e4e526a5ca090c85957a036e2005e88039bab813899d5a8f9a08c65da62a16d05f4d5ca1b964d080b40b224e972f76c331102d54fae5beefefa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h4c73b3c68671603dc13f25a7f87d2e1e4e098d58229bbf176c53621f60b5ff04294f6fe58018adeeab50a4ee79adce0c0c67ca9175b816381f8f8051e15adc46dab5be067a02ce9c918782be7b7622ba027eddee8db4e298c38ad3fceda07585605a1ad3f808a9e559a90c4ac5dbf7be192d3dcbe4001b003d5fb6de19e17cca65b6ce00fcdf8fef49a6fea59f0694259b4232606e4f5a827f8d1c8efe5628d5716cc711490397dc042252997a7fb094b9bd15e79a70b1c098b2891ce508542c4a71c5b46820f57a61bcad38e126493cb73c6741767657fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2a2f5675cf94b38073d735eaceb56a82962dca532ea36982ac71de38c83c8fbb802a08d7f2b4d0dd01fc7d351f482ce891071b90beaa86b6f9638b8aa5db3f846ea52906c0e37e1dacc14a78670243847c8b90fda31ade51e2eeb4dbda67d7c45b7d79c76b1106a79d05eacd595274ddc2c7acc3bb0d0d40d8c7a7da4a09c2be8317f0aa5e9499ab779b76df7c6660735d0e7ad91b4e2b86078d29c3d45a154c6596c96153d8adbefdfad6c13d3024966b991ad0cabd334c655615f623f9b799856b6bc05373dd746dbee3ffc65d10e99a32ead014a922c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h30c6e3219936882d01bd18a1763e4c11036d187011c6e6df13271a7b68ebe3b70bb29bea04db6c72fe2cd1e097aecd29740c25010205b40ed361707e03b8ad6f226a48f4d283727ee602d1343f72fe8e258bd6e5320237444dec9aea00eb1797c7ee38639b2d4b1d99b2dfb33a849009009246d07b1316ca2be497bc3ef5091ac0621deb0502d6ba818f0068f33d4b6566f6de36731e9f8edd0f93218f5485530e7ae5ceb6e22e34f13c85edd0bb1b6d2ffe76cdf841650a79d8dd5af09c07a5b5b8ce0102bd56ad2e29933afc298cdea937ca99496c1d2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h95c81e226cecf2e92f8498ab50ad0239ed62f7ec70a8f04dfe19494260b51c06e5423fe93b9dec001c22f7e8c6d5a997a4f9d86cc4658eb00d3f783d1d77f069fa6913c0cec2913975037834940bb2b0fb2daf4567ed8ae7d7fb18d395fe39d9857540ed88d3464c6b8990819d5f69b44e91d0a8238cd67491b47fb1d45b7aa0439749fd089e12b492416d3972934232962fbe9f2fb4759965901b8c035a94a119c67d4cca3467ba71ce3aa27aba237adc8f99e83de8f6815f4385a65afa2fe875d5e1b40873562b7d4f96669c794b8769cd3bfa5759364c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'haf0287d32f67b16e06831ded6e65118336ec9e3705423c5de6a4387ef720f2c3144e86346fa129d72d86cdcb849a343470d4c0b24527b6c49430e04b63b75f217607da39bc836d476868d51bd27e34150e17f299d17756f28e4542e7398bb2264b437dd22b653b3f805bb5d5df7089c5c63cab7085419d26eaa5db4f5fc5d5bd6b32789b554789bef464bb0c604b073d563aa54c9fcb8b69c1d3e371d5a7d1b5658b76f84f924e435f1af1b296ad26866e7328cbf89018768560e34fbb2d39be91d802aa40bd7a7c45521baab0a1b1384fc311e72d851587;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h455396cdbd5d00d5c67cbb680b4591cb057426b29767d1b5c270b63d35b0b274f0dd422c61a4d497e7e10914a2ba28d3c4d0b4caf78d698b60e187d91bf21dd524d5fd183b2c0c0174c8f3d14609d5ab2f638a97f3e207321e683b307cb8ed9df86cfcfa624b349ae2f44878c3af3f4a3004bc466b7a8669bb1d01a1d5e0995514a6d0a16776cbaa78790a9e6a6d42ece77668b2d6ef3ae1376aeb1b09c1b4daaa047596334b209a3687cb1c87397a0cde62e4d773c11ab0769d620a0d37b4ff37f3743c7429fb6dfdc24d960bdd7ed75a129ae7a7e04491;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb159dff3b31b7f3decf648a4be6dd60f70c2105935666cf520deb7c0049aa1e9833ad6271abdaa48af36be5dd800deea6ba0a0784c8340e6df6ffe5dfbd7fdf9b92722775bb1294af23d36b6eb365b782adcc0f07267ed19b310c0383fd72d101b5fc4a2b58b88cc4e7be9ef5c3f376616b9839a99a3dbb358dce4ecf7644e681941ccca4abea57ed401601866009afca5b515fcb687ddaf14e0799601a54f15aa3e7874f01ce937f73c41c62b4ad5f02d1450b27f484a1be700f6e7ed278897e338bb1d696d0f371271fb3b0dc27bf8b5b9bcd778ed2d64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h24bc4b90d647000ac4f6834de6e29dd6e614d69559244ce4094901a737495740885bd2c631bd80463ff1e13c9f6c08a27fcf9a2ec424f75f4cd4270f05d00a54fe4d3a1d9f4eb9c04dc43d9490ae38c5962cd900b885a153ff8ad9a47b76b9a07f55348be37266d80769f0026f157f0f10f76c2f1243f6b19886346cfbb0a7515db95a6606ba801b2dc17965725c7c65fe82544616682226131cf1390ec8b9d496c086d9a255765c70ffa753df256be91cce20e06c267785cd7b3830052b798c6c5befdf21d96033bf62f4555cc44a6b2afcbccc2366801e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6063a166c41118a4afdd887c7a526dcd62c7848233d9f62b4cdc21610c4f6ed083f6413abcc665432ffed4f62c9676b1a69e942dc762d47f432f18e69e6c6265753cda055bb0804171d1fbe2599acd392350a8ce3d153437f5b0e581e8571ecc8605f884d0b487d27847d2342be56725442366e23c68a9cb11b70ada3ebcc19f496219bb39985aabe3abb25699fe013e126572838b96f55ff30f274825d8ecdcd6038ab5a882f711a974d79667261a3b8044f39ce081e56cd19b14749c85366c922cbc650ae868cd033509d558c2f6be66ae9be31ccf00c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8d75b67fd5bf2aed66a0f229b06ec70075d5abafe03607730c2ba340a7b5569ad05e70ddb2a1c4dba03cc51050dbcf0ed10a108b1ee528e05592e05ae3ae47d97a94e59c00b6a56df6eaca5989dc6ea56d64726917c75221f8d9aaefc512cf3bf746777f71afb79c3d3f35050c3f8e265249997ff9ad71c0da43921ab1440962f9fc294b41ca5aff1d2d741c4c48a4afbe40a240e6501891b4c596afff7109578c9fe4f2a828bd9359227471a8db71e69d83f699dceb7dbe74053d61bbbbd84a6cc9244f6ef5cf188b87a607d9a91ac087d9cb599447c200;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h42cfbda6e5a9209d982d46650c3c2526ed9a448b912e70b671e6ae95f02c9b0b44ccb0c3a54ae9d36983ea52a4595a1c38e93aeb4f9a55ea2fa75cb9d3de701635c1a8144ebd9f46db7e116fde390707c9e2119905227fda90898f6b5b49dee1eb1279a0bb3e4ecdda6afece7502fa7d8cb0603c0769e8af810c422fe1b4445ee2570b6ea0a69b1e507a07d12c0a97a2dedd698d60acf4bf0ddb1e016b0473b4a0345a4b4d13a0e5d3bbb153dd8b01286be49d4bb1ee0294f62152d5f42bc6e7ab5c16665860a08c25b5578e10d0c9a770068a95f68545ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf882b762b02ac565e7fdf42672354910f9fb47e0ac3743f9d339130a72d960966c4454f99c842ccb9482446d51b823b5daeaec1579fd61a42079418a9203e61e5a665630254d805cd8610c00bc84566ac7b98b28e46727e120fd8e979d225962a89c11746609de9abaa55ceece835353fabb7abf385a774be314b917fef921f55033e7bd987eaef67ee356dbc40e01bfd8bb2331a061b049244496b5c9a70b2c50a96d077560bc3647c28aa6ce3de842d53c66794e4b236888d82d94de82276ac53ee50e1e0071b8f946b3610d35530c34d20145c051a350;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h288452ee8373c1b28459cfbd8279dec87fc5d8e09cd7836927dc17005e0a09c5225acb4911c7f970fee61d8664ac5b1a530d13b5ab999a875b428b41b01f3467ea1f0d9557d5d9da5dcec8bc3f12ca7598e02db896b61ff313636ba97a806c8d071f34fec4b97b4842ec3867cd116b68a5b023bb58bdbc177f269b33e0b713f1fc778c701391a272c98c32e9f499bf4eaf8d0c4f541fbcc040b1e876be7cbc1623439bf3f04c46422c4b850fe99a86612970a87570e4800d9121d5668e2fc76f72406282561bfc40ae5c1a99c1e4a5d167aa00cc62efc7b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd26e4a08a71eade910a430fa6f4e05202bf6ea78c80967e653334796051ccc45c315864cbfb4bd47458dbdfac43207bfd315b4ab94848c873b2fdd2fc999bb3990617a6154bfb147f35ee40ae18523f52696ab37c7ef04a213b538196d0769e1402e2ac9645171b3f519ea6f2a972c7c62b548f0d63d36dfb643865520c42c956370fa0d7598d14964a3e0a8e522141501abb03eea4f85b52587cb0fdac7ba0cd6a187da3ec6a6b7cbfdd0f6888421336da1d780df537cb0109ddf30337177086b56ff12bb311cb1a0a878adcb700f8442779e1555104964;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3296c20d77217efc73225f005fe78080b08ceae7669ad892a78e75f2ce3b68231a05cd948426546bb7a4d0f86f46c620e4547c62825b660777ccbf6ac70b569ed79dd07e5e2c1fbd13451f4245fe6d8e648a88afa8eecb7ddba785275154b13ef0ee7f7747567ce8725f36937afbcace0835aa5703f02b823d4f7e1b7da68b1129836430b3caf8bae11670a7a45e45bfbcb90907e5764c6dd46e20ab303b7c701513bd3a3a7aad58f5736a68e71179e1c87adbe33dd71bece9603f5b6d3417349aaea6b0926bd77db0f567d12e0f821b344a4f252fee3c34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2ffc8cbf338aa7b13e57192ea78c56ec639c552e5e10392327362a4d9abaafd729a69af48f33282225b5f770c28eba0c963f7e84f18f33760884ed3288e175a1a5751f71c246bb9d12f595cbd49225ad18aee1fe995f94901ca9c6f5ac0166c0f96a51d91a0ecf3c0655b08f8505af4d780a5cb44183de93e052f192b288245cea61dd972a671aef53b53c4452ff4274407f613047586e9b80c440543564b9ad1d61883a492e60e08ed13b174ece285560b0bb68bf230504de5f3584faaebe2450f30bfe5f38ae68a9e856087fc9a625c29628bf009e37e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd26aaba22382f8cae08f9eb7579f93f36201c598dea0101cdd3af7a51009c994182db20a4a913b76e4276a901382bb9595186f4eee6c7d088371d5c2906b5eade9dfd9c3d745d1fa4f426123c4fdaf8b4fbe5728d25b16638136bac3a65a926ea2b1a340991d4ea23c646a183238f09d2361a3b33e08ebf7ad2b85f1b22152c342f460c0e20efbbfa128de1f2b508a70e9e1d020e25a03ef8768d23225bef7178378b6c7e9d11cc9d8383bf79d522018e4df4ff1f64e65a3f30a3fc4cb2c97812a8675a9d145e880f5c59a91e44e9f5b2b836cb4daa4d833;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd8eb43d92bb9aab5ce6ac5e51b63796d026a0170ce99d2ee40315804d1495ac5237b733a9796c2db56e63b58f12bee7cd4a886f1b4a01e9d7d527c431abee372028b046ce0685364f66f5f9e006d9710fbcb00739a3901324d2669624ed1c9c8a8d1d5a57578d1965ef705979e875c9a716ce19b87e410b3726490d4c0af604e494019fdd8b9ad463affa1aa4db6b99820201c55ec50445a3bd939067a8f428c3e55f14bc89616fcf540fe6d88529f11b1289b5381029e8a5de8605c3627721a9eb4e02a0413dd433f38c78b1562bb864a444c26f02fe7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h70a28d92cb3da184c6526c9dc093206256b08f82b90a33123eda30e268b15711c54d449627c7d4defd5706469243fb15cab73830acbe0aff92badff57dd3d644d408a01fb650c5296cd6c9181e47aa6bead0349d693da1b0ba543074d61d54676be8df7a7da036e35f555be6a20793e61ad198132d27c80f4dc66cee42919fa60a995e1a24e144254c28694b5a4668df2f75e71bc579af76ae990fe82974f6ce4d675cb87248e452b71ce3712a4cbfc88298b80d3dec88494272b58ff5b1a2e1f031635db1415938173c264d6fa36e6f4f8e1f53c4dbc098;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfb8416bdcdd66db223817fb996daa6428f1014b41017feb95d0e83ab7ca55252b17cc8e401777072450892214b12f54f2db65777c9632a91809212d4d060d600af503fc67e02586bc1831784e1515682b3bab4ece78b765094a64f55b5b67eda63b8ceaecde5491e4eb23899d5d85d986e5bbe36bdc070f1732fcb8d7e6a1c11d13bdf1afbb8c91566165d7ac5b61c2ec220e56f6dc84ac05c6770c7b28e466bf06be4b79cea98a881e9943e4d8df90375017cdbf929a5072aef225ab519a46ddac7e9fdd0a2edf0ae6e9e1f41ea2866fdd4f653b99ff9ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hef8b200ecb96a7c52655a8245aa82de4393b4e09c6bd790cb39964f062007a787b2566f706d22fba427367adaececfa387b9cf6ebe8b5e32eaf92690967bf0ba7b705c647ceae738b3f2ad2b04b9e753d91ecbe45951a3fb248268e66f6339f930c508c11876336146d0a8a12e952380dd6a1fc997607fd6b8953010dbc2a0a3e11a326da63beba3d84a500b72ef5c094959ead66d7429112315af433d470ca7015c309fa6d4ecd72096ae47a84c5aa5848b615d12f6e1b71f584167c74a2c44dfef2c2cf2fbb46295b63e7e8dd3c7b2db27ae09401e603a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h851fa5ef1c532cbe69fd49765b30a28a0c8fd0c4092c3c57a3a141f95d4776624ea8d8262da2848bddad37f8604eb4ed5d8dc0f062e8022f6a6f86ae508941b7cabfcd7803fb50e84b5ec7b3db986ae9a7df5d9f07f6a1b86308b5d05b976679c2e2797d6551830b8fad2f39b0da6f6ab58995039cc19b02914b4106b1ba347911e77fb5926f077e152f4f14ef8698f5a19b1365c69af39be265e7cda652a33e842696b728750ead17b4ce525995e15e2da8a0f29ea1af4d1c0902569549f54d8a595070ace27b9f600e38424d626f1b50aecb6ed3169739;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h592c3beef43474eda10df6ef8f493271ad94a6a0c491a2cedc3cc5c284fbc5abc0bd45c0a72cbf87c2d729875d53558e52b1810fa89ad4a42233894d5509f10c3feff14849ec421caa100f4f6dab5339bf49ef61d3d1d98ab17a8c7eb90db087b11e3bce6b9a536b69815c63e1d7ebdbac4049ce9eeb5f33c9e79ef29a15edf01a717d9b8bc29b4253646dbf6386eb04a1f456c99e3c593c2720707f49b89310ca34120f9d1ca4371682cca28936381acf7ede9935fd97d94e1b82d9ee9e30dd4bc2129afb42f0237640794ff707411e87ba308970ec16fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha5d83593c6f2bc6d7805aec1c90355a4510d1d3b2c52dacad17740b4ba1ff6b827781198b8612f76d0d216916d14f27aa92f37820387e81de0b49cc5d4b466fa6a3e20c692537fba87595841637225cb58736765eabaffa1add88c65fc6c02ac3223e13543425e33f1ceae0af4c8b02b86eb35da3e93383f7a951e4075b8a5079772b37a3671557cc53882c70d01268aaa419c40f8792f51c0c6fd191fc96bb2acf7096e5f23a8baa70d6496eabfca0b266b7033940d8cb0f24f35c0b87dafb0145ef73f17e8ed3cc1d22d7b257dca091d43f75354659d5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h94090b4eedfc9e312eed754fbae9847d1a03fbb68e0f7e7fc3bc903ff8aaab1e39239d082d4c7d9f6838893ac70e3ab5868b0a1afb256c068c722360a333ab59a49be6eddf6910adf3e968574cee4a51863a47087a4a4af391f785c9a3886ed6c47f8ac4772c218486f5e2d5219e0cb31354121ba487bc738833db48c1abf4c5161509ef2eee08eefb40891264b261ad5fc916b63493df11cfd577d0801a5658684b08be1f37604274153b7a10a2f879d203d0ad9f608814551aab9a3b865a611f304960c20c77a19becba278c25ea629c640223e0b48064;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3462150d7e6a44dcfbc491c3e257e48f5a422075147aafc8b0672d6b5b94730cca0ebf26596a988dbf47c4dc007dc2cbf9fdc8a22c165685f1ba815c038249ec6f9c8a7978b1395b4e04def6ace5d3e2c8a8a6d4ee7513f50d4dc47513894b8a68cbcb40b6365442b7badac761f6bfe59262bb768c95ab3e0b06f056767578f222dd8cad408dd53f47d6745f9ec19d47a589eabc78a987a904c2ac1de550fd8460e88475d6ef921940c546138bd95326ede844dc0b395cf07808bd2192dfcb62edd91bc8172ae7a3dea737b40edd586ac5370a346cc9d09e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb3a1e8832bdee826adc714f883e71a3c3719d346f51a39edd9a38bdfd2427c15ed289144003c1975d44fa17d5cdab3cb90447b45570cf0acd9da22cf5f95c297fb2073d00f141dc5cee2a2ba903016d8237d64455cbb06d286eeb2975630ff89d9012fef480b60d18262f17fe07eb93cc0e5ae474d64f7a6281cb4928e270dfcfe7a8d5a1d7a98c9a8995193fb451005ad1068867bcacbc4d34c4e66b4747879909c056eb1e3a4d8aa72b8e08c4cd0a02f83d1d32431da3c731595d796e2f14231bc18dc3dd109aeaf4353ff76653212e763f98a18b8a17b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h26a95149da4a7a85167c40eee0cbf8aab97e6082d5e0034bde66bf9fe3627938ab911f201bd5445762719715a40ab99d9e54481cae2e344c38b3bcdd467e2fee6369c09ac92084342b140d36ede25686ee7136d90b085626750c9c8388334338f82ad3cfe1a91448b3c7545214ebd20608b92d21155ae841288974e3390784b8e335889e8cc9345c19a5bcf899bcc8ebf3b9f54a70e004a7bce4953bbfa9bb07cd9294f53167550b1487e0baabe9ab0223e0dfa30e61576ae48f8c559c946980d98decb6ab5ae097f9f139b9e1316a11865dbdd1fe9f822;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9d214ed7aad37f536b46ee54996c3352719a34c1e813a3275cb3c4ce91e12a0ebf1f8066341c2505d7c7b770a98471e2dba6c1e5801d5941326e493af24916a68594642eab0885d71fd82e90eb2a377deacb79f7b43ee672a9ef8183590c594353549ec8a8111fe6928397d3c8ccc6239c22adbd7cb2301bfdd7dee93649691341c86a79e113a9c70f1ba692eefcdb48904cdb6b22b26fd54ad9a6dbbc32efd989fadf95101fae7fddf79f86677e86166645a208a21ffc34ebbf5ba5aff4bf23b9bf6a548d81aed51456889d4c55851314089abfa6784fec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf4130f53c4361a1d2caea60e0f1eb2fb7e2570449eef0b758c8d210732313569cb1412314d52daa7c3b19cf477fed8f207cb23e0f13aca91b7228d00470f10d5a891914c85dc8117e31d1ce1bda3bafe55e2af0f2f8e491d3ca893a5b2dffc91a3797216b23a492a9a0ce1c70f2bd61616a8f76a15f846680665d35cc418d2d5479909fca5fd0f18afc929d359ca1cef9276ed858fbe40b62b9a1638e994f1a363bc6cd680128b52981ccf270f0bd387b1a007be1accc27fb08bf5e81187b08a64f88373e02bb185b6c61d6575d02826652f60f4d689a61c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h86181f5c6085c61ab357f22527ea8fe43db4164a179574ab96fd49fd271f32990c48ba9dcccd9c08cccf17d4b14d23785d0d5d7c8679a693a6647399680cfdc509c8c316de75c77be7714fe43019ccf200950a545335a41c7af85a170f7e4f4d4ee7467ae38dc04f9545b4d9f9a5b6734357546f89ecbeb0f679e6fe83123160c80ac941ade49645bd0a2cb6d912c85c2ab34693c24a0daefe59fa29eb568eb813a80eb950fe72eb7871fad8f928b05d9020803d10b27dc64f67ef69e24b13e03e5a2c2575e21a02927f27b52021a240a802dfa14caec3c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h615b1b33cd95e894c62bc7169617ad498308e29156ac4daea8ec9ab781f4933cca8d23d9f859ac5e77e7dda0078db151e2807af4f79cfe442b25b84337237a5aa580492683a56e8ebb0cc1273cb501ef6303472c8c2fff93c3cd308cd4271db46c3d19787dfba8931fc42d9daace36cc27700b2cc2c322801a9792f39f6cec46eca3fe614080def7d613b5ed89b029aa2cb0fb12d0ae62318ae6ed98978ea18743fe84b685f99a810015675f75c2a02d02eb3605aa5c6ef31d6ef2e592ff0f8ec47e7806122d1f869a24a1a762c4ea03d4056f0b371a6b01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h933221000b7c6d45b70607d662fcd7e9f6e53d5f9dcbc5c663aca17458b25690885351513784f9726342ae21cdd50d621b6844514852652556fd939c6ee6011db6a27ee36096e40ec7f02832f75a432121362ee37e43109a830da99fcc983d3842b461776afe5681b33a7c1f3d6a2f1940c14afd2a057dd18422d7b4b5c30fc75f3a5482c474251cc45376c8bafce305dad7a108f62e563b7f7fdcff0b9cb15aff906913dc1ee1f0f855f9b521f8ecd35c95ac5b2170f68b6ab0a80c02f91ed6662fd8ba985b10768954b843282330ffa27631c9030ddc72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha57e3cad49a1928843159ae62b8f857757fd32ca9e8c4ec8197e3432e732b18daec21858153670e798fc34a5f438d33ce83c4775a0ef08f6805d7fddc37acd051a33810fc5f735359a6d69738e08fbee0c10ddf92eb8009b042082b4724f43707d3fad16308986ee0066e00a0b2b8d819542bdaf7909a7542895f1f6b17111857000d19292b4765cffc584efde0bb7bfc6a522cfec44ec2bdad043f41bf2514c3610cdf15104a0a90b7aca15328d4d60d54a54fe22d70831dbed863f09dcb98be607bbb00fa055e392c8ecae9eb1e06783d9182962f4c5d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h68ab58c2df3eda934e5bc53d2e8f47e962a2a30aab4145bbdee95c5bb576e295501dc4aeed7edd5be6b80e202b2ab15b1957aed84345155d418eda2517bf79627bf221fdbf88933797c46190bf4cc49e3f3ebb950093207870c60e58031ec62eecb59923b1ddb4c69d78d590bf493649b19c28e98d2bfe8754b68926ac68c86dc658d4599338da907e5619a25b43a91daa672bf095455cea4ab78e7a30892cae8522aa6ee4f7ca5a0b84d2aa25e28b7e13c82ae15543988935bb5a776a36e57c30297918d20a866fa449ec547323dd27f5bd8712239bfee0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hdb957354486bb8a2ee7580fc505cf79dfa216b7395e9200304441b0caad7676a580674fad7d5ef98a43026c83fad5dd1df0c15a3d6e9e285b866b793369b440c0ea5f83c0f7923d9b509ee910b46646b47b0f6a691d0aaa5a660841cdcf7a1a66c3131ee7ebd01e7c9f8112a9317f1debc41959f264ff45c19de0f3b2fee026ea573773f5192d004508c673ef0a9a9f9bdaefaa09b0083986448a32e11ec1159298b193ab98972e43f10640d847b76f669442f1ec27cbad8940159e30d1e34441812de7ae5abaf5bd2047737ab02e15b75084f3997509cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h723755520107f6ac7f31ddaee715db79dd536b312a0a2cb644a6b295fb228cf606c52a224e572d9cf2f9b49a233d9e7c80b3371f0754a517189af7719311f5a77f7979c84f601e5d9b490e11d9f9b0389299bcb4be95d429cee0c311864e4ad086d2961b178a940a137a2f3fb77f9ebd29013952ba1603514abfa7ff9684065ed477875ed8bb5229524f7d700ebf1484a2a2336e36057dc436a0ffc3e2843ef227c18172c61fd31c7b8929eff6976d485c5bc169f5c8a84aec692a7695a567b375fd5c513e88a23eb51b9542de19cee1e4e8479321bc37f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd50703989e3bf3b866426e9c2bbd3d93ab7219e38be9537e9b75a205b1c1ac78dec0b101b6883c2aa6fc69ea032df3d2d67a8bebffcdd3e6f2af3d9747f9a8767485be451b72520adc18278d282addc53fb4c644e124ff2d4866ebeed0b791f77a5aaae0e5ecde1b9918817ebf0a3ffa3a6d8faa717e2e18144bfe87b036702e49df772060a27a2f7f462a6c3db17151c2c9e61a3359c5f2629d626b8c897d0b8d08b9777ecce55b52dae8a19f5a755efffd3e9a4834b9d54f5d28b285aa1c46e4df9edf1328067335c61ca05b15ad836f4c27313b11f4f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7db1f39f8fda4f629980bc5841a8f79351c4a5b5c16421b942cf18e42d265d4e24488da0088f4d7b3eac118dff4e684663bff9931ce06c9eb9194e0dab4c1e4b54438a97f26ce9211292be976d2edca649a13be0d60f02b543d9e591264fafbc7ddc583e5d2db4f282ab659a04efbca1bcd52a71c4a46f41b3947f212276f54775d3acad6bf9da39062ce5e9bcfe0ed26d5fca7bed992cc1afb2fe06ad62a19ef22928fae9e25445b261738ae3e5a1f5d79473cb953988f73e5db9233631610e326f0c1af2463905a8c85c017db372d38ea0a47b47dcfc7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he18190cbe957c3c7f641e7868f6c051812097f1aba2aca3f91aad1941a0d27357467c9285dd590ea58e3ae55375bd9c86179f7ac40d03ba55863afafe371a0b75d54d2eb6dd45367b77f89b23e1cdcaa8ea8e34e54c45d3992b79d8ae8768e8ff24e1e43493f080f8e75b3026530f93aa418811b6ecd11e1dabf5605956d4474ec56770f51c26ab78aaebf37a17ed96343bc466a872e421f79f0fb40f07c5cfc1c039d8671c5384d04d5ae35abd41d691c59db5324c89b514f3f9a8735f10e7c2c4c91b965e6d8bc9c66c51bc776e71880675ef79fc071ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'haf0f598407bffd931edc6e7358218f717737918781fd13452b1677aebe92f435bebad41f73bd266e3d99e261f7888903002f042d2d82fe92313483e3492622ccbbf831a486f022d1ce61d2272265b2a34cb8983d389f4647c2b36b226b679e00166ebea8dbad2edee653318a51688ee066c7818bf5e4e186a07d7b51ab53572cc6a1b69041bb95b08cd9d795f330bb37fdc17b44a905df29f7c0ba2c0d8cb682cc87ce8e0f4306131db61a7f522d8d8d64d52c9c5f7f10f86fa61ac4648f279289ccab96322ab15ce4563e30cbebb7e90facc1fb68255a60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb825844124bcc8286b5fd4923b5335c834053a934ff1ed0dfd64994f21ae1a59baeff0a668ce6a6d1b0403478fb6202faa111d1552da40815d6d06de57816a843901e028d6271245312c60a1e6fef3b255e648ff833a195ec4fc7bf8a694b5fcd73da33e84702ba2b8288143c6dc8ac1610369e1abbbf81b490db262e95eda4195a48751e036ebf4765f0f7d014a2bc48b9e56902bedd53a96a16750bd14f4696ac754df4a97a05b5d5eac1cb43f5e9e46ed811a211c3c100f152a1ab4171386493166f7224168ca57df17bbc40c59ad983e150ddef803d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he6218e7fd6afc5d6ddbd08bf1948f97f52f6e1a26af9e2993eb01521448563b36e9a3e1056b417316e821c04b60857eab53f88f3a78ec55b2a0753a21c2fb832e969c0198fd66a5582fe9688dd453bf4cad6c8cfbd24cc5dd22a7b5ce7a2668bd7cc14002a5c281536fa1e52a2f6419c2159fdb340702bae8deadb294716bd64d7ac758c6d236b45e0ced4eee571a63aae6420e58540d1c9024a2c2cdbcdacd48efe667687e1fa4c5f0126cb7805619a287785ab96249c12520caa4d00798ead5982dfe4c0dd61f51558e588ed7af78b68ada82d0c17be3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8a3d5a4237bac8cbc1274a0698ec7dee57f309bc83be5a7289254d7baec00c943432b222266f8816390a20905d266a3149e808e8092fcfa6da3a606fa401c7407ea547f5653ad0a98e4e872ec185fbbc45e1699000ce673b1952a9ed3668b468004683aed8fa26dd4a6f094c9f80fbeb1aa21c61b5ddf63fe3d62d44aaa5791d81881a5bfc653b2b5f63080551e5cbe925c0f9241bfefbd59f330087096273a672a4b03dc065e93726b9319c938aac365740d674cf1f5cdcc325a80e2bae210bfeb6074a3c9f8484b88ee2bfa7608a8c3fd17cef3ea22d6a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf78c45fb4fc2b97c72b7e7187a06a002afbe83032352fcf6bbc33f044671c084548ed9bdb9e839a40541b4238f86cada0fbfbdac897e29ad2861673dcff64bea42c2c3780a2ce24f1288cb39f81e65ce195f1047b7bc847ab9f6f7f67743d319007507df24be735fc2cda50ac5f941b7c3915bda5e084dca3c1a99c66f9a37c2953d71480f91406949edca30675af1043991abf9121490ae8d78c059902bca752bd158465be6aea16dd4c7342b8d39765ebf80296384deca1ef773073c6075680ea15be0fd1f981d2134e066d4fc3aacfb2119ecd5e8d925;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h10359fd2e1041b9277430a0cb4e5a4cd437135df0e1d466d0985bae0e4c29127a7dbfb4e96d9cb0bc988edf4706dd9a5c092142726a5eae50283868d9d4dcb9d95913213e285c74d11574c67bec040d05ae823aeb9ec257df826ca1e3c0390448eead2d77b141243cbbfdbb4431bf98ea4414a043ad5499fc985438f431404150390baea146b6d512c859b821d31182d6418c0a13701a254dc45c8d3ac9f743af5560878ef1db5b2426a0a66de9236907e67a28af1fa464288b6262ba10db016958bd4478c66178b42c6798ebb03ff2f4dca85ef8fb4982e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he49781e57abe13dfaf380e3ee2c3b2f3b4f73fa76389f1193086119a26b6ea5259000ca66082fbfcbfb15a02b0e20f5c07896fbdb536d2ab68b3f379951d6ac0b7c3407fbf12250d5146be91754833a5fc3eaf498c938cda6dbb71590745a9dc9757d7af36b62681fb2681c619dc004ee3911da90edcde2581155d3634a9a9b9ff567d626a03a5eb043af35f71860cc22862fcced50266ccefcb27c8ea737945c98463fd0ae70f1fa2327cd6f9b14606f934ef8622a0f5e2931a3942bcb752b66e8f95ad8197c465209af3a794778c2b30c8597cd04a0c92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2a0ff3cd4faced2b8a5754573f947e5757eef65ad909aa9d2eebb3df3e621a9ac4ebdb4103c29ee1d8a35a3ac1d8aefc39f49a07ccb0790be99a7f031a558a3f87df82dbade2428ed8ff86feb154901a79e6a3c22b1e98178f0e2b71fe1aeea8d033c0003973e8f8b94c31d7bbc36874384e6f7a7810f6276cb967cb910677bef68b08813e8aef7dbc43973aadfc08bb4b026e617c8b6b1f62652bdbebc3c1f57b350ebcdaffb8b3583270753731aef4816fe5d159608551bb49249fb2e15b1c1ce8a91f9dbbc319bcd4883323e105a5d75048c4b1c9e583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha9ebe720b1580b1642163c8e9431b7a91fb5f2c28f9e17665d7bb0f9c28d6d08d7a168d2d6557039424caafce7270f5ff6f7394c616aadf9c1c1228e9656407fb219d4b3f279d66aacaa659d81d9bcd9eb7a062b121bebf1deca0fce1d4069e95139c9685cb0af2884728214fcd7112a7e77fcb05d741883dddcd364d0b8a5d2fb63f79560fd6b72abd068950438d2ab1488d6173c6958ea23cde58e0bf2f49064a7a72d6f198a870517e5dfd376161301cee1c5c7efcea753badd692938ffecae7fcc96611c0b61f311bae72131e7c8c038c2b5dd508b3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha96a5f1d41cdac148f7cd9d0e25e1b52fea00135d8af6518242c21e18039a4b0ddebab02857876cf2dfce4479cfe9ea33402e026983f4da82b70b06027f42f56024451838f648969f9774a7c28d385085b098248ea3a229c7704af9153531acf140ab34d02e03f0f0a51265032663d7f6c1bf7712237d4f2dbf0f727ae944e6820ab9634d517bb53c7ab270d8d8c5724223d039b89a98a7aaec279bb044c622e1d5ec68ecfc9f704b5e91645b0f0ccd402332840b2e4c44e581a247a106841ac3fbe76d9538bc65255c342234811cc7d2b77a5cee1928290;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8557bcb3c268dddaf4dd86941fc70dfc817480cad02ac400efa78b345285a3e4d6cd4b2fb214339933aa2354b08ef709c249beabd4f72fa71a555a118166d76eee6037590fc63bb0dd84942ae6cde44b54cc9118ada83b7225726ba777c51136738f8f320551389f54255a75157039da79f3e6b0c6b14e5a90fd41842dbd37a693ff1312ee286f26b543aead64ae677e461d417ec08f04c929d1081f0a32cc0f72b53fb888ac61cb17f3a7a892f1cbf89700b3f7dbebccca0d851087ce46c70dc02ad361f0bb6506478dbe1d91f114ddee16d2398609fef3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hebf6fbf9abf392d6d4023b8399b13a558573af5acf3eb2009f7129452ae16e99dee0425da377cfd12838257ae2ac13fb2d4a2a43f7b0a83689f553b345e47b1cf2e7af687979706f6fcbb7066a13e9471fe11929534aa2ca6613d512164909592c7aad76d3ea5185aa0b54d3f15e013ac59e16339081e9304e0e2e589d41b5508cbc0cfaaacd2ab5fc20086518e5a698ed10c8f0344f21e51cf882e92b5f768b54a66ab6a3e621f00346d2914815fef7a70dc567887d355f6d3b3b3b7bf7a323a6f422b287b0b75b1bd0eb5c488860ad549988b4e62cad2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h291df00beeb75ef46087648e2df0bd40a0fe8e03bde390ae9a5d1c43175461148ab2b1d6a8656be6953b95c58e7381b8428e2c39fcc25b9b30af0159fe1e9dc914774b2dd1a3d3a39f9abaa355c8bc6903ff7fa4158f3056e6380bd79289de41c0f4aa85f4d1570bc4952c97dbf8944aaf47df2f88ba088d95b74b251b016ccc57b14af29bef6a6ff63067769fe2b3e0a07a005b16e9a2dceb1f82d1d714c8003471b5e772c3b13b0150fc8ba9f589887b43b03455a137fb89a6f622f2f26615ddcdf694a14dd9762cec25f05f21c929f479b3f502b93ec9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1e5aa552783cdd2e52134498326a756e1ffcb8c4ebdbc81635ff94bdc6db1cd43645c65e728b749b3615c6dfee6c0232d35a4ce32bafcba82aa17aaffe238acb106f413c648c2a117f5df6f4d721e37299d2a89592ea70c8ea03d6fea299937aeb7cd516143b2219c5ff1feeecb918bd986291ba344aafa695f85a64f760b0493a62d2063cd1d41ce120aec740907eed3caa223cf15674e0b884ea6dfa01a5e77dfc78b8ea6358cc3566ba29e71900a726c97b270df794bd668a6bb289212edbe4e74cef8da8261349e95dd4ca7bf76613f978efc428def;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h98276b8cf8d973e09363fbd84d21dbe04088bef7c176230575b29c2da0ca058633739a2fdd36b4269f0451a4ab4fe2f6b0c6c185d75347123475967a1a652a151f802378665694ddd1cf0f6ef4f40a7a17c23bebf3bcf02c92f6b8630a2f2a6ea2d78df22fe1bc335985dfe3f0f037334f19df057b4a1948bc65f78b4aa1a3223554c74682942a8ab093554f75083e4784fdd664b96eba91afa173c8fff0946875c621bf4a04f5574bec8aaa6589c4f11fe6ea3e0a9d8381c8ec189cbeaf0e409b7e01b5fe61512c41cea7032d148ff33193976fd1fb89ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9515cd3e4c72b16a256e48bf20a87138bd56a0d65b2b55dba6734c133ba0b685bdd4c4aaa798e3d5b9d17b39b2ae2902fc0b22e247e7c0ea088a743988a255663f178b0b0fda34ffafc8a0b6969d71c2740c33624f64be82a81cf82e9369c7e372c8567cab785e75e78896a4c728b3269b15296569c0d398bca91db88cf287f5cbdbd73d4f587d95ec78a3aad58c555fdeece5c5b58579e50ff87a9dfa93460122db4b74245efba4e8db7a11e9c5bbd0b7f118c4a1fe9f0b39f66daf4e178d7eed9f8932ae78d23120f5e790aea025d5eb7ee5b46e64a4a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8fead53956855c58835e94f79e6c6765c44284f759fc6691facac204f08037b473b3545b0e40e519a3c5650ec3425587f85b69d56df08d2ce738fa28ae2ec0f01e7fabedca75b9cedfa5441d07ba50b5cb6c5aabf0451df75fc00695cb18c13c4dd24335b895638e908c141bd87c1499ff1a2635cb7fc166d040a49d7d6b3b2a1828681a569434a126779ecbe58abaf0511f53048218e0ccfcdd68f1262a1325008b8d00e3aeacf1dfde9bb077faa9f1e171ae9557644824b65525aba2001b39f6622b53f1d2b377bef47a48ccc8201943fb781ea70a2f54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6a95b1e08bf8646752a3513e2199285aecbc8d61ca7aed42f6cfbce61d60e18e5d591d3a54e197e2f909627fff68825d3f6d3c7cf232cc9092ad9b748eb43ef4e5a5c12da3e56d89b7fb8ea8866dbfd5f0a5b69dc83610e376f35b21dc9fb8aa5b02afa47d729b52f935e658435a2a45272ab05508ee66456822dafd75c298d7b5ee658a92a4fb4b4a6d8cbc4108689f2482d4d7c026d6deb1a8179ebbf6c1973cdb64708455b2ccb2c7a6a7aa5594bc264fa6ab801c5217529cbaa3e0ec51b18b591d84b4579e0375b99128b62c4a0485cc5b0a57adc36c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcf71970ea8e65cfbb99ccef10af686c78fb45573c92a49c93883a62d6400c574bc9753e02955534ff82edc2d346029385df2f3d0ac6e0c5df8ab96cd6bcde06d23cc4b9f9f0f828d4fcad2abf4b57f72681e708d55f958a086bc5e2129b6417330faa7ca9dae54db917666e3043ac450014da9c1da7607f0b8e94c90d7bef3669c0fc1a4ac03bbbafc448df5304cfd16f4f246590e9dbb197633406d29eb3a070d3987ad3330b07c1b2816256d1f83f314836a42f86d8209faee3a9bb6158a3ce0255a2bf8bc031e7f4540d52cf782a49a244a55b39414ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3c43f546ffad9ebb2ac1f4d44af0b2ab99c4501c317ca3665b7bfdf58925a1a7209c330372e9c8eb1a7fc59b3421c78bde443a679ab0b43402d8a3b52061a0dc65830710bb3d23dd648c174c98c754a16712c13cf585ffa5fabeaaefd07f03f1003100991683f31aa0370f726e00bf5098047f0c50f600a7ce1958f6a0adad7d7c6f808cdd7fbff630dfdd0775bc068f6e355dbf5965800efb5c5f6211b3c8b613a6ee34fb1c8ac2b5eee14f8037d1681229946cef7154984575efac1d65ae49ec4dbf956f17413d5224a17df60ee2bd5815daa9fefb9bd4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he7a127218602114274e0d4c42c5f1a2077a28e42ef86ff09e9d520f684d5c8aff8ea101c32f2472276766d02d6ebc006285280204d85fb4f713581b05d5c3fe235ddf8e7e5146b5c763c999976a2ee198bee84c5652f7bf423fec3667ebbf96817a679845a8f64d29ea6211a9bb1e66d131d0a4fc93154f67e57104dea27344da55cb73faff7cf39393502cb4d4effcbc570d467fda9698e18eaf8761a6217fb1ad4530cf17581d75b5979f61eaabe5f82d64bd5891222e33df639df5575aa52bf71ee9fb7233c954b1dcec84449ad575f207ab0905e18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3c3c09e40dcb0b6b1dc9f283bfbf2876985822629a898df84744244c4d6a937dba3c11d5f899fb44124f2548d06bc8c0b0ab358ae9dd99f151385dbc2c9dc0475a97608228e5d7f29e0110173949686b83f9c7001e42e32a9fa4614aebe7d709f7c04ee1fb35966ee6f971e76e0e24a598ce260e22a54e0e7c3715546f703554ff893d7e0f4f8ad4585a6063ba56e0c2f34d2456b829bf70a837e68093922ce00572ea839155742907b3dae20d75cd7c055a4f65d8be70df07cdc1ce448b3c0a268ee7e5a951aa66ff83533febe87404383c12b634ef5016;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3b459c8ce6128b849549d93bc12c1a3c63d8a387a41bf4c436d9874e437f8880642ba5d282c40e0207c18992c7305f768979cc81b1bcafe6de181303fcf5faff44366d817cb7efb8ff53cf463e43584a6d0765f2e76db1088fce6c3179223bb527263e355a63f2c8d850b0d0e0529a9a3fd99d89841132aa132b5c710cd090894f6b7df3469a9a2e31dce14b08093db402967eab4611ab230ee3cc4782a0dda0ec83811c99101444ab7f50a8a3df11c1c554b99fe51b3c7c68fb5935211bb6e79cce781b39f2f1ecf098a93eb96330f5ebe7fdc054ce5294;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h803c1f21fe4934c0f69ca10220e72e2f800f4a1264f93a804d9fbb1693e69d09fef32eed25dbc188c05351982589b0df0e316f177d01177784fcdfc166291c2eaad089b3899b85293400935ecbf3b0b967750cf6e1f0a7ee82729acbaae4b60ae20bf2ea6fc75982ea21c0e66abf2c52260bfaa8075d93c99dbfef474643e09f01b2938ad64106e18e3e12be6acf861f3b120bc0f9537efaa1e52a49f6cd095d50fa0ab76b3eda969fc2930bd02c0d29cb8607c855815c343fe5c788d6473ea6735502e4984549f6b0e4858d2ae4f5132f0d80bc44649d4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3beaef3151e78b1b49d32da6727c083912cb93f38f0bdab6377bb170e411e712f0e556dd39b6632650e5d689d0bb54322bb218efbedee740fe3f9a8cf0265299abc2199de018a3f56b4095c8d601d9f0ff4cdc7de5bba69f321d2069c4ebc562e926d49cd79f6bb219c7bb13fa815c4b1d98d5d312c02793d9078a1f2f52144b49c5d0a29691867df11f2edbb9beea98c9ad332fc4b6cdeb3507a27a00a88e5c79e38d71972b384e25a442a261099162354a5b1b0c7c2307cac0e16d750310ded56e2a0c53933d667a8664dc0debd28e2d908841e6839388;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h60a2025bc675506d7a14aee5ef442c0c535b3093bacc8d318d85364b586ea4214291f17e89c7a7c53fd967cafd17124f2587dd9b3f54ee1229b038624b74adf36d89e43bb52046e941047bde8a05428287cfea8a7fd7b66a6fe44730acd7b5aad4fe5fa6e3772bfbb075a0ddcdf24bb70f4b80c1b10dc4d5f4650698df33569b635525dbdf4891fa5168070a5b8212c9a824c1fdba409e7d87b2fe4ba5b17d14769982c0a62032169e9cc47142add048ff650a18b6c6d2f2b7a760b0d1245feefd38dec31dab48a5320f99be6126f56d2d84b4d714280914;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5088230dbb7e47950eed676f5467a2c72c8940f3818213981bbb2f7877290102f7a86bc7e015dbe1bc2b9ad93cbcc22bf92029475c7f1febb6ef820f8028a946cfd2fea589372250445667dbb57f2d3f5e9b22f7aa1fcc96e66a512c2aae46993daa8da413d1a28622e284b1f489b36191695a62138f68f97024afb2e90990b403d98836cd3af529263a713dbe733066136407c737a2b7c60a66f078d17e079d7726ee7f398362eea94d08ae996326096133514457330994f728f90ffec95cbe685240ad817ba70fd783399cd070563ecbc40aa9f902daac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc77c33001228b103fb54354eaf1d39ded721d7fca686741c65676219ab2dbca9d01728f792326726a28147ac26a6b3af61fd81dba0b61a54f013e9e823c201dab732e20ad05d28997398a97d9d1b9bfec52fe99f98651f61d4b9135adb8f93bd44bd5b02a0ed3bf343fe128ae05ee4966a0b1f303c350c10ad43b002aee74a039fc8a708e5f92c61067c93c704a5f5b809efb62bf734703120905d398aa782859e70ed8e7dd8ca5244266cef4b96e25f3ba7b6ceed57261426bf19b6d76930f24450319e51aefbe9692b36ac231576aa14e407d1aee44f9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hed1e9649c6384ad58818ec4910ba86202d3429695a1333fd65ffe946e65d2fa68135f4e10f564a937b8eb8d9e1460bf7c210eb046dd86842a1432ae0ad34b76fcde302874f8a05d32bfa3ebbfa27fd28d8e846ebd1758f1054a8b27c5a751841cbe618bd390d6dcaaf8588bb8cc7bc57d0aa3332bf679f74c8683129d0e760027eea85c97fcbdf42be331ad3db79d2817b87f947fefaf611cf67959a81b67e0977ed5ea7c37525e1626cc93519e2bf7065f9d8fc4d0f4699192411cec0ad88a7541cef1145046c8c67052797c7593672d5f1305c62b3fe9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf5082c0515a1ee106bc93508798443f48fa8322cd603dfbea6ef5c15eab1c43946250310b7783aa01506fe4c32afcf5e6d6939a96d45d98d6670060a322b065760a91758c54de0947c4852b14fbe9480d42b11bb96312107105ff40084bdcc0e7c0e09a67f921309a42d1b153bc681c486fd1dd2081ed8f2dbcd5a853003c6db13e5d2480433dc09543e36a0e75dfd3f1ec1de50f7bec934b2321a155f3a5bdc28571bcd2a93eed21250b3add1c8ef0d661d7d5e5ce4611674d35457b58cba86432af6f872569c73aaef385e3de95a1b688dff902fb1c99b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hed37c654c68c1c4bf09f330ea0c295ccbad242b6b237351b21d67dca533091300a228e64da9190630f94b6388b70162e584d8f9aa76d4765571031afec134ebf10109022ef0452dff44de05c00b57dd04cbb27467759ae49835753e4a5e3aaccf53457fafcdcb05f131ec2a6f093dece01b72d6292bf1e00d9496daba201ea58f1fe7013162f81a960f501d0912c9b2fdfdf77aef7dfda709e8e80a52709d2fa80a5f40edfab4090ef57476c0a9ef83aac138bd42b6813819d0ce982e68191a44577ba134fad76c3c588dc1f8e4500684e4fecd07a8b4eae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hba842be4c7d243b252bbb0d369d69492a935e8fe0837fadeb243ee4f27e24c8a1bae91d5eaed963587079a5198d1e6430e619730065acb4acf06a1b0fe393b984fe21e058b9309981008a0fbf7c854788c91db28bce3f17974114371171b01c878136c5af754bcf7f1018d4d2cee1f7b35b007bee2e222272b751a9e8e58654e14f23d2ed3608c596341ddc63c46ffeb6b9738ea14672c8447a18da488faf32412417891dc6af5f1cfd1f102bc18eb820191ce36134046e7cc3164bf780a9c9ec0c09479bc3f38ffaa717cdd13f43e60fd153dcb72739654;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h76a1a74575b3df9f0a121be6be0a6eb6a94316f74083874249d784657f12cd9954c5bf7edae4e30ae85ab65eb3221249487eaca8b6e73c469985303d9d3b6ac165e4e07a4b6e99859dd6274646bfa2f30785e5cf4e698e7e8ab3580322bd3dffc8fad6418b58e64a531ea86aba9e544139f0c7a2e1326b8c2760d7b4b2b987bd28f424d1cac39ad5eb655ca31606058b0a3ae9f376b524667d290a56769e6e64e9ad94762fa19878238de16ec27b719f8097edcfd6833d5449797ea7adaad885a3d65de301d07ff276dd1819b9cb0dcd8152713ff7bcd54a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb2f70bd90b0c30ef59ee898689bce6f8d15f4ec3b4a136093e09082adff2a3bce1b29a5834ff864787372f055c0e91b6a51813fe6523f22653a90f0659c543ddc159bed2fa0927a347c8c6db31796c5d0d358b5d4e437987f5c6c6b17923fc67b7151d56e6c0a2cbcdafed23e4775a9833154fa8b6a9649b1cce59281c082d3eaa7b395ac9a37c14f0328cfc9e43b3ae04ae9c7edbd2ffe0ee5e843e4d9cbd4cd7f84d96f4dd384ae0e041998953cb8ff14c73f7dd5d93a08639c1f82e58b8baf2610ec7b89da2c242b030bd6354db8caf9dd959e24f61f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h24f46425bd5f8a02ce261950584ebf26a732b0e1f6aa8bb965aa232f6b9523461cdeb8f3deb8b91d31621199fa1745cbc7087f747fa7eb3a9a12aa948764148d04cdd3258d7447693c25ca5362c9fda8824acd8dc5285329be5818f63948d3f61157aa0c93a5b567ba1c8e6fba2e187b1ae4af464ca12cf652b38704c962624e40890a6e7d78407a0a94f0320461c84e521e5827142f38cbf47f4be06a41048f7dca0584bc3627b5bc2245d73aacf503729539b6e4bfb9fb82e20eb2fb9cf2a7035826fff1f0ccdb3ec4ba020c3b1bab1fbad9c0ab9c456a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h39826a0082cc22ee64d70e68b70dcf1c1c85d56e9cad1f662d63f05bb4b6136acdf84875772d54614b85b1fb31f4b9cd071a454eaf54f6f0cd073bdaa14d7f3ebbc131752c2e5f40b981381d2b29928977d9eed82ee777da0dac0b935a8be7f3bc5e4aa5dd661fa97ff64e0252c172375d81d23658b637baa6dd42bd0baed6a6a4c332d92d08b833189df8d76f48420a7504ec6291346dcfea79d6667b72555339f65d7f051b99a295f169dd6671ec15b3dea775c5142e7c4dc20da81ac4ab3d2f1d6bbd9471d78256904720ecbfee5a6f4f8b992ee47dca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1ab0674106b8136c40c6386ed23c243783ff2fc555ea98f2e1386393f0a271e9e2f345793450668ed12287a60c46fe07e64c0bf416a9ef7dfacfbb0252badbb9cb1665e86b487453fa6941d1ac80ff6e9adecbb90729499e53d66f7ad10f0c6755cd5fc942920334ed5fa0354b4142963cb067c581824aacbcd583fa80f2cffc315e126b85671f97e89fe49efcbb0f0b399ea83559b8ebe089905699bc2183c31acf2d3e088173b5566bf002e60b6c3043c8991476a170d4d18fb4828a0618181c1258a9a135998e0429f2bf48114ed2e3385b331c363d90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf49d4ab827cf373bf85498e9de2e20639b10cff08f44eee012735ce0e84f6b5bee42624bf1a521168cda76eb8db3eeb9ac2376f3d84acc6152976e4f58ea7d5a540abae4d9b8dccad020c0089b805786a94216cf07f25147b01c58d05fc128a4b6c7a15ce61bb5c118517fd04771ef90840d0f4cc119cde1a17f77fb2d4b5f1c757998213d1f0dbfec5a4620731e5635db77355379a8a1b5f6cbd3929b37e713b7fd170897eb35525c140ee96a4d0d766621eb9a0438a056569db8899e55d755f53b3cd30628bf222ba0da831bfb3dd5c8aabea3f8c86680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h521ea8e35e17b3cd12d44857fe265ae823a9b0d7ff9305fe8b727475ab5a4d9965e238e15effb3301dcad01db7819ba988d142da01ce300cc7d8876286f81e0a5feac079099d85fea910bf41ac1c37ebfbc8b4b9e11e194b53544bfd02da8e4e34856f420ecf55bee2fda3c2b5af3b38c3525c30bed5a34ec620a26bd95237b8d76669ed769acc8d246d711dfe1e0b78add3c7111de26540457e127cdda0662f7746a23bca8b516f168c78675d857e53d9d92b75a617c699822bd1e1cf93d0423a197254c794917511fc89148cbb110866bf94992e7044ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcfc19bd9961a14126ccca18e838f44daf39fe7d2fbab5ae86bbd707cac4579d876a0a1c7103014976a7e067dfc52b43130be5d172b48ae346c3127306c74b01369ee386c5e171ab5ca5214d5afd4601c472e5597bcc8222e2508178ad3c64e108d1edc522bdcd65f9b5b3485a262cbf9963e9a9a77edde72cc6e18807e4eb7309cb7b47dc939f03fac8a54187e67f8910d73f14d7a5a5118fabc6d739dffdd126fb007c0a5397fe522368d8af4a62dbc8467b92ab4b42c43041e177723ab064a147b8992b0debd2598f95a4ad50989cf0dc688a776f72a8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h16584bcc0c0f9dcec71ec7d8762459fa3daa9eff90e34eade0a782236b93ae7b25c4f2a0c8a70c1bf416824edef2f926da211b1bdd6fa5daade703f28cff286a5bbbdb57a2aa78e152a5f3280142ec7bbff8e66c57797c432b5e54cb242cef038e86836300fd043dc644bedaf7f4d163d6ae37fe654403f9da1443363f51b58d796fe0fb6963920e0dcfcff678927757d629b02b13ceba0327e646ac1d58b1381a418bd50e4430df7fbba88717d4eb4399eb7b9944e473c4b973d0ec61326c12d3b58b7b91bcd07106bc2417caa6405164b298b03c9dbff8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5812ffc59eb95c74a3270ec6fb071898b4361e89292e44aa40568f946e8a69292c92e719b71394fc0f63e08d9307af47d6dd875de8be3c835aa468a56486be1a270dfd32d769aae97d642e63117ac88b1e5271b7395b02992832ba266d633d42b49dcea78a5ea536447c4e44b7665c671bf4a42ab33b7eae2c507e7caf26476657952af12533833bd1b3a11ee83c479c83e7df64df757063096a5af162cc7844b8b7768939f6814d86595fd841d50bec530e78c09cd3200d3b76db147bf2e2a21435ce675e268b4f59746afbe966c81c7de4b1d7ef07d00d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h72ef7860dbff17532cdf5c0c0bd83e9e373875f7265d1bf18f3dd0d9babd6e5032f32c484f5377ed035e4a80e71cc5c851e596465fa5011a19adab739d20bd98f00733251cbb5c4558765230a0fc4e95b243d667e2f0a62c6fe1664e5b7f580cc9efdfd60f009e72ceb8ce898aa366fe2e07cfbf19f379d00f06c8eb4ba0ea85ad55353fdaf6b5a2eb161d555641d4124f4cdf9c8369b73fc34ca636ae22f5654536d73d6314b60faf6a5fd2abc0d6c774c4bd19dbc07508732a671a6dccd7009ec97ffed9a9240e5792a4b54148c54b8551621a3bf29422;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8e7bcc6673fde0d27161a0041f8d318d7003d80a5bb6b8efe0ffadeabfe00e2f96ed39aac950ffc2be626beff1d46f2958c6e4a142e4ac349bc2ad51c30aa96454311e9b72b765d973bd2336d7f3b399efe070de9ef35cb5038bb7fcd042f360b79c9883da0e8c0ed39ab0bf3dc64a59e78751e4e65c405823a9cce5d39f6a2e08d760c475f6988b09272d8f9fa1352183bf07c9aa9d5cf448949dd1cd8b77a49097fdf4dd8cfa1226a953f1a1a19ecba99e0ae4136b437383dfca1b1fc1e0f9c1eaad3a733c59ffbd2213808d585969b86942240b772470;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h63e2a3ad7095ad79b854efc2dd004f9d0faca527bd0a1dc8ec161b151dafe071225f00ca5a6c7f500307d964a6d54805aba3a7ed54b02dc24a0418f57d975e3714149a6830a6de75c79d704f902707ff4af27cada5286e09479e58b78b3e449c0536993a1b68df524527b1513ce55a0c18344fecde11de582af61fe4f6b30511b3a368bab0cf8c77c7323a66f86d1dc7faba4d42fec461361eb8f11ed0e07cb0b1b307e68b5aa8b28948aff667b16345cef114f47852bdb3f1a0bff24021934abade96e8ad95fe7cd7fc2ec2bc758156b1845eaaa2e18dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1bbfb9be1f7b53cd40770518eb55ccd3b2fe4ccab8c75b524a77f0721b37db2cdc21ccab2e25b65154db0fb4c618c04c3246d54581b80741e09ee2e50fd956fed8dfc8b1a52a886dfac7975f2b7b720e89427862854e0f1bd3d3d2b99d0d89315527f44ba68d9df87a63c4668e4287a472717020caf2bac80756d4a7a5985f60a6c972cc2d15f4e9039de41d780260bbaed5a8fb06ea92c897a87cb2b3a2c3ac7325ab17bf0788aa4c66eaeb5f727366a7c501748afe5225dcb3e609e41f6205511931983746814773c70e17dbac91a695f63589151a867d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h16eaf41cf72ed3f69adcbab1482988922db29d700266fa880c44bbeb691e3ed72caa0f2ab50ec3465369f8b6fa608a45bac7da5ca4f4c049d8f60e298ac0348ebe22909f9a4977d7b2af56d425fc0b1b122a5b56db2e1a7163117dfb97d1d6b0400a589c9f57d57925f9417a83bcc8395082e394b906f2eaeeb17ec7995a8cc078f637c04dbe22550699ccf07d0cd8653f82669a9a9af7ccfa51b050600a95601a4193bc5ad7267e91868b28bf8b1caab3e56f43328f3bc3c4cf524b1f3b6fe3f254fb493315b0702e20a78065e3fbee8d820a1f7e2e5ebc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6ab5ceaaa2bdb98fd45bad975f59a025beceb5a9931ebf9b0ff72013b22cbea3a31f0a2d7e9888984c8abd7e1d54418ac2616ad9af77fd5ae03af44118b4c07f2957bf74b6217295b74f84119e791e5141bf68eff6561a38cc4ae39cae62a837dcb9f0b84e621f3de1f1d8c3423d28a84a103195853e060c2e3e1a30b2d3802259e711b22f7106d98fd1fbbbe2513a254205b230837f90cad581f5f2b45faa56c0dc309a01a45b7bcdc192a7d06aa95d434f23de95c804e6a068272ca4aeed97ff413c54abe4b2c99fddc2ae13bdb371a312a89c7dd5af68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5b2461654a0bf3263ed5f293c88d229f6348f97f61d62f8fb408eacb70dcded733b6a9d3d102bedcdee68b09f425192d9113cfffe411f7635867ad749e25081fe08ef329fd956e812daa0c69653c4e45beea966304d7a9b8ab6e338446590d1815a9513f9500437875a69ce2da0ae94acecf7364fee14494b9ead31dd0382dbb65967299124b2cbbc4f946b3490cf588a49fc385f4d166550bb88ba2ee182dfeb7f970c8968b1020c5bef8034f24bd24c88728d30832bf82fb3723aae689a6848f33ca2db26ee5d4c81dd3537599131836025c5b55fdb44f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h16659056e8f7ac5e580d82fc63156b679955d8fff612a8b807d9c94d86d39e83fa168c6884105660651bb0b809e8c9c6e41be715a8dd53b7b7379e253938d15f35a5577e317e80d5f5f8d6010a34eb7d1768eb223e60b48224f3f97283d6d092dbaa111137b9b11e6023a5fca482946ed4e3f1b10521f0028c17a412543bcf4638973002618e939a2e27b7b90e7dac11d37bcf09909258d9de94c5c9dc756001d2e48185ab97f796c4bda3b86102cc8e6c39d7ec25c50f8a325576d38d12cff354cd318bbec921790a48609e2ee2597b116e8bb063e2337;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h10090e82e9c0f0f241da4df81ce21a84f5b9ff0a6cb433b660b9cbf5f56cd5bc56f7bb24d168b6f7fad109db08f75e8960dfb5d10b0f525f6f1c501c0e423abef539963209e804aeb14f1d647e58be99914f4a11857f30f9e03c8b48294a767939a777d33a7eba66bd16cca2e246283f0a88a92b74dd4ffd0ff8eb2f97da759a88d9204bcf87cfa2a3a7304fdda339f10080b31f74d03231e37a23ed7d32e20d61548de5c92e02238eacb5148e51580f094e9666cffb88bd83356d560d0623eacfab1f7dc1152b09a0917173263715e4078c4062e7162b60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hdaec8466f5ab7ca201d02e4de0bcc65419a5665b8a501efbc0e2e243fcbd3f85edafb84df7a886ecf90230a25ed018433bbcdaf879b25edc85a86ea96eb0597c69ae9b9616d5affe388e0b3aabd9226b88cf4848c08f05af84c10e893c9217092843ca209c7ed6a72e1b5e7b7e2752244e5fad511f69068b445369075f3887fa80f3725d5f9a59eedc877b834297a6f68fb8a8fbe8177498814b009c42beb97ea0f635b70ce3af7c51ed95391c14e8c9e4c420a7d596616d4f78d7edd128f29c388a08923341a88422bf8a375fcdee8e27392fac3fd067a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha12efe541684d3dfbbfab10b1c9fafcbc07cb915e6cca9ec30df2bd385cff863de79e2c118ef25c44562e91185e15beb0e6fc3cff84a1c1715967f069090b548931f72d2cfb100c56b4bd23f342a8086c1a4cc06a7bdfde1bf1830c676f1dd9466b8f0de185fa50d5883a9f25445ecd05e725328ea3b3f9a1b87f3518e96565a795ffc5bf0a23c1070f42fb0c4778b9423a751b31777b040e26c02aa3e283fad4ed3d833a230b8c94ce623d46f4f0c477542e37de5c3ff8ec612457e2cdc173b821966e4f193555733ecc3ce757eb068b6b7445059f72d7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h55ba5444e095cdc7a1fff4db400ff96c95762c807e592c9947e904cfc86f6bdbd7e5fb4735fd336bfb145c0b070fe76d457278cfd969a5fd8aff69079816284d2035edab28d2a7d7fc7e45cdc1b3bd72220ae73ace88eae11acdb00a432342cc190a98714d8a8de07daedc452c1cd081dcb194bb9165a29c167ca8d2d28e1511bec83f6d30986f1dd00bca22709f5bb517eb060fc8abc7c8b56efb986208f2aa349e233265f1f176cc268e69155907df846839d4c3cba10d5f1327a20d746190ba41c7f6f96dbcf0bf2f4d8ff61c77dc2297bd6801af9a20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h85b6b3dd3ccd8e341c022aecf6deced6d6161e4b82aedee6c64f4da1654b6121d4238a809af29245b51344b5dcf6fdec6fb702f7862b4f956b5ea9723d4a78f4732deb66371312536dd2e44b4ec832f66c4f22fc318cce356362e5e61c88df7615d18de017501a99f74954ae08dc964950df1fc2cee3275f2cd95482d91e3a7039e298f7bd2f81970a6eada1c60fd8dbdd13df59dbe8a8f3e6852132f8614d38dbc480308ea8c9c5215ecb7ed7a384d43aa3aea5520f2dfe01ce0869f0d8ca00bedfd1649ce78a999c290e9b3d3a61154ca18bc16cd8e630;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h50e9e830c035277af647159b2ae039954362f16dea8d67b2d89a21333267a410eb21f2e5447caf82c1b74669066a7a22a13a99367d65006a8ba55f8366495131a0f4a1c3eb058cb69f6fbfdf21de24abde258189292d44c057fe95989b474e674484b82e9363925a0c8ce7f0141e8e3600d8f831bd99d22711415a2bb12f3e2f80712cdfdb862d2dccccb316aef9c1f95203d2aef0444311a7b7ba81904b102926c1eb25f6e854341eb3f9f067cf7d2b5104293a6fe18b990478f24d1575cfc75fcd54ba70dd0866943016b84e0ed30a60e98bf6e93d8b26;
        #1
        $finish();
    end
endmodule
