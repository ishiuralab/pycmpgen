module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [20:0] src22;
    reg [19:0] src23;
    reg [18:0] src24;
    reg [17:0] src25;
    reg [16:0] src26;
    reg [15:0] src27;
    reg [14:0] src28;
    reg [13:0] src29;
    reg [12:0] src30;
    reg [11:0] src31;
    reg [10:0] src32;
    reg [9:0] src33;
    reg [8:0] src34;
    reg [7:0] src35;
    reg [6:0] src36;
    reg [5:0] src37;
    reg [4:0] src38;
    reg [3:0] src39;
    reg [2:0] src40;
    reg [1:0] src41;
    reg [0:0] src42;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [43:0] srcsum;
    wire [43:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3])<<39) + ((src40[0] + src40[1] + src40[2])<<40) + ((src41[0] + src41[1])<<41) + ((src42[0])<<42);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5664f010aad6b62fc66c5668376f780b09f2a6c2f5bb7e52afcaacb76fc37f883e20bbde1b00f618797ae605e68a4a764ae228d3f701b8158d36d03b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78695b506d67c667b4fd5408343a8c4fec0a800d79c46a6335f8315518d6e2a1537fb00e0f5fdbe966d43c8174725fadf4aa5bc635386d9cd5dbbae92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4797965b7ec0d618f531fc261f421c2412d206f7b6774df3c598ba71d867a9b2a3644c1f5d81f2c6cd7832b417d06f8c01cf5f7ff7da8a11d8b49c4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h420aab7f02e13e3e4ef23a7eb66709f7ce02c1e34a75001f9736715354a176effa1e9dbe33ec71ba820631b0a79241e90625c9c1c19287dc48b91a6aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h891832bbe63513838d5b900720beacb1cd8048b0f655ca3abef7b95408e0720889a424c927b1238340a05308b96ca2b1b03a227dc661bf387f29ad560;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6629b6f53a218247ea3725966af65148bca2f5bf3e9d5bd69428bc709f0dea84238be731bbfa52a27a2e0675669d2cbb7d3d3a5ce2a24ea13b9582428;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25a35d0f3ad9582627b53606e92141dece7405d1305b1b85b9dc07c5c48bc1fd48f32ba7d901685dbfd79b51e7f96e82919ffa1de738ebe3acccc9238;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h450167574dc4c2ca695ee631c227abb42b4a4af7b7216ccf52db4febaf15d791f16a05f1825797b31a952faf7466aac44a48e41ed4ae4fdd1446651e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb81e0eae998a1c009dab3bea647cd0519854c6ed5fad058dd281b65a694552c160508a94a7f2c26f7a0fbc4f9a55563d43c9b80941403411c6ce27f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c4c6265e169d411917447060606dc532b9aa7c54bb46c276ff01b8bc0bb7a13dff379e44747f5d49adc9f9c25ca8053057c6855676eb65b5c5e21dc8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haace481d5cf1c1182e4c3b0e59ba6329302ecb67cadb7c0299076e2e6fde79ef33430a84b2e54a9d9c72b3037db8b98889ef24ba7bb88417a3b22f4d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h694ac4c33f8ff6146e48aa159a3038f0d5e100bc7d6408653e9d41becb13c3073f1d8119cc3e3127974f52f4cf01c1fccfd3c83415793967eed6eeea8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34970643e0ccff75559ef9e95700fb4253e60daea38e408def355181c6fdd08a70c321110c3e2134d7c000f5b3d6bad18e8778a341431baa457ab36ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21c8da312d1e844183ce13343e3ca0da61e3fe9be2f8a5e86aace6172adc24ed37000eebc05ae928a5b72bb28fba93e0b1c08bbb44bc790e91bea8f08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h664347b41e6e40c60403a10718972baf248999359891a87ef293f177aa05bf333b540e4c40708be8d7a2d7f98a7bd0536b6394c0de7e8fc6426fde7ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d1fb747fdbd2aff17a9e863619ad9df5a099ff6910aca434eef96ff4e8072a71332cee8a4e3bbe6c33da7eaae5d24611f78cde7088f45ac6f27cfd90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14e5a48934678a2c05de2cf45bd2f759b65b7c3846ab9df4862129201631560f3b4ff3fec42f0624f3ca0414c5af7d37e1f476fee7066dc8ad8033402;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b13b2ff6f51a300a25eb358e712c1d1467b48a35200442f6a2111bbc8729357e91a6586e0401f2ab6d1d18f5c7eec589574dda4a46c4115a1419f0b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41d4a7635f3fa47103f975ff545b8214d5dd41953ad17b75c6afc658f2d6269ea9b3c0260b57c058dcbe50c873cf1e2ae5b691cc3eded8bdda5c67cb2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b95b249200259d6a4cd6f1b09c61e47f39cc922905b5eb1865cdc7627e5314004a19019ae5ed9678b5674885ea991e7b45d0f8a6cc03578b2f223669;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8c96029523182b60e0e8af22281d55ddffd6a8bdc6182c9fb23dd4de0a049609c4d7f587e5ea836b8af9712898800fd1706a493592912d38072e1967;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedb3693897cd3ab01ef5b14912b92e108d24602f2687e849e26fcec6e9a988dbe1224fff8df4b89318338e661ed2e3054e96a6c3478d4a0a03390de4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c37889363fa2b3ac108e50b7bcf291dda89481b476f34cb8405092848aec3cf77ce005ddaa686a0ae0084f026a77d8b0226223fa2be0362f8a995919;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d3ff8b893f60c090a1879c1e7e3828955aa53412bc7b904afef61178edc9c15c97486c862dbeb51b5ce7bf254a1ebe0b561b1052849f47800b5ac261;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49d61355c372a8f25021a19f1bf561e52a58b682d2840e367949bcaac108964d1a4c5e522d85abb37453b24d50a70a8dc705f4e28ab3c4aa6bd67a8d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd322bf757ed77c89834839f38dd6655c71ae376072cc3da68f1f3b237f7622864bfb27c418952f8ec301b20b3f377ca9c2726615ef2e8e48a1c34c54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49dbbf3754c2cfb97e22d9eee40a13b450e96aa3e772204924d24685c4d708e379d23bda0053ead85b0d1babcf04ae2efe7652b583a764189b04f15fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h563b89771ccab51cffb0461f73c159780d64b5af2d35ed0230c421d481f9406afcb3e9966cb580ed50c4a97bf4abcfa2ec0650d1cc6a20e169ab1186e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h570a095d98b8410c1bcf23ea28766b9ba3c443db329de453b88df169f93877cca065ee457aa1c00bdba1d92a7f07ff27820e8149582d8183e99cd8060;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c9540fafda020c2fc9e35dd4e599b9e33484c2288b6627f109212c8f526c94339605dc0c602b749eacb87c801a53f30ccad3101860da69638b12bce0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e8b78c7f69d65e2b5bd70afb0aabfb355dff1085fc04f14d1a3a843c358aa4adc2341c36e2dc7a51659349d5b8139b122268605dc34a1b7e72499b54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c3b7757fb879a0d0dda210c831ac64721f7eb8226fa110336f6aee1967581ad8d831933fe47bd4ab7ce8eef0cca5f275c72b302a5e60e83095374d31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91d133fd49cbdb7e1a54185695fad70e24d09876a9359e37201a4b38c718840f36f757cdeff87240a1e8cba1921973866eaaf2600a75a70990acacaa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8567bc5ddfff1d891751856792944a87629b3448d53116c3ba3a1b6cd27b9929ed265f937c80e2e4ef83a5c14b2cdd1eb7d3b7a8d4e102195c864a82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a0427bd735738fd6e311d4667f951344f4873aa90c9242946c6ac462df04d4e922cc7916eaf7a92bc7216f6c06fec6e47df5c2def88b1ed91782de7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8951432ae5bed951f64918ef61b4cb55a6ded2c9f8387969e1433dee68b8a111b9180f84e1be3a22a3db39ecec62b4f968d5c76df5d8165c26fa95e1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha04ef350369646d67745dd44867d58bab78cc4f987c0b7bdb42392a28f776ea2556168be0e898bc442bbf1abab2c8a47d9c88de5f626c49d5eb850c8d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bb4c4f556e99c415276d4ffa0936bbe57d07f24a68a8a42272a9f768ecb8a91c053f848f8ebe678379b9d9f1c2a1f413c0e3b653ce44c689ddc39e85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c8dbfd9b0a0aa25fbc5eb4b3468883f78de86c9c3eaa62e1ef00b44640326737f6b7923c81c45d71dc773a67580eb9b32020774989ff79208043c2e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b1f552914cbcc31e98b403692e45e4a7550b45130a565676fccd9cc1f888ae6158445cc8fb55cc88aa2a7abe221102ba4f029a4ac48a00b505de7e6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23985246628513d9ee5351182ba16b6c469dfd7a1f096c21ee0eb36d5d4d110ddd3bab8aba5c028084dda3190d7cf027bbeee073b5e9bc9f5e480f298;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3c95fd93bcbd2b05e84e8cf9d68bd9f0284ee5cd9a3f74dbde4aeb041bd4abb0190305de82c9fce914ece271d74784dae7d557e235999af79a42c4f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hded92c2ac843b023a08bc426b278d40e1d02932e7e9f811e0c896ee78bfd407859523f15ec52b4031da9bc2a5262ead460948db602c49a8ada4df6dda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9642f00dc5ee21b58fa5f02f9eee37065f9ab65d88185ba2aa34872820f3084dcf8f81a48b21bc27bc16c9a8cf2f4d4dcd35cc492e9fea94b24ec57e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbce4f182bd0955b19d90bbe11d5b2a7215e81eed6bf918631db53f976e4e506ac5862dc911c329544c434fefe58bb07c353bbd68cc9c1c2c46550985;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf116e30cdb265ebee6f921f3686ee706dda7c5fccd9ea5714c68312dd5ffe87c66475653098c222644d16e602f2d6a0e3a4051f004fe030a1735ea18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33553a5c666fb4ff6c6c6f914082f36b226a0132433a9165cf8fac563355e9685af5f0c5d3c9b671fa89aed03d0de695edef3e6b1034a414cd2d35a6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa2fcf2e072588bb9782c716c23958afcbf3937952b48f9a4df06a0f78b3da677a8e402dccec8a9cea49c771de3123685a9f52e3ea1cacfd4ca305ebc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c2a61c045c6bf0b847ef195ab2622a76fad053e2a0e3d8ec71bfe5af82b4ee4754324c29086ed294b24b4e13cdde7791dd2030f3595ee55510a4bc47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbffbe3f5daa84fb7e013f6e172857abfde3c86b55f620e207c17bd531cf4c571d0b14af087e5c41ba16783a31971d61c212c7b9c54054c2584d2264ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca4402f07ded8f91a96e9467f6c31d96c6e05423ac1bb57ec7a3dd71ef2515677a1e983d749006357bc353b6093078f4ae8450a9cd9fb0bba469519b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h631e3fc1796092c6c2a044ebf4ac24303412f37b8bad02097b46700910aa0a8134295b7fe3417442d1632e034d8ed043e2caf975b468b331481207027;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32e5a72ba15f4914496f6ada8f306694f9756ebb2454140f74901e27df1a0390e7fd19bccf5ec0f35b65be38776e5bbbc4d3313034f6108587378796;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacee341322e26c849346bb8e0b79425be5552729dd53ae751a1f9be94349849e42c9ccdd5e26279e2b7aea069475173872a92d18e05ee94c4e3f7a2f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac4a5ce0770fb41bc5c8d7bab10298ce02c36ce796390d91958cd40ddff4bf4342382e83096237bc2f62fd7214460c54d982feb6d91fd2c9740cbaa9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h649538a2db602b7fd3a0fd7593c577287397e50a243cf20342ff4035121eb34800f4356a1e1235ecec9fec0e959aa95f22dac2597c2e2ad10db36a719;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd62de0720ee231c7cd5c6cf2d591b16bfe6925e787cdb4422d42a4d03f2a3b0381433887dced45598825cbcfdc2a2c00e246ec29ec592176add2eb0b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3c1786b65a27ab160a9c4622f79afdd7ca235472ee52561c8ed0049d8ec67dec0ab073961809ee978b407959fda8cbfde972f2343121dab5420f8715;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7b760f6cce024c3ea86ece0554505d25eb7f2f1d4754421fb88b72e6e66700ef27c4645b3173f53b9d1eac50dd63af81496c3e58fbee0c8a82dcd385;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93958a261ae92de5a5e0b1f92359e978415846c496a2b69f50b4197b2e6bf1c072dbc1a91e674a82d5f3a9f36516c8d7c5ae776582ce25effb49be357;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcacac10a3a574f8cbe9b169abe044f0240e4e2442c05a27a4001380d7197d228a928f2da1cf22be8ffa2566bd8414d6e90fcfdfc5c4a5ecc3402baad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1564e76c1bbb5babf4c95378cb8244f3c9cca628faa559846d2cf825e5398dce0173725535c7687a96722f977188247a862218808579dadc091aa16a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haeded6284f056f33c6d1460df9a40625e83c2b06963a0a17dc52a210d4f498c5fc7cdd7be35f952f7d9385c6088a3eaa7f5377e2dd57dcb2b72e38308;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heba8e1a1b5d9673a52423664eb23d76e5c937ef58e2964456f4b7373a9371232eb8431d3e7baa09ac60b2174e6cabafb5916ebd30ea0eacd21e636523;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9224b563b68222967aae8c74afa8b369e32f15c8e0a2541bd40fd76eddd1266b11b07136aad5950c95201ec9f3cf010a510311f2dc62edca883a21b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h234b26c3f391260eb25b31623687c418c3b3f445d787b835250cee4427a1927eb9dc0769ba35501aab6638467454ad607632da4fd73fde9a9386f4051;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51361aaab5d08efcd6153d553f20c6a9f22ff7dff01bef33b90986f70bd8fd45c90e3fcfd9bb87ce44f561bec4af559b16936e3b4274326b21b175f45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8adbd62e2a9442d583fdea5c0f27bcdaeb1bde25be645addfcf3bbf131d87caeff2432938fbe5a43410c11a4080632a2018d792fcc24d1edf3cb94d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he99c495958b5ea774ea97df73a9f7d8cae74a87cce43ec94907647acd02bb7201b8fb52d68c5cdea60598aa261c9f4c5c0875087d156f6b327f252ab8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97094e9fb39cbe2207a437075171d2f6614d494b79acefe4316a70780184a06726ca48017037afe32bd54ce3b278bacc7cdd25127335f2333a6a9ec62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ea38f7368e76c787cd04eadaf2168bcaaff5494d355d80827b0b5ae91763f9c0dd42ab4a86190f8b60e361026c2b0d15e0e43a1f3b80ed89c03502a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85ea491f08911b4267dab4b1c1e18865dbf65c76bbf1b45974e87879240a9c5dc8db68234f53044e6dfc2df80ae9fff62b597099ab8c2d0e541652ca5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5326acfda36842333cf146ee8a8cb664346955e647c1bdf1e4431727e56e4084e2c02c3fec38b2c35017410d097dfa78d48b8f3175a53d33535d8b5d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd034eb5d3978258c67e60ae75831a0276e54c79665aa2ad1f4c59f33c9ea0d5ba22b5ffa66218eb7a6a5e51071ace88d4c9ff5dbb88457c3e45ad3bb2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b99a55719aa83c15066ec4e8a1b54f8c73da3ff87fe8b225284a72698280dc0fae829dc017a178bb306733d21b1122e1516b8d2f9c25be93f02a4a34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda2ebffa746e2d96cb22d9e208afc44a63556618eb0409fcad69ef9b6e02562d485a3e2f2fce7a7bd693c817d11636175ef2c541f2084fad1faf963da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0550c0d3ec9944ad53d63c6ed0f140e0ee56034a49325bc22d43f3ca5127857853c52a3e786f881358add0a452060f28651b2f297a573968403c6f70;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7839cae0669099bf7a1bc375dfe2a05b1130922f2ad8bdf9e69cfbc547b41f2b00dbbb711881fd37c040f50204f155b314c2113314837e3d8e438035;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbbe0d72dfb71680f8c2cbfeba803fb0a49591e4cf38647ce666e37b1c02ca6c552adb62960abd1ce3164489a244926f7f01e0fdeee86dd4efef31bf7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9f7865bc6349d319044f0c2bb8101908e53ea0be8e2abf18d2850ba8395457d38160e79baa373ed0076dcf03fbbf3fe9cb25f552473d4747bfe977a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21b590b66aedaaa23b531d046ebfcecae7c2f8aac8a9c2dc368cc24ba8cd5de69a8b50baf7912a7150b88bbe305282632abbe6e5b129f9120b090bfa8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h339da175bbadfb35355567c12c97aa702306c45217f5945090aaf56ecbdef58e392cccf184ee3be0ace422ee4b4a999907f1a2d5c2abe39cb41578176;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdba6edd573a0392e075578a2969a24ab520d608d12e57b3852fcee3e1d7e8f69c959e0227544b029a92228172cd6986cfc0ff0814ab391cef46c67344;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90f65c41acd960319ba645c1f6493e586896d47ddb4d2b290f60433a77836e9b9327d5657e6598f7c5c2a28ba463c25932a801207d2e58593e162631b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c284978f4c51352c2d6be664c70718ab7296980223cbd535d476c73f1b4a899e6159f57de26c1cf285dc84d9eb2430da16d5f4c82d8f23231f3b4681;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f3ddd26c5b773adc10824b35d0d9efb83f916e1432d8bb4c9e3511a6873761c0af8f1cb51fbccc295dd22d9dd89afe88fd2dcdcd7eb0067efccc72ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h627bde78013a027c6a8c769ca2366c77f78d368f4915cdc1c5d2034266669d4d3291bf3672ae3049bf5881594d28452527feac42be44e0558c8f20282;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cddb92b100778172f5ee9116248d40d3d94a8ed7879259c509e0509e4e66c110c72156ef744e5c4b5258eb5ed966b15513f577b3b24f24cbfe577ebf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b80edba2665d72afbc5c5dbe6006202175ccf8116241f95088166a00671f329226122bf4f0e56a8423f534dfb3491b9bded1f263450000bb89ac20ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8712a39df8d2db852e157da1da75ca81b06404e8a86d3084a3515c8d43e84f0d0eff587ab7d635502084786ef10f89e759e927f3f85d60d46f5ad136;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc687e8521594d989846f290a7cadf370eca85fd61dea6f1f39df2931efa84bf0dca09fe5813492001319e6ef24e28752bcd7fe497f34396c0fd9a4b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb02d0bffdc1020b73d013056fd365b629541e98d0a5b505600e681e67f944220a4fd4730aa75b9eadb3de6cc0f0cf0451f4c6d78b6e00a45c253465a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61ea303f25eb9621827d0a04c9967bcce82b6e02815bcebfd9ca069282a910b00a296fa5a652f2ff723d196871fea9a9be45231fba30aed00fa638b96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadd327c2b94f981d3d2d6f35c77e87e991d28a7b690f88587e241a54994108b4aad60e75dfd4b830b665e2027a14f6582a2ea09183e3039037c96b7a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cbff54332b6c477bf949e405a2e22f2b5a1d350d8d68ee56f005d7edf072690d265f76bd14cac1910f734b3f4dbc754b3469db1454797ab695e13521;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca7cc1b85480ab1bc939fbeb27ac3c7d3bc00a21bd5eeec8d05b5f29b86ea86266c7a85ed8fc3c5b076091cb869c93cd600cfc94e282b63b8dce59e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2769748ea467b81f28421dad68839d343563e16664b437b9decd42c9e24147d7c2820b42b6850f53230f501f90993c5b0a8060f45483ac4e037640e0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa0a9e4e19883277b773e6db07b551cfca011dff6be1df6cf37d64107ca715d4633d716ff1178115fe58bfa53500f390b77d2903b36a5b5a413cf057c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf396e342083ba48f77b79f7d8d428e92de00300d580fa4ecb0352821835d3e4402d13e0af0d4496ce52305cf29929d23ba99aabc84dc046361f3a3c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6eb4b4a9e0f015d22a1e8ecb91f92f7911fc805b74636b0fd12fc7a4376744411a696d976ae9197683953f0956c65258151b075ab180e5e9e0a291743;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90552d18f4368f26b92d5872f93e90cc08bd0d630bf57312c10927a0d6c5dace486a235ab155b4716505cd776ee00d40abb72b5ef4531b66cd09ac50e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h156faa6bdb157a422d6ca3cc8d75891b62d0710828580369d603a18d229794b7a5c530e067d4bd46753fba12116fd8b3fb5ffcfaecf9d4927ccd69c39;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5306bdf90624cd95d42b0f7e378ea1deb0b269d33e541161150073246f8c3d0bf0f9f4f5a73a2e295bb7306866ebc092c681801f7f5e92debc56e854e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d1e40c12b32e729bbaebdf6cf9cc40a70af6a8d1d5d56ce3d46a573b8d749dc6709226c118bc2b1538b869b7d782586a131d9c95fd8c74768a9db2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he189d721c03d2dba3d02df2cf83efb70ae53556cadc9401fd61a4af38e0394076c3876f84ab347528c8368f7fb5e4b9deca4c270886766e0c385afc53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fcc3fa4270b1f550df240da6814ad0f566385f6eed788cc9adf543726ef006bf7c6becbaa242f786b04bdfa7ae82211059f40d913af69530b5e8c7b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e60be4b1b87feabc550153ca68f0fc58114652aabd3052941dae629274f7c55013ff2748e04ea9fb1143eff2c52e4a7266d2fb85b8b14dc68eb89519;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe92289993f880a92daad02fc13bc4867681234a949767cda077617fe329da29c752d1d4f5a3a75a5f559ddd77d41758c7d650efdb8f681bb6ef1046f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd57e4973b92f4b306b28775657b087d0322355394e52bbb17336c7ffb1d34fc80705d5cedd8d143830baa38b218c53d2d95b7bd633c15551c1d4c0625;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81d3b7fd01e982ef559b0f80ddab3d22d2b678aa47d5af93cfc6374cd0773b141c1e55e13a27ac7775f4d1e44816619c4bba6ed6f0f7e89c5ed80921a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c6be21fbfd8c00bc5f2bd35ada14a2d05cc602b0178b4167e0fb4eccabd78cc3f6375d3597d4c2a62ea91e29f9f256c735429d07a9b994a0150b3294;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15c3713ab4c3a7769c203141cfff6d81fdb6c70684a3c1caa06cb25eaee3ab7a50053cbb4068f5fd69a1a80ad955de11284b5a0a5b31d8fdc5d6a008d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8fb5de6bc7a5223f5e9c11485170cb7f53e7b1fdecefdaa2a46237f04632949fd1f03229e1fd599567e474674692dcbcc67191d9cd70d1dc0a80bfd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc603d825f71326dd189fd308601aae65c502712474221572fa99863bdd5557e30d56cdf3d19bae7bc7cd5cf84b49ae1e7667a18de8633b9bfc161cfc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca5e0a96162d6f52be07b51dc14c3f77c13cc5f4f26f65a8a46ae132477f9630affe857d266d95561361f54c9eb770db3a7f4c65f0749e9cc43ef5e02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fab3a18117e8177e80f53a8391419fdb769a0a2eee81492ae0b34fde738397d1194744de2201a618b34128526dde9a132348cc718009f8c7316b220e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h172d3850e727d1fc37667898d7dc8ebbe30d269deb88bd028d7a573231f054ee0753e524b7347f4d4dfd5ce736bb3bc4953c4547d23a11bfdf3cc418;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cd43411bf5a3811ca92424d3bb7f5373268ba3056cd7b24086ab0daffe0973a947c5b016802b5f33b9f03acb1769a286303a74d747d1f309d4f6fb03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he271f92d751c1b2e714ca800e7156061675360eb09469386b2c9233372bf4c3495f4b8bedc8908f800d02e078813d401c5562c3d2fa35b3129f5e0a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfae6b454f68625152451de0c70c7408e60f00520f9d06a4da4c3496fcf3df0bb95a4652f1fc8af352cc6875318a804f1fba6470709079e04466908a10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92163c0b6d47abb4d7b59fcc35a34d53708d9ee04d65a024899c7d93733d0933fbfffc55726c4bde6142db102275682043b26025ca26ee9fb87bf31ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bd8f083086ada49205711931c07b152bb0a5ea3178239d1251d8ddc1d164005e379cf6b8fab47de65c970d363480234e0f117dbcd49650a0f915a665;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haee6628fe1793003ead3c7aebc8cc403e821f7953241bea15395b3e84a7557f7936ffb1788fbb543b48c48b33d217751453f87ccabf7f92ecde245daf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7522c29b47626efd123c1f396e5988ea4e043de7928092948b2dcf35c22dc46adc68254bed8e226127deb930d42e947b31dac550656d308013fab8f63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26c97acef71068fa7d214b142930850fa3f1adc945533bcc3bdce06f42ac7fe211d5b9cd1abdd9a27e44c867d60518c4cf11ef4a826d1044e00c36565;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha914cfb1e3f96955cfbf515d1fd1afabed892d1f492b720c7f6d9862746e96a3a7ee649c43a56b574e2a8fabcd22909d8eaddecdfb75ea0dbc5568239;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3254199e99a7e3e945eb6d943cdde23c508b592160f0a5c478ef9118e547f8b926384c2ae110bfba9e15725a8360261187b995fcb0a3c27518a420e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20bbc3b0e700957237679d5edca82459992ecdc3e5d122e41fd661b4ed554bccabfb17e56f69f4b7e4a088a92d417c1258e3425879fea5696951d1a45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb069b20e85d4b2bc5cce3773ce1c1a19992ed4b7732e3603eb5d4314e04021656d41a1d6e10ed4a9ddda84248cc1a494a1efe30620557fc08cdd26691;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h982afe91cb156099ad29bbf58b4ab6ca8b6a5df7c5882cdbe6d38f4343c5641d75f7440ddb296625652d45fc64f3310137d302103d9d977f68721d477;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h445c140b739a360a8597d4e5b3fd97dc6020411890e1d2214dd49a06363a1e6a17efab5b949c555e68be38776659a9f5403bd945c82d1a658785597aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h701f71b4770c7f3d7f42db0699c9b5d1409100dc1c1679c58aad0f57f436c721b0e297c1163c21096103d088ab7d18f8083d16b15fd8224208f30602c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a481fa0e66a07d98df712b4ea3a3a18faa02dbe12a4a8d78665443531188e6a98ba675df01215b77c8641f583657c504547ba179737d3e5e929ddb03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb30afd463019fe45f49269ced7c0d3f6e1cdb0c4265b8dcfdd0c90259b0093e5e94807363c9f3f2e51db94712c02b84963a2266459e06651b2a327ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ae9ebf0ad45aceb2524b115265f6dd204db27a53efcd2d406e5da71d514d5658db740e1f48ae576953f00306b95ae467d36ee9afea3140b59d3c4430;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf293bb4def023f1589c8f16fbf42a23784d35e0f79ffdb8b432cdcc8e644c8c4dd01355ae0422af631278f54d50d83b02f02975472ec3c19175816061;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cd55169adbe7afb3def4ed6d72f2c52a8ad25245bebb83039b5bb365ced6a2c625ce5af4e7e9b70bac963453bf3c323fde35760634f8709ac1c3a00e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda982e5233b75691bfd2a2f6d4e492d32a61972015574022c86e336a4ea1c40aaaf652cf9f8d10e54df748ec4a71f90c328db4b6d0155f43ca31fbc07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d0c133b14f50ecb46d68a080f41a17f4b6ce4293f1fd9697cced85979b8caf503c87b30b5377fe41394129b2fa4ea60027e9eb3ff5645505b96b4272;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde9d7c42ac0a0aa26439d22b56d09a226f434c577276c67e9bad6adb2cf0874f6bcf4b13913cfa126f7ab9424711aeaf50589311c2507f305370d241c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60e019b5d6065e63cc17e6eefde6f27bd4f45fdbccff02b2cf26a891cf3dfe7c9815e3546c35e4ac85550ebdcfbd2d7d5e613d92711712f6209d14603;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefb96671544a4107b65b28b461ae88211038bb7589d5913e884d46d8f19153100034c3d4fdd9655936173bba952a1cd1c626a31e4c4bd1f64eec266f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbc479d313fe301d65901d6191f96dd83920bb3529be8407c5a6e1fae2d6e87363ca8b4517d582d02e19ae033bab1364eba52bf82bc3918e87f32f4d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4cc4ecf205ec117019d5fd25a2203ae911d8fe200a78db115b3f952dc37f0501f52fdb657850897950179f2ec7a90aaf682eda177b5dac2435fcbf03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h490b97d75d379609651aed638d07e71104d073823c265d289069ce04d22424c916e263b1f006a8bfe892e965bfac00a3a994967a722545b2f1815eccd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6289d3aebb39d54b20e69d3c694f19d1fff4af61aab1a1677de7389459f8da45951b80303e4c6673fc60c57132e0084aa8dec6123d7d8362f8752bd23;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h535a2fdfb7824015abf57a619c3c512c633eb9d0f932741090701ab5ca710a2cf7dc505b4785533739004a2f7eb635af12627737e8f61d58162ab187c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94bf340cceec57d2e9bea884d10b45cac4339dad8e087352c92ab11db6fc0b7a67af8a7f2a34eb8f8c26a18af6c64702793bbb3f952185dd095c4daa6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc02ba98fe10a7b450d703677c8de8848546564ab402571ae0c71f58454ef611cf302e8e57aaa6371056aec3d8e110c2b66caee02dc7970a85cc6e6a8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65676c2610defe98f9edc2a90feac8c632103ab10b3ad3dc8b396e3b8336633a56444a425ed0bf91e9d6dbcf3ad2c96782f0157e8e90f17507710842e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48fc953f76d7f3c21d91b586ee4b407870c3d306e6a4581880ad79ee20f2414e99f5277eb957b293d1fa33d6c5ac0628abef614bdecaf295d3cacc5c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d1d2b7235de43cf4c92a6a23f4c08901105231f959625110fc5d069dea8fd18eccfe831584f1aeed142d8b2d57e40e4ccb3b7a7b6ce26cf7e5176fca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3a1e8c126f46e71353379ed1a324933b1b53a4a194b0ed76c9d5b6dab19a15e6abac03a25d6bf051d33792e4ceac8f601d4cec60d897a6681a0d11eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf0dde23b971d3c9082c330414ef5eb022f5c7dc672f64f151a1d1895380b6ad329a8cb0f7f032710b7bde0ed84d2227290ce660a42194e06f00118a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fc4a16d79219620325697a11fba1a477ccd57fe559c6859eab4e719a8575f397c29fa72e9dfe9ba46bdb9144f270c5952bcffe4fbb1d9f626918a097;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a7825509dd44d2f3b269974b72de0f6cb6e2ce53b6b272451eac8dac5894d76d0dfa4330d3f5d72f3ad03e2fab7a056e10020653c423aeca1d00a97e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b2260003b404260ad0b86219ba48509b06ccc935b5cc07f425d0ba56ed502c44defa5de0444ea840f8326ae97566b0c598e0ffcdcb783ffd57f88244;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h143dec38202650a6af0bf498e35b78b58af75166da7b34d543916fb00c2e4379d9cc5a56aea296bbd8f71ed977646e58e5fd1c3547290b6ff74684d12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99cd637241b59c873a45209bdbe312fa363cb352f7eb7ef930ceae6c70f6640a1e130e99ff645783868090238a0e087d7e60aeee88dd3eb9817dbd479;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39727a6b7a3079cdac2a164d7803e2881c7b3d46e46eec983e02ad55ec4c9c44bd633bd3ec0cd664aa465626c5c16871f2cf954b75ab075fec624989f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf529d7f6367b0e3d95f38406a463aee9b553cc135a36bd6b1ed954cc2f1456b508d812441ea80110d6677da8fbdaed72c26e8e0453720db11fd9656b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec19ed807e1f663ccb5157cc96d9db4b413fcb42c4e77bd5e4c58d835a7b8b99bdc7dda40b5eac71f2deaefa64503461400e182e242a435247df3209d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3bcf46cfa94a9df1b77fffee6c2032cb8ac777f7da902c5aff451e8db5b83651e0672524fbafee1e8ed89267512490200c65d05607381d602fbc6c44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25f0ee08fea33641eebdcdbf56e2aa707533fe782dcef8a2f579d8dfd0bd4c288ca64afed8b4d284093c166a1fdb0fa314b445d35af5a6dafedbd2448;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c407d380790dd60ddffb177894a3508d2429074db08c159f2f7fa79aacdcb4bd9c0860803bbfb4eaf86941bedff4ce23d151ee48c01ae7ca00635ccb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3ec926c2632e14dc7d508e52e231cf8b7fb30baaf757228cfa1135687bee00d52807f0063099055ba4111666b2ad1b7f2de8d08bdf299c470041f156;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5418a7138a35b56faec97b704452ed846d4fa2e35335a013baa664539daa4a0b97d9012c95ffe0c35f338ed62e191a5f39704ea6693a4bcd796257bdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4212e4f15e6756a7b83a80d790beb0abbcd2450581904d87da4bf16bdbd28f81a55ab7b06f1a07b07d72e4f443f23c4608ae2f2e69b05898245347085;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1f613a618cf4f17cce7fa881c4792b7fcf8cc44aa55857cd4fcd13e000cb52d5ce63f8d31c1ff324260fb620d4995a7004be2b3771721f3114133f8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddd922d70508954608c889bd583a750273fbaaea12c496d357d84287e4974d0a5248e3606d0c790d3783a33752ca49e2b58e89c8cb11cc6b7c975b1ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd295d6a2b162c8d800be555c7c6ba1cc729f6b28315eb367f574d641c0cf7da9dbfb55539860a7a310213c7a1c4c7daa80c6585b698bab8fc061a76a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd227d64d5e25847d6fb3c4ee63a44ad82fb26265e5df3ee4906ca9ddb78086cc173987110fcd95acb5e7f66b0331ee436743b228a8aaba8d728b237;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e6d2c6bd6c8c5ca6d29ea4819e4c70d295ce02d868d3249826e220d3acb4ada0fb17712671f1f27f38fd5a1ec5b738cee9d2a42f40e152fbea8b7724;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dc319797c02ad08a8ead63842f5d4e3b22cca4644c68c719c662f18dda873edf8f1d6c82e6dff4ee83cb80460be21e20dbd72238f018db5d9a05999;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h892810ecca6709d22b23700b1352d2c4475c6aeb841cf7acb67d2e923056960b46dfdb8bbcb2177787816c5bd3ebec3fcfc39d0975d01d4cf3fd4a315;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a382d40743c6f3a22c04ec23582ae489613271b84d78ff8478f5a10b37ba6ce6fc7dcf9210a8dbdfcabc21d0a55e11756cb6a6cb1ece82bd594b2459;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdac78b3514ea6cb4300c3d1bcdfd3cf0c0a8969c9b8aea1dd13d8eb3d9c527799079c3a970bcc210be1c5fe57dd97f79132f28120e8964ccf9635e0a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7659667990d1744123839125a8190147eb94dcaec48451178668065abfbf3ccfd6a431e7e290b08949fbf2d641d1ea91c4ba11c2fb575436453df8aa8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3c29b2b47477902f60cf40c6d0c656e16b30ff4a9e9db74cd6328e922e6118947cbbf1448cd79a01874b698bf909185c7a42c2e7cbd1baee5d2a1ba1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha868156dced7271ef020f32ddc0fe9bf1fb4c757efbc53d8b7ddcb08f8c39f0a9501af278bf2046bfca5f021361b220a88cc0f76615d2bbc636e991f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcefc57e95c84c61db90da8727e8b9f1040de430d2807771f34b21b3bb835f17a652c3f5a27795ef56fd5f9658ec5ddc46cabb27b08d17f54af53acc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c501376fa6851b21c7c4ffbc813878fe0ee01cf034583dab259cf442c9571023b9a4ace9d91ff7a3971790123fd4270a0357a1111f3e74d246f4fb5d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h811425f1b3dad03a1c356e680ebfae05930d2c193663bae19b55bb12669b33fe428a02470901ffc5080b538da1c4efeaa03b12171cd8405b0e672f265;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb80e4af092f55f6f90b3a951ee7b49a8e76d400935d22552931b930bba04aee3907c1046c1c3bb38b4d9ac4c6eceb546311611bce8f7bf301de8c890;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd23e67ffb274b0180d108bd9a53bd0e51065bb9eef9f8a672eb17bb9d3720cb043a1c5ece207ae81809d03becb6413405b0bb501852e84f987097fdf7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29f672b7b27e5ceb688e2a5b6026535d3d8d053e3145ea3d9c00b114df4cc7409e0a1d3c8243f684292fe4dbed658657153ff929eeac42d4ba20cc05b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha25b98d6e847a529d390b510094f5a3126cb90074f9179a1c44ec7e87a666096b3ed3d87afabd147913d28d1febf8241fcbcae7887f364718a2310d72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfef83b1b59ad2bf85b29776bfe9041db64f80a07e19c4d39b33fa5e043ced9b76c1b16d523d849b1bfeaa868021bbd67e78c008740ff337af655878a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c87d57edd107ba385e1bda391d2685acc598b2bf679fcbd83d14c2bd83d56963f2739f959077fb9e276a9e4bb198c106e5eb3424973def21b3f22f37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77104bc246638f1316e997986941a6a58ab6d0fdbb9720567217866cb5272c8fc03542075358dca570c269deb78c67fa1f840b6e2182b3c29ff766d01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce50d6681e919efe5a4622fcddda5fc0426ea89c5b5f69224174f236d179d6dbb24991ef0affffe68f97b6d4e41fad7f94504adc8395396b48776fea4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha89e32b23a8bff85a4c51d21cf698c27f66b0fd86e1130a2b3cb3f18a2deec3eadae40cafa35348d168547b54b86e7b45d75e786b0ec98ee7104a95ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8e61dd269f680eabd4896ea7f0a67d1d23afda601ae56ca495339607285beeae4164782a1a290a8f36f3a9afa97f7541601c7c06b4f5d031f3ef6e10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha507ad55d5a06723be661619dfca8fb33b2e952a173e5dee15550279a3790b7905e308b96b0b09f3f36ceb2aef3a2743c18dcd72193095938fe0305c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbccbca34e10539255bcbc6719e884e49dc28dac6948731e535e10ea6b8b7051c45f6bfe964782315902ff7abd2c4f475df7bc35fa7398abd476bb417;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b76bc0ed7624a6fc67414f564c4ada1f932faec82baaf13f694f162f2135704a64711a948b2dcbe4d56257a1d5ffa7c06f49afec8f920eb64930fcca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd973a75959f85cd157bff21a8614d62611200aadbe00f844716727efd44faa250e587e32bcdf2e4a75062ce274f20ec0038fc09b7815181db8be353ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4a35551b337877bc6ec27c9aeb3ddf234fc322a1655f916537bbb821e8f86ea8b64d50439cde9d9fc86ff547e737bcf949a6abadb0484cb3558bf85f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a8e82c7610424866a430180060c29fcc6b7e2f32cb7a16af53cc81c5132e063e8ef35ac1996022c0e2cb04df639bcc4b9acbd38533ccf0003a1eda1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h537e65423dd004b6a52de0cc950d928393583edd383b3bea94396cdc7a9c9c83a23c19f48f94a5eac5571e0402349f023003294df1c5cfa9786a9fb32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb26642d3edf07e4bfe9828d8f13e3a763f37bad72cc436d73cc39e68188fb1605667ccf6544299672d318129bb975b66c4cf09c8010fb8b7d37862f5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ec8486adb3b367e27f70a269b6de7eeffcfbdf7947ef176e6f15436f614ee92b9b24b7ee54004462bc7037fd87f2b39c4999801ba44a536bace662b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd70f1af295a69cdcfdb720be870c5c84c8969683eb793069d0e96540ba4d8a1a36b4ea06cc2d76da7210df912dabd4d8d1b8068af6ed17176b2ee3408;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb5b72692ae07e5ff6f85bf5864947fad92ab1e052bd244a67a6592da089fe0f7169e35197b6fff4b7d2017cf59500c6ba327e5406375b3f6c09badaf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16a07898690403c37d1efd8f5acc3e993ec9029a4b3c7bef2898fc12ac6b86565ce2bd89f8ec386bb3385070f42c99b298b624ef1097c6cc0f7c7f54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35a8dea4b3310eb89d88c4c8735e8d5861ec13003f60f3a49e3989ce7dc02312e9591fa6b98f2049bd35328b9af4826f1ea7cabb9558a59518c6e2ac2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8185b574cf5b3f4a213d2d9aba11186b0bdd645f2f48f024f9ca3b5f41378da40139a2a47ae370ac9ae452970cbe07c456a23a168072c03ce94a5a4c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd2a275555ad6d2facaec68f999171d228745e09337b65a3fc0c1ceaaf646108597101bb26fe4de8f509255f2236857a215b10d3b025aef76942532;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84f04d52990b4076bf3255294ea4c148bd1b8d72c51438f7bf9b6e0d10b2afcec079f62d089de5635ddde52b2697967bcdc64f623ce820e83fc29fd8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6876ec4c66d9755a81a97fad7ee322d605d02bf8deafc91bad5f34ca1d642ad125d33fb1a9a5e8209ca46c79013301eb002cdcae130f9dea9f6a460ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ce919f1f10afdd1f02b3cf6c69ed97ab26b8535cc2a2388139e243aa453e173c3cc49f818a9386e71ba0826a79173a5cd0feefa6e50b1127ad3fc542;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ef7bf3637ceb29af01611b1dd8a2d938ac809b560b0e00b1c8a28d33f298ef30dbcb8a6b8f0b5f5713988128f2d814c92691d49c926e09191ea5ba5f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38a363b13fc14224c5444b7a5e63c97b0bd8c112ab14fc866bdbd197a5ae942e31254355f495f8f519a2c0c62d53ba642292335381abb2c65f697e1be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc10917b123385a91f1bb48975a7e885b8110e1f1181ac15531033cbfaa08942a71368f13d3bb8c4caea2b7d3c1179fd25b2412f9e2a502dfd983423bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63143bd6cb7dd213a6f04fd1f5f01b8d442d977541f852ea681526f3b5fc0e17e3b25b9ac78d802d5d7d5df7c85a5f4192c7d319b533fc76e38679164;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7547cbdfe2b55b75535686e1874a573e3042c1a05b0ba661ba8553908975479dda20d8845b88ec378916fc51c8c4fe02bcdbf9b0cb4be1f4be44f3be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66bb2151d5208c2621f67564ae022995d4a3544a47911f08220b0b685b8f6e1ca4ef237cf8d6d83505ff42156d2173557d3830854598cb5b44fca4716;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd128d2f7ff3cc5d9ae1315b3324444feeeaba13b552459b2a94659bec5e6a7222b833e10e1163e6e6954b1da122edc03e05ced05cf542987cc3ca57fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6300c122323f1941f02923616fff124dd85931ea7c64ae4ab9510778060cb340a1dee02862875b823163034ec2a3dc9c525b774bc86e309015d344013;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4d92027ab7338d419a7334607c4b09fb8234e8fd96a40433cff10167b5c115ab1397cdaf331c22f4dcbbc2c3a10ec501107bcb433511e5297e3dd8c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c778ec3369363fb45f6bd3bbedd0ec099500177800c9f4b0156bac94f371ecbe10d087481f5e214398366990a77b76b9e3c4714269929243ee0e93d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8095b1497476c78346e8cc42bf40f903073927bf6766ef80b15a0f620ad1c9939fc93cf0301ffc8d10bd4d11358d856e232df0cd7e27e4e88648f5530;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habf2a91e672c00f06a0c0d01bb5060a5a50ed84c8f82e8780114903f80366a2ba767cb3c9a4188929a199be1af8b53cc65f37996af231359a4a9d94ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h104ea41d18c47f85926d8778d047cb0dc29210b76fc29e0d9dcbd1063c441048415396e426a3d3b5ac6eb78848341e1731706fc1ef28196fd55c5a493;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31a10a9044bb1cd8c2bcd986befc2b40752a4d3b769f4d8375c950723b9d3e6293e4ebc5ca9f76883f72ec6b131e19c06520facdb8a2ef9deac5a5d82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcac3b3a2354fd7c2e69c8a58d1665ed6847d991b494f743e1e7fe65593f8f1d2ab66ac1ffe078b870929d867d770807d31356b742cd89d662362eed74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h278584703c65f7a9ca8013f8a9504522eb5bea70fa56213faf4ac96a072c9eb9ebcee8a77075167f1812ee422d0a01ccf0c3620bc6a548b59b39f800;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48c793a37ac639d6117cc992202a64cde409ad6ba0518920f0feb06d85b1096e8514d51f95e245432c9175e18356d2712cacbe69de04e0d63d2a83cd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h252a4bc71061dbd82e9da8ed7fbfe155f9b51e5ba0e7ca1c2799248ec2762041b078afd5fa15168f5963a52418dcf3dc9ef457391ea3e01a6267a436c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ea3771f6350049f36f2b1af33934d37ce3383152e43474e99add0a30bf6d78784336b8ca1fab2cd5683d86344b788c36c316c1374a603edc1d881b59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3d400bf29174bb7a3a59c3cefd9aaf2c6519dc84ec4e84bc83dbac8d3c111e582f61e3830249ea6d89171cfbe98a0ba28e7e1190d2b20be1347ac983;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14a1cee73efbb716bbd1e593ee36ff52e6b830a5f255a3aa2973d7530b5d95d74c29ae85718ea16e25dc54f121c85589df122a184162ef043e5365ab0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4a11265e05d5295449b0758778547972e0ba123571242b74d8644e49f79e0aeab58a642bbb03cacab72fcbde3da08ce4a36ae20db4767ecf42d78234;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3736e00ba25de75ef9e9a4ef3f979a165f8aba4a5870b4ea0ce29d246c628886994a2081c87fa6e15b97c6d5f887a89d6660893be47959edb458f2489;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1a821d01c793000fab98fbc5c70cc32d1b259ef55cbd55caae2143c33059feafca8b05ce80c7389035583a958b3210e28c216d1d8b80b60dd8891174;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4008f71d97c54859439755aade6374430245818c21dc23cdc5413bb1dfc374b4d1c73b8d8ff256d2c3f19f83a68ebd2685424b74111ec7f31a3844342;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69693dcdaf7fa2e29cc82e3b166d4761c67cd06f54e3d313eace85f4b0894b032dbb9acdc935f1d69ac8e5ef73e6474028266911cf49ce59f6e5efa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc50fcd66f82edd41e2df58384a2a9b9e80170707da9618f5a20565cf406c368374dccaecbea696c84420c0739280970754d0670760f689cfd6cd4aae3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b98f582530cd7faa1218ed06ec876f7fa90451aed749ccdef4989ba8c81356287af1144566105412857f0bb194d67ea6f9cd790a50b0feb8b0835856;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b44f8d6df1b9f4a547050f195b1122dfeed953a4ac5bbda85856a048d0c289cb65b2a890caab0e6e9bb2509a0521d9a2076f7c3c73b817ac3d638e22;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9c991adca169d00ad38089476edbf4a49b837cc052cd4ea1d3cc483cf0aed5e5756979553dece7393787e455b66560e877217d4d1458d836b4d89423;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73edc814a288dc28ac33625f8ba85b92d168b733a19d0d87ea71424d2fc145f7abab2d0a6bd44f8dab0e6af2c56e49cc7ce6df53ca252e20533a83a23;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e70a3b93dd8af27880dcaee16ef5e68109a03d5348d691e02b42d43ffc27f1526496a7b68eb29b00a09808c249cefc83c90f49bea9ed93920a7b529e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf91cde9b6b4f548b7604f651b4e7aa11efdefff52e2334d8629bae26bf983cd95eb4c0357bec097e6932e4e966d97f53959a30ba632567910be86b4b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h469ddab01a866d41073c5f18557c386bc49ecc3ead32fcae4944aed48991937e28b2bc4177c22f701a85a6c0945c8ab16b7b62d07ea9c9dde6d80af94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e24f26696a74cc9031e033d6b0fefdbe2c86615a1aff704dfe50080248d38c818423132315c7978f1f14ad961b6ba6e765e6d87803f603648fbc74c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc285515c2a1de8eef522e7e9669bab057842302eee989baba52cdc0bfc25db1e75009855ccf668ce32c96023cf6bad69bcfee3a0f2c7962765319da5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a8e8b05e2f292b2a63a0a54ea628882eaa9cce965fe41ca62fa0f9ce7598dbec7c7e593fbba3a97eb1d39114457817d49bf39f78571a46bc8750cefb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa9f31662d7c520c02c1eff3c671dc17bfb74efb16545b0a52ea1de2cc739569bcbcf7f0aaa2be2356ada60049cde72e3c5e76e8828ae20b3c9af60b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd7baa56c64e8256550d8ac684da96e5c512c712ada291e71506371df4f2754a3f8756d9061c4738c4c8edfc3db245da2ad505beb7c9754a8cd5b3ce3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33d5af16243375d0af5024b7375ee83add57b83b91f5b12b6f7fbc3997a7e9052f3eabac4593be8ba49bff5a3f67e77db352ec53d515581f398681e04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2899a57ea568b755389c5ce19a8618f893ea4d0c9a779dc5b12a82ce893a3baf16ba6f8148b91b21c4c14cb3decf9ba9d2e67a0cceab3a224557198e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fa1a61dd554e716521adb554b25223b56d260f7d39bf1e9172c1bafc7e1ee778119b73124c867ba34f0a330b670f2a7a76736f0351362faafad41760;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3821583aab9da86d9d6931564000db1644d33c106bb35970eb429be0242c3d5f1d8c9c2a1bfa0fb9314ce12ece6cf088cfb44574ce9f9c4585e2f3b5b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab2661df65304a471e47965927bca40612ccbbf7fd295e7af0f1e8112191d7e1ed35bd27c6a2ead02585cfcf6b2841f12dcdb6dd10b121880e37de33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59c78fcbb147295ad12dcf9c8c2b5e979e8c683c4c81e8845b3e0bebc2f76f82d5475276a9651d28c9719328d193b65b9f4f79f2644a6ca67b93336f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5bbc62879c3efbf40758eb70fd1dfb453232703489edeaf4dc53fc891f71333b662f8903e92b4ed424356293cc16875b022678ab9f73653b3e05f2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h878d4699f0f187793e2095d7993fdd740a91c4bfa44643f7ef901f4226c3924a2b2afede0fa6d358f0a3cf930c94d6e51bb841df2d4ad7bce40d82440;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6836dff3a0609c18d153317dfab1854ac84fab2015bbcd5439544761a742c156fe8a531470939d49cc08efa0910c4a0ef213118a4514f18d185f4221;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61e6cdfb87f12a9732ab8ff5a929b44ff7daa8f7cb02a13c00f7f937ef5ae58ca6246e68b614264cbaef057611a27a1c5afb287046bf61f437211a117;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5a966f45ec71b9ebcc68138ffa0badd3c73cd700626612ebd7eca1401b27153e9a6b13d76ad7d6e1adc99e14dedd745ba38d1446d012218aa9246280;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d24f0a18a237daedb84783b5b08ba9158e03f0451158093e4140feec0be78e9e1b224963931a613b5dab47c111c754cec7a5b886519f16c6abea4f4a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8ef10103d2ee46909fc5b869efd570c1ffff629f9479c1ddedefa848a7c2d9565c55d3298a23ac80a507aca1f5caa3b60fc20b36fd583b5f5e9cb856;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fe4d3ddbdfd2221361e4518c52f7d450cf0753eba25b1f82c13556b3fe0f5ea390b8c403989b02b484d647daf3ec98fba3cca21b50f768ee1a8dfe46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19e134ab31e93a6a704079aafcd5c1a7fb535b539ee4fb96d05a910ad2f8772c4539c752d0b2c50677440693ca63f178d4bd70738de6a9bbf4d31c02f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e40e3475ed19eaf05b14326567d9f7150f64879e14aea07a91aa36aabade47a9675d7bf581dff832a17354d344acfb27e2024cbcebd95051b96c987a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3560d32d97d7d24dcefaf2cd10198789739f54e5e88d9a97830ff68aebfe9b70ed995b2d182b0b97382c090192f161b7911f35a58bd43ebcc7f748f1a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdcc4a70d16f7261477deff5c927b14678296dd05536908ee637928d074113e6e823785eff6dcbf80454afee64825767e91ef5c1f0dcdf2576448f82d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ee93b841213655d45293f014ad47296297ba030bad63220dac532ccdc4f06d408a01ea46ada4dad12c03b0385a6873c72dcde373c84e1557e71f21bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdeb38adf51de1ce7540ffe59b889c4d6aecdad0e918520c76fc84ec07bab7cfd4ca01bcd325f5a3f4c39fd7029657ed6348852eb4e6aa4826059b292b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10df041228b27219efb5f45a3d048e1b1abd073a4309daf79f55ee1820274d223a43f8ef80247747b3144c6f36ab762bec53433c6949cf01de5759d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h372890f82828d7f2a521e7d647372ddc7b8a86889bc5b1e215476b19af4f4e8710346706f645cbd377bc9507ecf8a0d0605e3896fbd9770d1a2eab3ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4485fb4c8b90c5ffb5426be7c0ac0eecb571fd4b8d73155790809b38378bca85e67b8cdcfe2dd07a7d0a5de5c10a1051d38e832f784cdb95b2bdddee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b4b20c63aae718803f26a6edea259c88f15e0b018f7eb0918902bc664449b20159aa50f08174e5af145103f243bdd787bd2d8ee75ef9b63aa4ea5bdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c114c09075f21081ec5c9f72aa52a7b04daf9212b4740c8f5a943cc719d0e5a8231d3133878cfa536f6388ee9a003b21adce2a3fa50893640310c7a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b994269f01e5b97d3cde06a3e7411787ab037b8bdaf5318259d5b221166ef634f8c4789574e1a3aaff82346a78167a68bb2c111b739e0da8b007877c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9cc6b15c2b11ba7603bfe05fc12d5032aa9b71467f1f968edf40fdefd149c4d896185986f4d5e71a4c0b764f31b62404053c0202f2c0d693c3d1fc17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5388fd0d886656deaeafa30bb00b5fa49f462fefd9978c39c527ae84de7105d42f4efe00a4d9513e41a83fa262cd3f305d28d595f838231318201a002;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa1d81509f6f802a3adc45d34aff5f9ca6cd28705970d98832a1a1e1afafefc7fa77f1f799a9186132ac4a9b795236148c2c2df8093fd46c4e44c6fbd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bbf20e675a5db89dfd72942bbe3c025b57af070430c6855ce7f8e77942e298a69ecf5facee2b6ac42a8001e593650f81df2f6db4ba657093288e46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52f990a2e7b94bfaf7b862b498b9eceacc97da87d0b24151b14a68bc77c52fe8995b84d06ab857b1e4c45cc397be80ec74bf2b009afd8c3d5178577d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacbdd8285869d8769ea32ff5986c46d24a21fdab1259a0277e99b90f1eaf9290150daa9ce05f0db5d76a686a023ad5120e4dd86beafd42c6ac178edd4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90e53486952903f1cf77cfd25f3cf6e3954513a4a938779230f462ff587019804942ae7b33881be7d30c73de6b23fd608a91cb525af3ac1d42c0e62a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf804157d6b2cb278038f260055b853293592be712514bc1a6decc84a10917256b81273803f7708fb03b81f29b160d1b2e67d80267b4669f971495b6d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11e01a25814af594bdddb33845e5581dda33f365b597f73ccb93b707bdcb344bdcd4ce1d88371f77ce1b256036f2c3bdcf8f8403ed0671f0392761d3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h989303125736bc4866a92219ee2d75593f78bd35d9a2ca8b84fa6b89df0a4c499d3b4887ded2858653dd30ecf8e498ac25728de6bdb44634ff3dcfad5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36e948dff299168ed9d1685c42b37414462e6b8e5c8bcd0a4151cf9e93a97668d4ad39b0db4eeb70d099a9f275e8e5b70716756d3540d26937ae18bbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81af80bf162f7ee4382c0df1a8eb5a82db32ae52e23d5d067e1f8237b0fde62554d2b91cb397bcfcebf0858846c88aa8de70172c65b23368cc435c98a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7d97ee992739275ce238bebf58b9e3ed4376b773a0e1558cdd1d1a6883358ecf6bf6d0e8f3cf748229e44691285bac7f1203792db0340833c85142e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h760598dbd61788f10292ef7f6e0ccfb6b8fb482161324ce1e67eea1c1b5dd838ba759ba3240bc86e531289c91c375a74984ee7304cf69bebfb4729fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5faec3f65050fd5c3e80a930ba9fce13ed15d94a268f7f8e86fa64e9431989c8b3e641de2bf0b5c61651afeddd1305e0e2209111acfbe40ad68ba2b37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8ff0a0446c5b24d88c0b8de32b8ed8bec485f78792537b6104561868bc7a25dc09a53e6294f214e56c74c61cdd087ef1718a138ae879cf8cdb93d981;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1152c4aa00091c000f0e41925716dc1230e34f47e9346bbb6dc60ee13dcac4192c7adc655bc7373b41d93b66c3a89339a3d53fdd2b190bd3eecc3a58a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb03391d6dd095fccdd283f281f8cf1874ba989b266e15a1139d3b79173bf7867db30369e36f804c54e917469884f020e6c533f8e26cf3be4d0a740d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f05b745fd78f59c9488f32ac25df0e0bf0358fcfd4067173ed871a92136b575e873d22260c2516ebf79a7087049dbcb25f65c4242ef9e7787804c51e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hded00d2ad723561472c3266c2ee57e84bcd6374f378de07d438b202d2c4f5d5a172d8185030af95a9a2d51688c06c726f9e7e5d98bc1bab8c9b143219;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h225350cb238f498515c243fdca55a21a601f53591543b06ae095344baad3e6d3a65404e5d23ebc6370d23d105902898cb8cef5c991c1a1b50f2bca77a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c4dbfb76845d5062ba6e15dd67018215dd2638a67458b10db6f3e3882304327324071b6a55b7c93a36ac9f8de7dc4b56830007839126da1dec9bc670;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1305efe33d83092c214023f92e6e2f2fb87da942ac997372a5dd4a415b6864048e3136339c0d4a36ffc748392cbe3dc9d9bce969c60009b75a10b4c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h934bfcdef5a68202c12b8b5a50e473d90fb043635fa477fba33f21ea14f5f99f049bcc0f11ed69268679ad81caee929d3f731f5aea4b40010760a0bb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37607f93147eae5ebdb77b357cf0b6d6c42835c9d44ae7f6ab1b93d826a6643a30d18257fd8a3e1a2e40e673477767b066d5d17cf9d2168f1f746f1a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c8b03207993369db51ab2159c84914ec025b8e3a9c86eb5a6692094a7d628ed262cba3a599a49a129bde9bb11402684b7298f0cbdb70117fcb603225;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a75f89d9c4cf8d4e64ea152b7e8dd1fddd4fcf1d92cee9786717a51861599c7813ea038b3475671bd499a3ba262a12f360ac3728c595fd9f0426d55e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8f14be4412e921f8218628d51a03b94f3bc71b21cb24f3408af07c5b1ff539179674286cd01f41c2ddf090b76e78445e2ff7fab51ad7c063be73a75d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9bb1040673bce3603a98d41fe733b13781b8e8a2be61d439f7cb64c523b612e07e62794eb9291804cc1cba2efd1a666e9443fd7621f3d8fb49866193;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b3c4fd404e09d495838a66837131a7812b8d4e295c6b02efe89ab1b7e20f6e435380f6780403ea064c9119c338b8f702c413bd5eb69be3f6106bde7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5e7bf457f0b7185b8a282d4949037c15e7b1953953d514a9e9689898be86613770046320f66d887a334351208186762fb061900a4eec482d23543a7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cce0fa08168bd52582812118a1e2488b2bf000df0ad4fd040485d397ac370b2b50a5f2d7c06c70a333f725c8ac1b12a9526513456fe1b8a55dccba1a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf1b169ef6b6a393a5f9bb69c40cdf75104d88cfb05bc3b06976d2337c6249bb21eea6104e8789f50f74288f95b82adf3ed5eef10f0c20ea9599a285c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h472016855842a7653a3bfd8c0a4f16a61c5e18b9214f547c430d0e86c625f8eba12af6f9fb6de6d49aa24432f1f7d2f0c3c5c473604c3ba9e922e0a46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6524a5cfe07730245cb73e2783f2ccf1bddfe09b8eb4584aeb371c9b4aec8cdc450243ba835520fe2800c488fbcace55f6d8d5d8b0e98abf916f41d62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ff5b8e6744947a5b337501b92188d16750c9155a6341acec978328d724feead817ea6cc7db30b2400d6a8dcfbf9722ec83137a207bb9c20ed0aadcc8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72caf3d06baa959cc81c750a5fd33e35b8d1997214043cc9dc73e17d96331af47d593fbacfa8916b65411acb9a24993737a4ddfeffe36658f4ab21ace;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6100539f72da5c67b83edcee9529c27026574cdcf2a797da8b345f109c63c9e8761db3fa3292886264895bc2c5285c357850a5f1085442d857405f7e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac7aeb5c27283bcffdcad2188f86d6e6a3dbf9df530e3cdff4babb168c53ac1774a791c2d23694c109bedd6bbf8ad0bc656f1f09ec6bf4f29a849e40c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8097c95ce1ec51f4d0313b20a0a496169d14adc693f99d30d0e7303929ca409a51fd08907525d215f3720c0f1f507e439d0dae8b1485f1983ac0feb9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafbd75a6aa02ee4be88a54aa95465f3856b488270c1d33b3254006c5cf7e7a56d18c2bba0603bb10f26ce70089a1034a09c15633677f8a6c3be6f8560;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3a404d1baf4a2634c2d1e787f5059e2236451213f1c8702633ba78060f0330673a705de71899cc379a48bc918fcd24066f2094cd65752549b391615d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2af9b6fb61198bc6cf733030060252e8ed7e1d11026abac56bdf238dd19bef3872db2978ed9314872e5cf2ad1813ce958d480623e5d76a8785e1d7c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7555c8593c32b0bb4c2cfad566ae93265e94c2b3f9eb91afbb6198a94819dc9906e45d5779811efeb64d32cc93187b0eb6df35443b10fa353e066a93f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3dd0da2fc8a3139ac95280981eb996553624ef620a34ae2631e52791125340879971c073a14632bf7778cae12c3aa17bcfb766290e0ff211b2002e40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18afdea7c35a794e299bab9e186c02077e0544efb3bb78b0013b44747c69fe558ee406e6021f6074a77b93d644a81de65b3f97477996d0441a6b1b9fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha40532ac1037b99caee351aa61c7d8e5975a59f1089352ffb355faae799ada49acb335c2f25794d8688e8a2cdd6043fcced7de3964093e2c78393ddb9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2af5a41ae9a54f6ca318c171bf85c5a4a8e1934dc3d5cf33774085e2145983f4ceea254f39d0996d45e9937c4398b1b2dc6bd220379534f6f2b71d506;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9b1831cb952ea1f34635624c45badedca565a5cca2f9f18d913dcd14243bc207bda6bbf4c34c6b0e8cbed8482b6bb78e01fe16d740b0470b28836fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90aa2e57bda5dbacfcecbcaf9e94b4e86fdcc041aedc332ff6398e196bb9e5763e7eca674e7e6cc0a4201738cb5162433046a1a7843f632c2ac08b848;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa05f1ea37562d72bc5a874427f0e0dbe6cc1a6d3a14436e6da321ffa48e0d49531e03f9e1d3f493d3c15f2cba9f3042feea5a13d925342bec3eeaf6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c6d8252c5ed83df6d418fc1589d02d936bd11fe74fc3ea3bb387ab7e99cf41fe9dcbbd9a5b9e8a7b4ff5032fc7e3ffe5503c76fec696bf1dc7f9d809;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bba17cc64fe8d18f33523a424442b0307cb2416777353d168c1e48cd40dcee426cab2dee82ddbb2d8c5209e4ee8791b006cd25c5374f5a175ac4deba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h233fb2006081b3eab813e48f3161506d0a9589eb2bddf9f52487648a4555fb3ad25fbda18ac36c3938db050cf94d76798f341e724003dd1882a0c3600;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48198ba9aca9c983b801bc6eb440c917b92fd091602cbc5ee13f5786bcca4992cbd18fbefce9d1eb252703a2e128b0bea5dcaee58d5a8a6765c687432;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70c9728b6b636a074dfa9153f930222e66de344a19f488ce2cddabd27d6c21ec360ae2b2de6c573b66e2613323559dc4cd7615a53be49bbd1b795809f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1f4318a9259f8ded8dff6793a4d17f50081bc407307fb74f69dca211e43d4731fde6a32e406b6fd53e59b2b6717ade89ee7cf524008de168869319f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff637fafd631101a1ee447bbe0c58d5ff2f254cba49aec39a0a0e1cc48818ba4824efb24a06fab0041a8eda1085d75e9e4b02db04da703f22b2b40b4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1c21e0c0e30553cac8d43738f438f31a530d021f0c5f68f49f14b51226abaa319576aca9ff9a7d754ee9ed2128817da5278cfdcc65aec8c2cc982170;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cc42881e659932bc07b2a62f3b3c9588fc1e655305572329e4bc56c98e73d32850d7bf909637088fd0a509accfb5ef5540649d7fc4b6eda5279527c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7febb9b965f2850d706cd3e1026b469847ee3377e650a8e507b2d3217c0cdc9b4d54b337873ca6a14551e1acc878b8388f940dc4b90259970aa70e55e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4a155cffedcc89281f9b787d9315397e796e709648e790ba9cb18d7eda98be53de51dbc43f187789d6f3ff2c6bb26a0793a821729e5e52f9ed573d89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f7dee78b0c65d4ea6d5239eeea0f99ce6697a7f5ecd72006962884d61b15b1a622830482cf9d269475d11f5b873b044695bb4577af2f349b8948b9e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb870a62c31928e9773530ebf3a28b14319c165e55d1ae771198ff3fc0ca821398656311536feb962c4ecb9afb699faa8235a21b28e36726d52d5b42f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdc98fcb6e63bbc44cc7c9bda93a369cddbd56d8258ccd69a1695f6010585cf7baa4cb04dbad72e2b89832242402bf50fe27c1b651a02d4762c65279;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dfb3f5d474d6a1205ce10c030f9fd0c231e58fa5d2a1074209c0b79f54534412e4cca78228b7c167dfb23b2aa07ea8f5ab4cf1b97f8571fef91e8c25;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h513cda67a7b9e4e2fae6a8a924d96f33a3f572993465d6f8a959cf86e6582c3ed8e2c468f4ba4e86c17688578e102debf1277cb52c975bd824a375ed6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15d2903215b936b993557fd051da431a3287b75c0e7bc22f78035c808aec8e3c67ad19fce96d9a6d7fe0e107b7b84c0457bc1418d54d3e1c95299d8d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59c3da7837bb1d766c1a735725ce12ca2b3a0fcfdd64875291307e91ffb2b81974c6a46b1823b06c0dbe66ee2af73319d95c45dbc1ef482f767f10e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h706e46533b6674fc1a8ffff0b55486d5a6e1d85ac177022ce81967b210a381d8a8737e3aaccadf95399a3dccf61897499060c75e7ceeaf3240924385e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ea1523197d6186f1b45529f44b891b483ae7e328e34933da01ca02c6aeddae70343042f816fabdc817939fc1295e6f0a22d06f5956b39a3ad66f53f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb012c9e440062f67c35110ca6dd8c9bd78650390252cbdfff163b3a4249e7d397a16c86c0c6c97e9f4b5460a4c178319c8354597863b6f2b69d7eb27d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1709f97a73bf1c503fb6d24def3835a0d5ab99fa7f8d7817b758b0901c255a785ffb0304f5d380e591bdd2901b876a1495772ec2a8610d892f1433c9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ce4520fdb5d5b6598bb1885a85aab84edab514adb433a9143d6c2af643439c4d23747579b900139c945efa6a3ae9afcbf06e2d4a1beea178d6395e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d50e06c4ae7a725890fe38b59b0957f44bbae218837ff7d9af451bc84fa0d2247136836f3cc3e3187b861a1ab07c9af4fc0d5ea9e17d2cd405d410bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3a6a66f4e7846fd93a0c00d05400223f49a094d9ae70900c9de3bf1a786ad03a4b638065cfe39e2346246d9cd0e696f2364fc0635face1c6b92f9ed0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12cee54dae18876e7d63a9bb22dbaff7be7fa876eff67a81f61c1b60a7ddb05349fe81775e80ed245d839d5bed86a25ee46ceeb559c208405ec72bff9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbefb9d8df9761a291c9a7c27d35f9dbc375ae3d2bd35ddac44274b5f8994c18228047ff775ee19b632c6427757a7b6ce49971dc138df1dbcf1700e947;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f96e4cfe7d1936b4a025c245528280ff76abb247dfc347b155d921eaeba154c3391dd7c4249e2d5b804075983b2f15c8cafc0bceae35dc7c97d2f10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f8c0d013dfba3ce072c6b45e4ce5a39aee33c408408a9969d5f5bea0ab2e1e0458fe721407a9d79e2335ad80dac711044b32df730738f58b61fe8249;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h671c63f54e01cbbb840366d22d757d918410da673fcf5b6462152c6bfe047e1b3e5549ada5ac4ecb1b067d6b6efccc5dad7fb7a0b8e75519cf5d0f1f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c568614e20b73732898294ab420bff58da13ac11f26f2071165c9322ae0434164935c76f63f5beee7a7a5993822eb9d682243aa0c14d458cb7402cfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ecf5708449a0db62e7da2bbb959fe989c4f8d1b49b93b170e9dec76af085272d3a9093c050590463a9c1c2897f95fad07d663772befdf4727a042d73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa98156a8d16692107ac2f62742cff628ef80f352826190ee8593a553610d645562f5490ef05e6a9c09f7d47266220a0e2d6f14afa80c36e7d8e18314;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8eb5b60ffc240384138bdde613a5b575b580baea9b1b3e3b6d4dd1bf9b82a7bccd3f145567bd38499e87c050b441602673dae10403a70df7ebbed184;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8df28f4435ae0932fa38199cdfb0ced9f205985983aaa089115b78c952fafc1b70f06c9e2dad0b21475c128f13621398e663265f1cd6ba65a30a88e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e281a6abd2195824b4cb319c9ef81e875dda06cf160287f48166c73e306c7db84a0a04ab01450c3ff6b784af6f3777786f7114cdcf571f61cbab2568;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h248a1847048ed6df4b83aedae12151253185d54d73fd13b8f8361b8955dd0fc0a922967b9c17e5b20f7a59fc92b8e939585301f34b060f6a2347a102;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc9619efe17c5fa9b7d86c949592d8a78fb7e7774800ce70f016c0ba5f13ce7fd9c68ea9e4189113c9b40fae6f01e683a1be5ec32910e8b659c3c22e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5e3de570fb027df69377a9b7eccf1165a159daa1dd0b07d7b319ce7967125576cf7191d69b785be3f83ec5a3bec463bb4799c402957a069c23ab30ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8f3d39ea428966a7094c43d9a0eef63d52519b9b16470c9e2f0a9b692a8e66e3336c195411ea421f780b8b4603127cbace202388e48a92ad32c53a9f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77f58138616290b1ded9c3f7498f366c657c8330fe1b00e399fd6c799860ad8a2f082fa9d82bcdd4813dde5dadf3adacc6c05b94dd1a09f38c89a039f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d86f7fa2ba9b09cafe1b4ff1df0b1104c5ed919360a0292e7cd85fc7e0e60ae9ee24f6c3861598c3a8fe9e863e9a0f31e66f1501979f638cc01d6564;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h758ce79ff1ea6340b80f1866d5bfde8c9eb8fbb452c670d684087a07fe4424a8bb809d9eb5d6f14b333df27c84beb4a1f8046eeddaf885376972d36e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf556af058a3f49b7c287e681c39827cbbcb37545f10677d6f169ce97d7c8d076a92a4ae8eecdc98b3e6caa1f23ac6d8fd019afcaf961ec90789890b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24b2046ddccd50f78581c41eb645b445edea17d8bca5089f5cb6c502a41ea609e59d5fadffa9347e21c564fd7618e374f9233ca1a39dd2593da859410;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6509b48806d889ed6e57b787423f1bd78870799348d72909f94839198c708e9e58d5e7e5e0a88cc5933c5865cd7bc098d7625270c3348072b77a9a05f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6838c1a5754a30217f3af3e7ac6edc8f363de70715aafc65930683b8155b93fb88bcbdd9e0108b761d265176f20c7b0bd6b3b7a09ab8655ac5eb57ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc187dd3a4c1e91f924e2fa3c5d941746699c72dc690e5278f7a9b9f2e33b885ad0e441e314a53f62b3a5a728fec722b8a93356e1bfb5817d2fe6d0b6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2174c7b9fc6a178dcca95f2ef96a45d3e67eaf4ddd318a94905dec3b2c92948745f440e89ac9bc54727aefafac0e38d67bd165ae0b79f9c8f930ed912;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf2cce9f51031f76cd7431cd5f82a6bc556e6d1af4a6924449387c71a9a633a62245a950b799306fd6a5ab444cd9df289705e7cbaabe250c55b904d32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h297ecf7e7ae7b03942f2bf44b16244bef47365e0847443b285ad9432ac23fa98dc1f88e6752f8a31f5cbe588a4500faecef1e111f2d181af19b003cd8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bd3432e18333a3435fa9d318627366f1693071b459fe2023130932899963319f48c2cb4e4e30a88251dab30c32d67c2273afbb44830ef2ebb7cd2e72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28f5872cfc833bb78c0f80cae138a5998c8a250de07958657444dbe043a6b5e49164b1ed5c5c62883a248dca947fc8c736aedec4bcfcb06f24e5fe67e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb90f4a41ae749f9c03b3250f6bd7deb32b9b35a18c0f1c3df9227b57d0c70f815eadc7c66511b44c1133992150f3c06e4b5672c220d68ae41064e4fbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbef7b8eff9292f291280c4e6494230468888e9616c57852ff99e00b43b25ec31dc44354878227c9e3fad0c7c8239106be53e627bfa5c7ae8d679eced5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17660d241198e92ff74a5475eff7f99dc947b6a395f4543436c7ca445d1492042daeb7c5932acd9535ba6eaa5f6cd555353d8b365e28d323ed86c814;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93810d6e3e92b95f0451e4de08f1e36ac2b0ec0e6c92d229c6a01e7e2bf2064d901a14be38805c3e5225e16014fdef71e6f041a9c4725a023000d6ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1732375f9fb8c3addf2689b51ba7e8ae49b2d3189db9945cc87c6fc0a2cd2559aef41f0f6daa1deb4a7f83dcb31073814b39628f282c71d8fe8d1d58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbac60c54c29d1e5533ddac49793f8d5336017c8f34d07f9a38b7ed7cd760b1b4474feb0fd863e15e3b5871267b81728a46b90558470444af8dc17f08f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ec639fa1c01bf80ba7363737555d838a01a78a7ccd25aefc6ced41a697cc6870e742eaee1ae374076293cf6a2bfa36a1a1e84203b3cb2ffaffaae6b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91b2a8474aa02e2cdccaef3fb90d906c2b0a0c3ff776f3ec97b925ad1fca561640fe1644652e72b9ed9254b97223bdd6c3384ebf8e6248dc19fb8efd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57efb28ec64d6f621a1a0de0ca7f72d543a36b0dd1b40512b9a7378f39a795dc6d38d8b2380a83e72a25f64a81d012a97a3f73f6a9a54d83d0d8dbb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf529b8676de07e15b992caa6ce7057e413863d8b48d025f21488f4a2b9ff89f1f23517a87ddadee0368be498b8e84f55c792064726495f0ccd20aa727;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7513d2a3a2146e2263ff515ea58e49e0192cb063816700987344c638a1359a1bc7f72b6bd283df6cd9a1e34fa06cc6f6949d609c082762cccd18dc01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71af9f9d28f429fcc69572640aa59c7b4391b9e91e2f7953803ee3d0f41f5c9004167a2f6a553c3e3e2ccb9ebdd83e2da6824d01d63f69dd4f9fbce71;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c81f9dc77cf126f6b7788652cbea7b8c3e31533c500188a8681795538465f8b749ff999c5a820edd245e31d318cd09e2690fa0f4bcc4833f364c6609;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf88a9064c8fc74d72fb65c4b6a6f4f8e126cc97b7ea03ad262b3103db64b444cc3e62d303a0b66cb2d7963ba34e8a51185012018435c0bcd0d352f1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha80721b7a189c89f82431f5b34daa22ada697a452695feb85def185044c2c239e2936ec093ce0401836d02e4881ba7c8164a5fb058fd822faeb2646f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h299779f7b914ea6adfe3c2007641270bf651f657c60110d6e46f89359ae648245ae46791f904eb3352b7900a49080cfba2cd8e852e84836e1dce387be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85f4e7cc1dfff12322d29ec8fc9a8d643c2ebff1d0f578a49817dda06fd46bddd17e0fdde9f08038877fd3f8e016b386ced663cc869cfebecab55338;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f5621ceaa513e6f88a6c90502b7775f8dce96bc3c4a5cf845ad853bfc2df980ef1ac0521112d93473a7182ad6b2762579c87e60830d653fe2d7b7c3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52ea70fd3daae8b909e5ca36dab5890eef8c9fecae7881b9f53ea893aaaba9e7ef15570fad3d3ead2857da3109381fcdb4ecf26dfa86542a15d0b2141;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37ee0112b7705bfd8b3164c706eee28dd07d5ed6d9ece7e7f0e93b76d76e74289b8ef8feaea26490a2a90d5e75a6f851b2610b6e9132b53118b3e6f98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b6554be6a43dc803aa611000472753f6fcd4a14a32166d8656bba3a926b74f8f2c361cd6855f66a1d5edc7d5b49accfa83ccb893367f9150d2bec5bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8af6a34d1211d8f47bf0caab4a2dda88d19c6d821b043701f76bb56c50ff9c8e2afa7aaab39ece27ae703584aa2bdc0d495e094b6f2d6daae198201e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73861599c21cc428a9d4f3a11da49cc46b014fe76a793237739efaf418485c2bade83ae916b30c75e955a06429d47ad8267ba6bd0670ff6bbbb5032af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e474999960838ce9d7b1c2da1ca7c882cef82f52404108ad141202c0eab972a1b8979563e9a1af9336a20dcb69cdf3e2927d4419e12d9831be2ebdba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14b6c23e14a48c55ac9c79f0b1902ce6f2fee5018e5437cad2aca64bbf5e47c600dfe1b547fe138e21552829d1e926489d67bc354492e6415472eacc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f63129f536cebcc12913a8f76c3feb598f1dbae281c374317bf2a0e71b8fb65e8bf52ce85009eb53d8b5d286fa6065de8bfda6eec66a4816a35d4b48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb80a4ea7e372bebcc2da9355833b1c9c8691646894795d92bb9c273f417b1260d804792804641cd2081e9669d75a2aaa39ca025c983a77725ec22ad79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7829036cbac81ed40392284bfb3946ff9b34b589ff79b344052546b1008906e326446443dbd5c67da4b44df32107bddbfa9fc7a48e48620eeb2f755f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c7f67e114b3d788e39b02e3334262dedb0487d3f97fb4bc62e79d2bc34e36dae9866a8bb73b727711568fa4e7759913c3255797990b8170476c10b4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h190eb310b6521ac9153453b69b2927187a7b192b6b4739715ad23d390bea69528dbe52765f624f34c7111ca1dc94eacb5da2b5d3556e97939a7808ad5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ea17f02e7df68a5740b8b46bdad6b34ffc8372656a5aed076f550af034a45789c906b59ced0752771a64fb8032a9b290a0df1891d68de705a3f79e29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc13eaf1c5fb3c1e62245278a7ccdee1d10211b5c3fb38ac9377224179dae7440af6f94349e9da32f05efd560fec3e62ef161cf46813c91583c9f28e4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6760c036122bbf49af300e830b7cff673e4ee1575eb8eaa98ce208eabc72234c8cb56fecfc325fd721ec6a226f6dd3a587d96a11b202efd3ace98473d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f6a68967d2b286ba7f51b4510a4b8c2c3bc12313c26aba27d9b113a11682f0b0bd0e9301f17b956ffa34540c13f9ad2745dda63ef2f0a1c469e94ebf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h191dd0e81921dbf91b612a738e0de04e0501b8c9a423daa3a95c199e4659b8bb438505beef35a3ce1bbe6606fb9f56635633e98fbc84062f55063d1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4530fc1606e07102622d70660f6d84d3a93df4b09079fe2c85398a50de3579d138f2a9574d88faff23ecf9b6030afddef61148b216b665699e810bda3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e5a0a3469d8019a5275e64bab4c272a4d5a5fcef93cba8bfa8133301bcc68cf8f78e36bb43c009d065bc519d4f5e8863091e9374e49af03afa4debac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fbae4456fec5c26bfa52e2ff437a02ef7ad0270dcce279eb12ce084fb404aab5fce2cef55b3d91634bf009bf371a50d57aa9f18736b8950f9d0ba9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fcac19acbab4a87eeb65d0d27b2c67f15e9cb9f6077cd4bed8b5bd8468f03140adb6cc4fbc54ec3420d2091873e71a7a673cf9359990ff86372b4532;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1514759695741cff1fe0a53b84612ab3f307c04309d784b5392f14156fe965549a1ad054dcada68456159912db4972c8910ebc841b4b4d42cc3a66aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d41188c737e3fc8c30a6591291fa5e19c8d309a423ea387f6eb99f41fe998b4a550d51a9d736a600aea35549f7a7ed2673151136467c2322f78c3c06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf24047f9694be82163321976713660275e94874375ef75f0b1b670433642635d0316292a580e26f7af1882813f20cf9af565534b68851e232f7f1a43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5ffaf46af1fcdca46e297cf47f86d8703f37ba1f7558c8601d0abd083a3d90e94cbb910588d14bda68e2191f095bf051d6de2d13633e476587116b3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadd3ded1221bfd24283c1fa6d6c9c948483f008c0a741b74393cefc64d77bd277c282948beb27f5d099538bf4b57dcf2dd3988f2f4db09ca05657bb2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h583636f03ef33456eb467c487b27e3259b1d18bfe6270bb8958eefb116d7803cf0ed727d31e8839e77a720d095f52dbf731fc3d1ae68aa4834c4269ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he39154777c0354c9229a4fd2a19b42c09b343ff9aa965488f6eb020dae5ed47e814ae67822357db6ea69785dd64fd66cd9779fce9407744afb2677b13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9629d9897e8a6bce0ec32bfe859539b70817592dc06c15b4c13e868d489435b2c04691af84a18f079003160c6b14c4a52c6d4378c622befa0a1cde3e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b3831e025f75980c46d12da5d76547c7b117ebf3902355e7bfa37b145e017bfd87b71bcc32effff7ceb547b20f884ab872f534e4225413c61ae66e82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0051d52d47de42fdf2cc6729a309bc1d96b6fd9a419ace29b6c56c52faf5f5f6f61d47c9df11c2ae6ea8e76bd82a76d486f62d02c845ca8c88ec4a6c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c32e4fe136b81d1143481d28be462a69c028ae3c5cf7fcbf7d47779a6528d14cb7e0a6e4613e0ee63435af5c017024221d1f90121198f0933afd13fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h218df7a7a4d8d8f09ce5d67925e60a8c20e7144fd40bca8a03d413a5190d0a2bbcc3f1a3f7ce84a05e1cfb3cd7790fff8c81d2fed5e0338dc2dd09018;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he750f52db63c5281b2c674fa3795cb5a1a8c84d04e056b7bc9cfffccb8d920b0e2233f73cf2779c4edc73e44c20beebacec28c1daee826673814267db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h731e884d4c6d350147237fc1ee2ed88c434466a3061c7de410c99783c5587d49052f3fe4b070058ca5a177fda30473af20433fe91f73f84b3ab43feb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ff1d4b75862422ad0a42cfa66a5f13b22d45f6f32372e5624520f675efb8acb98de53f72529f9ef6fef6b1e4f58449dda6a55ad4a1980aa8b515470e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78b924f36de9b595197060b81477a642831d1013d3482780279014b8b7519f668c5d1c4649f39458c2b3d085c34146c6f919cdd316ac6bcb035f8a055;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d0b21b0b8b1140c48670d5aebd6e0523aa0f6a5407b0635b833f712e13a0bf270d6e85cca9c9cf5de02937aa2618b82c4720d80602e6a5feb0394fab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27addaf8a4478bcf28ef4695ca83fbec4c0205817d5dcd29ebdffc0ac42c29344a0ca44be6b21da5aecf6a89204760160f9b04723d4b28cd257105414;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd724c2ffc805a6b9c1568637da2372f4825fd04f9cd7d83ef59c9cbbf39964cb8458aeaa37679b2989fc1dc8a569f5eaee5311ee3e454c57f2ab0bbe7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20b67020546e28dbb7c90b40c8eb06435c2d9394d475fe64100dc7d687d09d3c366299332d4711e6114e52b17af95660fc56c66463bf6cb34acab7b9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb71a760083201c59d1f8ab0f579a77935fd7628f5d9ebfd311cf11c113c3316ed77c5497a50b5bd58f9bd0dff7a559b0e8ccd71f772d2e369fa7497f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a07ebd47e403736fd633e654d628b1929a4190111bf0f73ed33328d985ef5eac9eeddef5b8053a21adc9e2151a723a9e971914e3641db3bc6ebaf305;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h357e70eaf02bce7ff3f2f0efa826742781c6e0f039b0df4ae05ee0ef1740c54a3efc5465dceafba50424398243d179d53b30952f3883a44d59a27b496;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62523259daacf01aa60c0c2857442b9ee6ba00beeb82508eb9446aef7cd652ae6e10346fcbffe055eed92a3474c08c3acafc20a44214e6ccc72e1e14d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc98333288b4f7c2a0d3a6e0ff815393f82dd8b769cfde8b8ad9f9ba42ad2bff436eb6559d3d8adfe7cee6bc58b3302d2f0e8447d749ed33e07350ce0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf162387df1d33a1b0a22a34aa6a3fb84919095095bc1536e4aed09f7188a66f9353fe48cab87456545573ba796ba68dc2a38b79756a30d82cf9afa0e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2bf2320507396c89f943f89fa4f9e9a4ef089db60de513a25a9ef38d41307bc5a349ddf6f130c6e39f760179844816109e29aa313fb61254259966b7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha982fd04a507d12fea9a4f7b5f99b21c3f1fe806100be476312acd11f90dc38964c9f393df6c6473063ba8c6699c70fc397c3a7dbb7c7f8c14f7b783;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac4451e258ac1e4507ac5e277cdacbb2a1d0544b9c9c625776a6b83fce7ce57e8956f6d1624a7b06bc7f503e3fd8734b1f7bb830f6e020c423ed0a193;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bf1fd3701bde92b9147b724388b91a7b467704a81d5c51958c27a9ac80ab5a8285452a0352e1cbdf8b5e978bc9f036714fabe98ed8b7278f13f93c42;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdaaaf5ccb3c435eb693a647aaf9c3e827d6c326956cc840af87470f9cf10101fd7dd14f91e4b96379b1d8b9d529a7b96643d339cb9805386f5f80ed7f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76187c92d4ea8fbfbbce6a82cc941a98811f189a7669c325c4039471099cc991aac05e03d9bdf253c55672a281d6fac53fb97c05cbeeb12d8d7edeb4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5186b169764e2647b47370b5ca0d0d6d8adc0a58af8cd9ceb8e4cd92d75f64162d1de7cfad0dea018f2567b3537156619a0f246c4cc32ad5b2b3fb197;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd663245a9cca7de3e17f3a6b21c306709d1aacc87f58e3020f8ccd8ac135f3e0b90d130fef125e74e86492783c9053bfab9b438f60beb6d25e95c09b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd687ab618770b84d347c9ad435e34a6f29a3e9728ac674cfa18a15049dd47eda1858588269b7f2ea8c6e4b17498b8b4e580d08dad81e65f0583a04715;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa9f56f6320642f50caa787390f7d05fbff5432515f7ffe943bbfc97913650d9c3e87d023e13e69ab8f1fe3983d86727e213645371d3f3f65a82cb385;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h886218e7eb398914616e2bf8986d58c60bc43ea38c88439622c0ec75fc88abbc872ce877d81d0391e8585664e699307afad949c9b21df138abb37e5a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb8a66edc432cb020e1e494045167a3ccc87c92127b12045972803d3aa57f3f2a040439f63ffa3795d1f4345fffd4d21708b27b5b0ad660e6d647d20e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35ce1178aa70add7f6f89d24b5f70edf5b86b107fedbf305114933916cb87901a23238fd0216fbd1abf5ddaf9be84d31424350ba7b2ee0a1ba886d8da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h999d100c0b925f93e1442f1c1a653102c3eebaad06fcc65dadce9708e6e77eecbca57793ec3134e57eb74945ee77d1e1359274f7920b299e9f3b88a7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha51ff504dd5f976a4650de03b9ad84abd30017b599eb0f39fe918fc25b10e31e0f32e76bcae5b993841c47b01d5e510301617d5cab00c5fbfd3ad9f81;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c8c80ba1592289406a22b8146b78128ee5528001d4cd5f76b716118b5510397662ad1af02e9973149f7e9f085a27325105a530d92926cb7d1e3626d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9937535b80a3a78ccc4adca3fe0a326ecb777b1217c3ab80064cf1925aae2013f2cb873ceead53a0b58e4eb55c2b81f69fde61f52fd3047f21b78e71d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5126428a4ec1682a2b2d237f513db37a73d6b7346ad8e007dfceead847e95df2c34f0eb61c73be0c523440f4e6450adc759cb551683518167679290e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4de9693b3aecbb0a5a463c272a4cb0a1fc58219350cb0aeebd115fe894679e5a6c80f83d185a215c24d93543ed04eb027265f0cf781e34c51d3a1466f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b03bee695b486ef40b703fe9f01c240c496b7856dbb50e16d2ca09e60a6eb0b5e1f0994e78e465d1ecd014138c66f8951e98b64a86a31d06f679a793;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef1dca56eb98acfc4af5178c1aaf951483e92745756ee289b8458738a58cf32c05b54b7ade869898d6716972a15b246517e50abc2ac4fe27a60f6c069;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1f0e5b8425be3ca25fb48b59ea42c3ac0e8189a92b25a96c463741ed71f9a39edaee6737e9d734efdf2c02a07a146f012bccee7be91ad6f084198cad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed75b9a43c97914d05f8f6b41a8dea2f08aa3d1b7be9be671c0b1f65840bc635fe1e893b18bd19ee8d12903c2e2bd1641871fd96b50b1b26df7995fbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf1c0c2b70d2288af2d2251f3a5ee7a9bf3176bc3dab2975774298882849058d783e38a452ed3c714b4b8adce811650f523daa3a27e6458adc000f269;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6931ebf65ab0ac8293ab0d0ac977fca52da189857c1e803d3913151bf2ebd88d0c47b982c10ac140c3bc0b6b96e51e9de70a101606873f8053e5280a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f82310db5e1476fb5d6e9947cd894b31087d82287929daca5ca04baaa2216545ff76eb33f0de90d213402f373b4d94e4715e8ea4fa84e11076a5ea74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cccef28a8999ae6a2e68f54da81a92668235faee6bd8497c914eff119887fca0b3548c454e6abefe91b0c94d33ad21a684ef94311ce9a7d33d9c9c00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h498936dad74e0df6de094456d299e7e31eaee72edfde20c2dd2de1b54745f7df754f1a4bc27fac07f31dfc172c24cde763d7660cb70e8034e039f4983;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2f45fe9778ea6d188da7d9f57772fee97d0fdcb71757186e3df8c328cf65bb4b71b673dd84f11fb4a0bf167af4448bf4cb6cf0a6fe08c66471d7a83e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92fcf0a72cab13ddae05dc5a61dd05b9d152ab108b6d6182f89dcb063b8f73fba9b16bd7ab2b87259f48c6295df025c67b2e98ba85c0072f8ebbaaa40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h847b073257c47a0c689c0f5ffa2498dfac94a9da6b240e74592b308e9bf17b5451dc78a2f89f8df58f137f3d092c8c5997c03eccdc63106af7cd8fb61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had0fb8d1b667135726731aa5271e13927bb2ce31bce4794445f51a667ec5857214e4a4418c76324a79f8352b179e58ffa004c139097c4a8d78e7fa2e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cb639fb3a89b8218f2de636fb5f8f9c54cffbbddca44ada444e18bc9eebbc591c053a8f3cbabd34c25966e5ab86535626c13b43b630240db9f37e7a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd216dcbb99fafb5224955bf956f5f5c6da4136186125c9cec13f04824e5d8fcf0ca3ad8fb69112ac90e18ea28e5d2deb97051a3aa0673d395a925a76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h980aa83268eb244f05617fd5f9f6118609d053b3afffd1f184402acfc2f02d9a556460e571218e76ee9704ef887d2bfb4ac4524b16f4ebf181b3ba36c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd43ee05b3208d26c8c7e6cc57113d60ef9deadce9beea1e909ca7862e56f73ee47da5a4283382e6e8da86bf859a71247da2d4810fec54cf7de749ac7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13e46ead87f5a2c50ae7acda62ff951e889e681150762aafd80517a0527a44a5452be6912da2641e4ac14c4a6436b300643280bc454b9ff9b76ae14eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he089b61009eb1960e386703400563a1825fff6a84d98a8acbd389f37a5becbc5809d4c0e3cdbfba2b0ff8d411ad01fc434b47183830225e59b696f02e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e8acaa6729eae22ff7739c66fc0ce7315c9f40e7d957426cf02cd504bbe0a1afe119d25917703f00f3afae4adc4d7fea6b20127ce834eeda5dc449c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb75ad2bffcbdb2fffc77c25edb3b048ba8b099ab31741506b32215985a95f3ac4c01b54cdcba17b40695de7241c500dd50f78dcff65f9942d06607e6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h554a14aa6ea380523561323f83ea469ecc8508a1aa41f8b47bd038b4072baa7330c7015a8d56581f8e7ec9f26d77b729cf0f6fd9a812308dcbc31cad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25143f58f2a968b45029d09bdd7b8539009a284a77c2bdbef6b6bc77aa68d56d2b3a85288ac0b0e3849b327cc0f5c62e20177c81496b5faf089784cd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1d7342b70464717ca2117045737841e122032d04d6f5eaa5afd5496aac1257516f0a2a196b6527912b804b4ec23132f7de216e9498552d4abaeeeaf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ecca69739dc6e9f9ccc627d9662ab09e65a60e32bf790d056c90d52fec9692c223136b5bdb025b78463c8a5910846257384a804403763ca72aaf2ecc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbf728c258f05564ad93f0c509fdbaf603f6a8276dcb2b867bdd901929e819f0a90619a75153f8a0f339b293233395a020bb82239ed98c08a3612b1ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cb49c3f7eb45c8e3b1f723a94c8efa8a254d8d14037179a6dfcb45141ec2edc42ae0e840cd934cb5f73fc2f5a3d425ec2fd60b9014105acab090a904;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1208e9ef367c666ebc453e7beef008ccb8fb5cde56ad8b1252887665ee9e632f83f1a56ba93c198f1842bf1e57a826ef91610b70c940be14582c29f83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef46152647b2cfa8d400bc03410a3f1e704f82415d1a68deed1a3dfbe835f3842493ed73a36680705dc1c80df36a120ba5c9c1b15b4772a0cdf24bcdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b340fa66c2b5890a7ad650085eabc5dfc2f2b9c3a2e94c9dba70a4780904111223c247ac87464048fade2dbee952895c7b27560964fcb30ffc0bb18a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h341c77eedc7255564d6edcfe61645af453319290814953cce974707b03255fdd20f6b14c8b1395a43fd99a423a730bf219372102136e0142d5823631e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefce2a4ce622e90944140f2ecb953893319bde14e101b1792a36f79eaca53529ccdd284cda7c57b5fba476cc55f9336b24c0fe86b7b0e71fac90bfcbd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48cef8eafad045ee731108ad2f227ada80feb79af2623ead75a8d641087d323c90e39a7ebfcd217ae54d1b30b24c18d3a33b2b1063c4c1bf87f2ef997;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22225b81da0709b5c2074237879b50ba39cdd7f1f7d763458f4ca81bba1f7be9354f1d95e4b497af3f1759385983b4c5e6a9e1cd4aede0ab3338ee5e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2860646eca449d79c5e1cdaba4042bc8232f722a9fac6d53017c1e50b10b5f73c4b3de7ad295711f78698395cae5b87f707dc45ab6aa260bd5289cbf8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d2b45611797195c771b50009d86e16aa19a7bdb1eb07a86281d3a87605674e51dabde9398150ce4383f11d73bacc4a63d32814804b21e4fa20f8c12b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h555138539eeb7a97ae14ae7553a78dcc1ef3885179c37b2d0573657061c353bfce2fcdc299ddde088cc969f0bd8ef46de3f57a5efd9417dd2bcb75eab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78e5092047172a2b7652650697848a956111551f48c4404c883026e49e75fb99c464108ecfe84d48b8cabf5e8fe3f87d36c560d8c61605f9efa6a259c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha97029c3686294764eaea99f3b0ae02c9b04deb505acb805571e849ac9fda0f1bdcd807b0ea93cc4e7ad62862bef12a10858b1a7374af6c246533e6bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f9e08af11a619fb3f467d2440a8a1cdfb6126e71f72a2cb78aa769ec103bd7218973d39dc61b31fa276690e98a11ba6ac217da365912ae65f88b751a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb595019f50db08bd57e4b966f4050448dec76aab478f68f86112a995308aa2c51ba2d5818548f00e352b3284415edff9f90a6def5b22cc8b91e1a57d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c33ae8d12e216f33fa38e9f1ccacf95a1aefab35324fa3670652c788f57f6430e6d8528ed6f5f9d135fa4b5dad21ed33c5ef18815730a78ffa86842a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b94d45c200ad752edbe1b73ee237c911da9bfbbb83a09d88bcd418c56a52e733256e190e5b4d0ad2dc678f3e24449e3a967b38ddf007e44b0ff2c09a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h182f8bc6ffd293e2279f5f48e336c854937d168f39c12f4ed231bb8e87598645a2dd5ac7e03b5089c2c1abfb7dab775e944d6701e87bdadbca99abc00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fe0d5507f999b0c64efe81fb6f23884d7e3598317f009ad4a10bd29bd2ecdb63c8c16d3a9856bdea8c1935fc5539a55f9c41b26d908700e6ff403cb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78e7f633a55d5b2cc7dc118a07de56fc63c10f73602644e2bf992a97f2abce14466f8b12185237f7d5c660647a5fe609265cf8239537e24c8ab0ca3e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47c4fc58019b98f69389f7462e07b2db935060e6e687dce77af7bbceb14dcbe552b2acf491b5c48c5b66709131abf1ee69252ea8338f2a59d6b0ca327;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haaae6c47e2d1436bc7f4abb1b393252f4949a47f50747a9fad17c6d1ae20069345cab1bbce3fc46e41357325b2b96f9998002ffa9e7badbdbe2bdca49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6956f9bba57a90cda14fc5c8bb47e452e12345cf09d8ddc57c299ffab4301d27b6652da831a902e2ae7fedc18a3b3308ad1ecb3b759db3516a708dc7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3c356740e265d0656a783c8cfe66fad473a99db52ff1850fdbc2c94238bc2d7a12a1d77198fd742c6dd85188b46647ef5b1920c6dacf75a200952739;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53c82dbf2286a354e47be5a863f92e8d7bab20464f1ec2061d699243810bcc7e463b0a589b9537949e1a1c3eacce95f42201828a65d01ae82b44f461b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c35ec22963b41bf5589d6b3dc68089400e9961f87578a247ca00be63ea62e725349198647e5d46c3d7627930c0ad7cc53cd2465e28bb1da667d6a365;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22bd0d599025f96ecc3042993cbe8aea1ab0afc2c8c78e5ef6c229cb90dedb72f0b1ddc63efd8bb7f4412a42656328ad81328ae077f992a76e7d0a425;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5cd91b1b0de8bc3241dc167a7ce6b912a81b58fce078bb5940059a01a83df1345086b5a674a1f41cc55afd2ff341c7366e4f66c807e5c94b43c5eaf4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h313f7db5c721e64780f791fbc61e94b9d7acd126d4e3f5f9d09fd88cd9ad1d65b2305f70a48cdd43dd3a4ca2523791441c0b5dfdb12bc45e02f5dd90d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43a62f495fc0368aaf89d30c4ca37bef2fcc563994fda4711207ce998b6b7e249b9305fafe746676dd2cb171463ee1d2679553187eded6b76de96fce8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50557dd7915f5e704e531584de7602dc53f193c2f780b9536e4529323805df02bd1a2140af70f4dd2792c6638876ed2c1bf344f279356de7ebf58ffec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe60b0d113d18e4796685b66bddf359fc5ee456cd42bda0c469f63e317041b007ded38aeb12f69e612f008fe4fc23762f5dc2f3154ba0cd7d382403f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35efdcaeccff793d95313c5899d0ff915741111a0e5ef79c305ce549a6f490e473f206808fd0c308090d171998284dc5fddffbfe8c00d2a251d7bb2c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h755cd27c2373d0b1ef4ed75cf905b430a0f84e6185dc3a9d050efed2cfac4104ca751342da737cb8778e8d1769a7629fc30a939d3af776f4043568c79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae882531ed6cfbde6e1e6eaf22f697f415bb98c15ae3428b0f944c7a5a91948f0c7f7e7285f437bf2924fe0f7b2ab9a5dd8323aa878b5535edd8c52c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9971f099dc9acb300108ceacbbd12299e272ec6715a41d9008028ee4f0baa312cb00a1ffaac288ed9a2fc38ddb7371f920f72e12b715680e96e005a4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6447a1b1cc83b05267b0942005a43a0a8f3cb0730d6c2112aecc117e7c0cb482bfbbe31b636558e884c6928a8b92f87bf23add3c67a8edaf1b31b95b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6af6fecf62f6c3baf4d189b83f1376d79d82963b4cf0ae33ccd0e235eb742cc54862c79fb06a93811a2e50dd5a65f33208f2ee67bdf54b02179b6947b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2373150a89e8ea90e20c8334203564e133a74b8f88a0285c3eeb568cfa4f2150c109e33abb6fee0c8a0962b0ff7196255294e1e7ee40ee1945a7ba16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5164cc02892f1a8fa243da293990954d429b10de0b7b99695c7954d38c2e081470913f15e3e8f61ca884a4945871fc0ce839b3ec6d0902e9cd98d6cde;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f7f8012d237a6f54cf624d30dd4d32c42f0c8d7207646e0341315543bf4d1c00869f4a73c8d4450559e1a77a5803cf8031861778a5a639fe797e657;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3252955cfb51ee56cd827ab08126a02ac3a6228f7730ecccab506800fc9204b55410bdcb4c6294b58b84056866eef8e8dbe949a0e43e8519a413d82f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13cbc7bdeda9a5afc346546d2184106e0cebe5a814b32071cd9feee27ad92c9f8e9543a721ec84db6c1df16ebbe3f8f5749bfd13360d0430afb8e9d36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8ffde91e91bf794e76aca7529ae5d0c299ce62d59a546dcd74b95f566591072b03537b714f07481d227790cd5ca0a98b803a3ef6a760ac9050d4298b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d5b53c67a37524adb664367a1c2b727fd28f0c04219ca880a7a6ecde5fe87e6ca27a22ce87ec3603e6875eb594950b4c5ef9b11daaa460787c04a2b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61bf642ed1a19fadef50fa98bbbfe4066f72e5d210d46f02dbd8d6adde86d76d41f1121a06790b68bfc92bcd39ad6f9d2dc8d76bbcfc9f39e60d297f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb071a5a5ee6aa2b66094017c14c8abf0848774ffc8f887976b69238f5708a4ed4856f3d3c4490d0a8b892968b00e1de24b9bc0b03c575076d13c1c51b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h801b4a8b57156d846f51e4bfa9bc97abd9d68f39b6cba727c7786174a0c8f8b3ea6c679161e07a2fcdad50bf0f4131e915bb98ba6d6995ddd30659901;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e0c5de0e6fdb140d0ac2a1c2eae4f469cf91679a28e6d369cb3d7fbf56dd57d16ac01e2509b5b0155a76ab617cd8666d613272ec2341783847d6d6cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddd702c228c6cd3a720735c118600082c07acbc05022638f8698f0445b61b94c4a48e435f35c8881df26dec625fd4dd80668c6dcbb36af54f6ccc69bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81153d90b66acfb25ac88745887a3a444b0200484e0bf1d6cf1707cd5277117469839b7f3dd5cd3f99dfcb28fa0141691fe468d63d78a847ee8c45e7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9704e6a2f0729f49d49531a4cadefa696d70f837ffca9e28012f0555ba0fa2ec3592c8601f00800ac1ba654f2e33965f844cb3be34b59548181221f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3f2b025e043efc5bf06f16a77e2050ff7f04e3820ebf8983e8d9f1ecc17ada39d9eed690471bf37f129f8eac72b65d0a8eac7f510707d0226b228c2a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4867ea331978b7dd8978feddfa8c6486e4bbb28277945bb9116da61fa5608208855614b12124955449f7e973073bd607701d6632a18f205286e5f929b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h299342e6499992f33becc120900dec49a3e5e2df69ad50d863eff406b2cceba5b42a19e1525021757cdb17e295273b4af019e03e8e092cd3a41e05f9f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60dc1c145a7b358b29fbf170d2cab814d737394b5170ca8c36a932966f3cc9d501c3589c086136de41a577297eeb224ce7b06fee2d9cbe5d5ecb9e2e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cf1927ae815a78132db3d6126e984e1c3a18b834ea1f39f28657bdb0e3ddf27d0ee9c428f7e85f2bd1ba79aed997cae8acbfbfcc2df5d062aa8431a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40a1211fe97e9a601e492a3e44e84cfc413c1e2128b6f29b24307408003a86bd79a9d2e601f2ff58b4db3cfbf1ddc7826cc7f0df28af50509770943e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4fbf1419def1ca03009caf7e33495ec7e93ca0ca83586416ec2c9c7d0e629f63a799e9ad5b02b014f40105303e834b8ed2db725d6f3fb9e4327023d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b641ebc1ee0d3a38c33c08a2d88b035d787da710cace00f2fc3d1e592b4db231957ebc8721c4898ffb0f55b666082a4c64a6499138a86a8767074d58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf03a8c5fc3a6435d7297e8bd4386e2ec070ee44b47a8212260a9255771c1d8f527635e478f072fbee327b8989e133d63b99ae4e705770032d6734e73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6aeb8d7f1d82ee41bc9b2380145cfe3cf71b70827f3bcf420f7b4197e9e95591cdb707fe0f857af7a707412c26fc977dea3fa29afef6ee3066b64807a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35d2dab57fefa033d47df9cef7d4c2f50a302a041235aaea26be68fb2829159533e9265d0fec198b71b02b8da10f9e5f2f840d4f7d8449e9e2d2cacbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9b929f6db9b3f7590acefe2395feda6510b8fcc4d9df8f45daa089c2d1d30756aad95af3b8e390ba2e5771ff9a9dfc6253a199e91a39d1d28d9aa408;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had11081a38b473e1e34bb7512a8117bb1f90ac38d0bb00d9d0f9775bb734725b2eaf8f24bd8b0f558fdc335ae1c6f481c0b43424c328c7812fb3c775e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4204f7a9d834f9d229a2b541027f727fa1ba27402406772f7d358a6bebe6b22f3d01f4d354a424545a8369a1788d69d43cf94bdf56ec3cb9094c0f997;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc81f2bc5e43d5050153d14b52d3cbdde82b4e6d75bffc314b70e6baaab61c65fcca3628b675c40135a2c9261969134259ffe2d01ebfe4b082651a4216;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10e2eba524238f91eee48c95cc8e1520a96aae494630ab0fec97789a4fce8b5d43ad659ad2eb2d70feef9d8b433c049cad433b15b664a2016ee3722ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf21384ea01a74a4767df33dd387e1502aed15b6cda2716736a5651b35c7332f99b1e843afa09171d4d2c33a426c77f68164f2caf2d857616e6b55ce93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc19583797d43805db1d0398aee91541f4e2cb6e9c3158a9dd7ccec436b993d940ad1bc7a641527445a9efc119e19ed3e73812a0197a6b654d02dcea3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffa6b8695fd100790a97ac01cc0d75f31b82c6578be676755a254a28db29526f5eb87e92f80811f3ecc4456d6edd062a668e09e421cb81059a9887f14;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16e4cd97f81ede43ee80e12561f358b62b92877f4503e13471e784ea6def0b3027afac064f968d68f381228d30d4d6ce412ee312ae7dce1bac3beb4d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc92e8aaa13e24a49ac37005d37d415acc4c17f20e42338ab15bae9a504dc11f0dc07bd93d3f4d98eef531d46492e76d6c8f329964795e97e28b936d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h810f11e3440b3e6196085671696838f713edfc3ec41476f138836fbcfab15dd783609f0211e28444fdcfd14b7c96f7ea1856739c628cba9197a8f85a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a117f6c56cb43c1ae1f537ac529ff4fb63ffde70fdf22ad37a76686cf5c81d09659278318c6f9d88f3496dff3d05e55627d054766caf8f745776ea30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74de2029c65ed42f6b1bdc135a8b77e6cbf04404b52a46bfc6b5f7bd0182de367028aafcdbe83a74935c52981aafc5aab166dcf74cb9fef07bcbb9cbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6dbcd6051336acd13ebc64c71237036c5cc3874b73c9a01377bcdd7cf9bfcc3d54fb1c8d3e9b24968df269cabcf049c5e779e0b9a66f6801792efac1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd428fe980a928d66c685a2e56dd1bfdc2c648ef9ffece1a0464c5f5921de846385120d5dc19508513feee11fc34e8b0dc0d88f12f00b5518ac7d28dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cfae2dfdcf32267fbe2b7c73443181d2666a4bcb46c55e477b25e7102e3947c6fa6d7783f302a0f8606b244d4eb012d623b0d7aa40dfcd40bf9a7d21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d2fcfd04b17875b11c753ecf67ed20966e1e8556c0c96b307540efa4f343483ed54ced9336a0e2e8537b14d10458534b769cdb672d326944c193dae9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fcfc48995be756ae16bc1a8d87f34fbb632230ce269b127d2a637c98245815e1918e748cb8bac8f7c4847bf95749a7eab011971ac13f9e10608c89e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a62d44ebb70b28546a39e416ed406d938a14ee35381fb751ce29e0566f58ea22a3d96054d40aa4ffc5ffb8dc2c7635a8dbdd9b89c5c42f50a5cbd96d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6692723a8e58ae35ea02810e9b0dd5e10f6a9b25c9a6f6dbb56e234a8e480baa6dc2032c99f119e0248731a7d0fc6b0ad776566b91a4b475a4b009c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a96c8cc04dd3b74af601eae35e1503925dde7a7fd8a75ec81578db0873a1b134e8e34766a577fbb7aa752665d6385b5675f26ff1cc97dacbf59f8bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h986902534528463ce2fee718a7553ddad08138608eb7b376edd8c8a0d7acd9c573192663bcfab07fab52f14638dd0613f904db473e8affbbd873dc01d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2a774d1790f226b4e5706e4f0b42c485b65e5220f52d36de52dc9a15d937706202be6b4f7128eb96cfe8f8fc3c12f02fe97e3c42cc87d8389179d53a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59e49a373c048d7aa137e83f8e5e402a797c4f56f1616f3ae6177e498f8a0218f3d47070399daffc2be5151333e84f0d3faf65e541087c541695e1f99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99400afa1897d9def3d4edd160202c39b585190edb3268b63e560b7d8e10cfa758039a5ffaa2de4e3432ff1cbacb79f4b18f3dbf73836448fcc4d72e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aa5630cb630e79e2bcfc4501dfb660389ceacd33f68bd041e4d39dbc9eb41c512d82d6c9d28adcd3f9d1775763e9a01825c8b2ae3f8f71caa3a66314;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98b2a48ca70cbe359cf9bdb9f021e6dd75a7b1f8375fc12d775c846bcafbcb7b10bbf75b84edb9d04582d91d0252aefb1af14f75b048af75710de13b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bc3b25a50bc9f961439dc4c099043be39ce9633c7b906b4ab59919a1c7f9f884f10b6478fcece597747d799a577405ce2ffea0801bcb62a35fe17eac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c54a5b7769e73aabb92b05eedffe10cbeec009871a21664ad2c0e8098390cfa5192e6d7cc473ab7545ebcc126707d26f0502996feaa8d4508900508b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f6ae6c4febc376a8fa4fc37bf4c7309490d8c42445a6e7a15f8a4ac1097dcef41ddd41de16ec566c375b35facf2d22fd4a59f0b56c40a56fe6480954;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha387fe34597b8ceae4a10c806acb017066744d879d0a8d373588d70f67f02944fa3a1d30029d783e52fdd318d1245d457875d0440c4fdaed1c0573c6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2974b44ae52b5c73448792f4b6b346874bd00a2ce92158f7845ae7dd68b17055b63af829a68a341e502872d1694407c52b9ca0fbd4e6d26cfae905e0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f0a35869a1bb14e0f5f5da16a8e1ff81e089b26e54472c049f23c68d8a5750a32dc016de6bfcc82e11c1de97aba0eb030ba03954c05c3878ab382cb7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85df3c40dd9049b0141fd936c847671f0519b4848cf880d6fada53881f52fcd2618926511ddc898cd3b3878eb1dd4e2ad1d97bad00380dd91e6c1e559;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8399739ab0106ad3d88637de1b6c82dcf4db9d8cf774ba35f9af389e63b04f65280da35da151f9c57bc45405db01a26ccd5d816dd15a3e45778ac1359;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d4fa89d58121c72a11e3518946c5f0102e56a5395220eff63fbffd11c021a8d31c7128e550e698ca124fd0f82c2251f838b8f63b0ccf3df203578402;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h249196251f5a94386c2b66239789f9747ce2ffc4ed58f1135cd554e866c2db79e35f62223fef8428487dc4c72d3f2355ed6f0db2f3bcb37aff26ebb7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d542063a2b61005db582865f97c3f738df4d49eade8f7bf7910e6118371ea26d758c72834c574078bcaf27afe4feae887b8da42723912af651697b92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b453a8d3679c04ff4ae0d0eb7f5a5ca40ce2013d3b6e1ea05ea71c5be7751f884684ee7ab36460c1b189defdc87f7abe89bb87a71f66b13138299015;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9e9d5f2328f3a6a548105dcf82337124f260b9fb33d6ad01e069be441c81d356984aee7935563bd7e2bb1119be83addf250a95b6593277744eb67f21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a3d2cb6eeaa2fa25925a8cd7a5a981ef100150b421c6b0fe845e4aa2bb6b50a1ca16a73423790e2a80f3109d69c1f8aa927fa62b88a70c256aff0f4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79074fa06d16f33e1584bee076caa4f3e5e47a9432cdcd0d1a91a23a1b0096f75916e88c317373e2c1c44576a777fbe67a5329414bcc753dc789694e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc5dfc1f42c3c7da631fb1081c7442512a43d8af0fbeacbc9ef021febc2db0caef9f5abb1a341bc34128616f535b8a2889d7bfa20c2ecc22f32aec96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he905570f10299e7f0a52fbb180f1c61521fc7e31b5c6b72c5c589cfde42e54231d23b2fba605e390d6132fd8182eda1e1ad054c1b981bb80a5b63009d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5c21b640595c78acd44b3cea0a3d2a8ae293090130ed1164c947f5cd21171a6202a9418f21f005d7bf1f98088685777b2c1f0675d6f82aad79b16993;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b60256c498ac2b35e1c546215270ec8dec4dcd9a2cd94000c27f5622822be72bffa5bc0db331fa98f36c84215b8769eb566e28dcb8bd312b68a80fbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h337a6989d35e31c6e14e4f2e760d83904e6d92e342211ec8a8c5b1cbd1fd671de8ddd0e5d9c1841f8ed85e9df6c5d687cab12fdb650120a0691d11d8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcb7bbaa85eb21c1372ca7e1ab409464f1a59e7442b6ec5c19236fb504c95da7f1e723c9d5ee280688bc22dde99b80de2b7f8ce7787ad5fd6d924ae67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87eee7d44fb4f18b2a8e04f485e144b03ec4235bca1092a2b647190eabd63d27e67ecf960d12392dfee406f3420d27122a053c69dc43e7b25c060bf53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82a8832008a4bdc49c5f0995ba5de85911063aef4afa3e764125c72ccec2bb67f2bc44a26bb0f0df85c394052b6830199eeee06938402a4b2a59a0397;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab015454181b8bdc1d2c128d6a178bf39158ef0cba32b89a050964779ff856d5c5d2bf270a027f2e6ccb33d1d66b8baea4feb6fd93571a4bd8352f442;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3cc2df08c5b6f21baf39404e33d4828c0c4d35ca4b19d2ab8bc98005a3945e9807849d57a5d6f45723bd5bbfcc8e0142a4c3e4b57dc87f1541eeaf0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2c3cc98860d10d1f618f94390b58749ebd67ee006ff48598aefea2082274f609474499e3013d5f90469d6d00ec2dce418465fea18514d5d762bd4fd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h124dcc3300960de459525ed1a6c3ddb10bd4b48c6f8e0024ba6c4555c36c5062b030ca29fd064a23b7c66a8fa98583e0126b59dae1dc658172c67c690;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fa69ba191756393f32107e71bbaf7e3dbd4156b03be86f0d741bd1109d33b80314f9be3206d79b6a62afed62bb58d41a656d9cf634647024b0fdb549;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a493f3fd3a03af20e0f7cccc1eedea739fd89382bf5dad5c5f1aed11b2c3c0e16bee04239a6aa9c3e8c08d55bd1bce609fcdce5463c6c9675ebe91ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3cbfb709b808e8c6b7321cd4f58e74c5306dd032887b44f85b5ad45b64f89845245f29f7c7c5eb7af527ae6c4384aa1ee152d95638bb571c4e07ddc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h485ce415cda0442ab1d591ba583bc5a7ba88007051efb4e611f9a5b795bbf3d7c4b112d777da37572c30e54e1e426663ca2b63d227d7dccf80f0d002d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2517a3511ffd40317a248dfc593a0733105ec4817fd75566140ee5e05d69365bd6e7b88d3bdd2097628a1daf4f8f60cfa78c8589e8c530045a6c15c96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68f4814812e5c8027bea099cf6d952222eecccaa844ab3b82708e1d86cc45bd98eed11412fadb12433ce064686c2b1fb4662ff61e468e71a93f591fe4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff9b1d982a9fb7c219e35f5d48bd7df855e16987980f5a9989290858421024d40d5056c2c9f4ecc2428a97ea14ba0e96b04ba1db7ecac3022ea9b942b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86e84c853dc9962037f6f05bcd8c087d8761d3a77db7bf8f9cc720aa0c849cd914e70d9831a8996eacfbe178b2e59f9ac0749fa981517391f5e324173;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ab6a74a7f53602c795b7db5f9b0fbf3c32dd3b8806119aca43bcbecd710a10f21bff5a599dee5cb26ac8458323646d20f84af1ff17814d43c24b8ffb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4cea0bb21cddc777138a1a2a0126c8ff14a08ad0ea8237563cdf5c7a2c42c73e00e385d73fbfb9395184e29bcf76da4f93478205875a4389ea2f3a60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf30589ba86dd50a0d8eb645550f85aec2c1ca5a78c06757d4c9f418b0ff50c325177ef76eff0c845f6d0a00b2eafd80cf88ce865b35c2df73b6e93991;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92c68094e2cc6a596be9461427dbd25985cf307008d579fba0792ad71513e01dccad315474c9f7a5884f980980a5c384fa77c431f119578a09a4e7f18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb00fd58473482e2908e198c420e79374b3ced8b783292077729635a20358da4caab5df5c42e142100cf56fa828faca8fda6782c0ee75382b938d394ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdd2e0aea3d2da81f24a3ecb2f27e2896874c6b1283903b69873f9fa15d90b5ce819ca7c7c883d5f1a7855bae757cc1873e813c299822620c74932a97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e50f84969f096089b83bf53f3b3420a309ea458c2a11543c5bbebc8b0920f44d7c0db3a68a41e90319c68ec9f789043d6ba9d7648bff4b271a5b4878;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa7064e596dd5f6b3e65a83156f182ade5f972cf8d2a92182a95f88a2107074590ba26270574ae022b05dfd62c2538d99e2f966319f4af7b68810a04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h710fd8937b04f54ead619be731b7fad98f8ca70694f10f152173e77eb79e017e05842480b7998835804fe95e40672063e8d8c7340ef349185a95ca790;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he114d055edd138e161199f7f20e4c554daefdb5191e5e5fca8694ea864c8b860a028e5b1515e075cce4f4cef16208f3097329fb7e2f5f4455bb4294ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2debdc9d6b75d4d6e12c917b252d9f8807ef4858801caa39cda32fe8d470cf046ed70af3d10ddd242ac3b86858e8cbf9ed4e7df906c7cc72967d786b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaaea69656a88339e811ac820ffabb3dbfcf9a8fb9c60171286e101c931eabd450a344f85434b7fa162b393484888733747b803db65c77bc870d1fbe1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7f6998a108d0eaa455f94cf4a4a3fbb057303c0a7614f85ea522233d8ba24c5d95703263b02e231a0bcd54aa54b5fa308f2232dd149ad0ecb0b6030;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd80342d2f527701548c9ab6f27d9f9ff62d61b277095d0b8e7fa5c2dc490ffc22cd278c5ba3db6948a4960490ddbf7bdc6cef6fcf86dd1c6b8ef6fb29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h435e978c7972bf44b93cdcea9ee6df1e6fb2a9656fb9441aa85f4b73623c9817f1acff38d9dd8777cbeee70bc591b7482c6b0d8348dc2260ea1a527ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a5e3ce6e0f41ecacc6663caa8c3bb3061240d1d8b0309137f88c6e925921cd46787c24b35c7b0761135b8f533d28a6c2aec37ce17e9ecd5110ccae51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6c1c3e09e42c3958b1d16271a3c256bda66ffd5ab9fc428c842d1eb5e544ae69c3f58cfbbde1675862df122fb1a39b47ad67abd35a2a1dcb8a35d993;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdc21e6e73a2c2fdc96eae7372258e99d8cdfe5b379f71b9d40670d898aa3018c89b5a71998c0a4324ab4868300686eaf4fca1ee74d2ca0139bb2ca5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha744a82aad9886de0635c66ea38be401c456e60c2bd8c891532e4a9a6d97d077adc2e97886dc2cf90e525d60c8f5ef073c4aada9a9f5b9519f1486cd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b6c6badba6b1ce4a21cca6dae7ac7084a3b2eee52de983707fdf4286c362ab496fa576c46f58ae75c0e9a0ce4e4cc5d774b36049c4bf82de365822d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff539bf61abce1f2baad95cb59c5a1fc2a863073d86ae17bbfe24cfa5396e40ffc54b0e3ac9ea80cc744804e02d227fcd62c8c9c5ecdb7cee8f2c5a05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8fda065a9ced54249d4bc6b172bf67144899d7a661df4721e42340a91f479e5d05228a372e294ff8b1aae20055ba3d3b49fd203de311c482a924fd40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd076066356bf990f1b8ed6c996bb6fb80baef6bba8209b32f6e3eaa814fe8e59b6b6d08864b40c79dc6bbbdc1ea2c1dff86c8b6ad51091f30895ead17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77ce7bda46f8e9fae4ae49c6f0196450c8fbfe6d434e6bfa78db5b5e98acfe17077b3556e1f4cc1c69d656cb8fa4bebcd08d3e43c25dfcc2771270363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0274ce6473656bd811732ec1151bf72b6110409d6d9753d447960f07d109481afc2b3ed50fe7900b37eaaf625682866e0081677185ae0bae413b5b44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e4629791a46563c767557f88fc1f69e71e46e2a8c447aa375957228d84823d419a97439539bf39618a53da3ded514568f85e24dad18131de2ce0a0e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefc6457f356ec3565171062f8a6756acc178684259356466acf7c244e988839fee98f4461a65adaf2396ea8bd694c41c97316476e4e50af981c52662c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f983725ed8a44cec577c27cb95d4853c36ffd25adb6de3caebd3716289f70e7952a3359771272c382088d5bed3d36b5618852209f1d4892a90b01e82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0319079a67ef135e6267e38f0ea75e915608708d895713fe1be03d28db59e2d3f1f3da047ef5524900d9f02cad7993e027ebd4c5c276a480a66ea1cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63b31ef0027b96e38e90c016ea6a6790ac96ec90dce67508a81c9bb581e31f006d9cb94801dcdf23aa022deb60c751757377858ca7595ad73d40615ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h655198c774b090fbd1fe6affe52e3f4f8ee06dbad97eea5cb7c7530dad5b71eac18e4e21209f7e9ade46d31c418def752f251e3028fc8c6e4f980cf4a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h757abfae2373899d7f847042f1e1cfc2631b9013f727c414a62bccc79d2870dc49bcee374c71b13a68f518a8e5a21c1800f79c7221be2d96a8db60824;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c571075d678b22798e08c18d6aecbb4912bcb0f364a4f71bf9819fcf0a90842476f6f73d091b8408b646b2abeb15f54de2a546e6c329da56e8ee9a8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bb58fca52491054ab4d9ad0ba07b4dce76f213f4629ad8134e8fc2e0848ac235e6e8f09fea6088e5ae5ea2ecc5614ddb0f3c8a7c0bbd23325d52c7b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79febe7e60a9f97dbad5a2c7fed5054665b2489b3a8e618c57a6238876034aea5094b4961df2e4c224856c53177abf6c8f5e97e3d8448f99c9525c13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2bf244150179c8ca608855f97ed858436a5b239efaf0340f03a0553dcdbcf8fe80e78a1c864de4353f607c4d163b732dd62c0392bf36161acff2b33b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h737f924406d42169383c10ea2c7f76dc014a8f979bf5724e2406eabe90725c038dfd2d26c82a7253c1bfce499d6bf93a2656b27841ed1f6f1108feb90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9bc1716e9368c45045d30f627a18f63da0113d1c36dd1faff30261d6f2ab4b8d2c84d6de93265d786a564fe95f6a9a4ae924da29869fbe5aea5b6ac0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb34050620e87b0c09227bd3629f64b6293be45c8a8670055037c55c6575d3227335b4071eb3c60583734c0a6caba43b2286eb5de6a4ca8331e5ca919;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0f7f47b8c95c1717b921afc081219f1fe0a6a409738f9adce3963e8447966110d9fce5c6f63986ab7cf9854ada5fd2bdc978122933b3f25679a75db0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe207114fbbedb388904a548e692d13d93f4f97f8659e36301d904f391e7c1f069e64783669f24b6879c22b85581fdad2c99e5fad5a334a333cb48f7f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc7f99939ecb468af2f4c87df21a096f15ecf88a95e31e85e5b4e180ab322346003ea2c6500b500e12002b046d7a579a8d3557ace89efac35ddf4da5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hece7b017e54c42dfd9387f3ce5b9b3d3f55e1f4ebbd9ce831f85c1198ee2efd76721f3ef735c4eb249a6de26fd27771bf33a6922b3a546f50b8a16ef4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7a40d82290526b4157e7aedb7ca518236fc550afbcd4a012773ba796c0a2e28626c9201ff5fe8c40c36887621360fce2ebb28902d95f84d8a1bc986f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb0cad3f8a1cebe5629a7ecf9c825e71e9a2936b69b945f0c9dca0d0c2fbe87ad01ea9966fbffa9457ee885838923b3418318983135f520afb0cb2fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb8b380a3792f8eb0e1334b60b42d20baefb35947859fd9a29a4db81aac7f559ca6443c488a451e7e6544b188171399c8afbb54bec85745efa6c07eb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2b5c231f69cefc8e7560cb64d7bcb4f104ae79d6bf80c6fd2368d706055321a3c46f6accb385693d1bab2b644ef79821090309e88d35fd3e81cb2a5d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0c5f6a082621321a69f6c9a145dc81e09e9e1ae124e3a4f5ff81bed4a40519788a7bee778dc986f8fb46d3e0e7d91ac43d54ef721e22562cff30da4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e7fb14de4a66f00d9889c989393853a8e346137d18fd43ba0297a4049c24bded37da70716258c0d51f8e4ca84307bb9da2cc001943ce032c53948c65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h431d3e6bc52b4c66ca4c06d1c5db696bc8c8134df3ecc5e4b80c52cec34d88039ad1c19bc605bf089a44a04558df502f0e0b21e2de27c19a2027168c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha134d59048aabd843f0727349e9e054418959759cef5c83ce8021074998c8d076dec337fa861443af74ffa18b4ca9723dea7714aa549baa124bd5316f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b0c2c7a9d624f367498888302d9c04876706e3d67b2d4938d741a099ee100f2f12f56120e526b98cd8cde8e67c4efa00c7a55997eddeb47202156ee5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa57fc0937c62e3e28f2d36ab44856ed8a66237b473e5964cd867ba78f7deed7cfcadcb39b4f97a2a355a3ff5694a7b59e3e5a62d750f06a1a5a1a393;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcfbde30748f400d6bb31862b9f4963e2157bfa64fa685e78eac9580a75984386d5ca5a4b9abd0566bf6b447f01deb94ffb8869185b91074b33b32c03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75d363833a3bee0750a5a54051bb49f96115cc8f5819130cd586eb8cf25707f76dbd3d5fa65a248c9fff4c2208f57b5a4a17d267e13e2dca6aa69d6f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h364cbd8f675810912de2cfbc458b03f30950bf363ace0003c6382ffcad4a06d67fe3271702b03fb17620e4b05e8baf555dee05c661027fb943a70a2dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42924a27295bc7202bc54502bd77c8ae1e5fbacd83015384ca3e3115f30b088d7af5a9a9362b18297feae614ff1b20d5755540cb6e5ca397e5092f673;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9c5f34226e950f8a1ee9552f5aec4097c867595d90506cb0288f94d31d5ff7cd5239c6877658df646f2df1ae99b4f306505a51c463dc47983267e7fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5829ca469a5a7e4211b7f4754653710b54ed64fe43e49dd45868c29f0925ed223a4ba95a2357ab7ddda20a0e94dd3f24b0da36bbf7d65a738983d35cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf331c52c7ffbb67624a22c6ded1e4c1c312b7e279899cb2b6522d8e33d1e144ca38000fdb9077ebbbfda693cc4983c3d1116bd12f98dba08cae97cc8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89dfe02cae2b268d34edea037931217eaf701cf236b11bc279c31397bc9596a57f17e8c7baec932e2553eadc436fcfd0dcc69a7a1d606048c694a8fb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h675f8dcd4778ec54f95c13060970b25a35617643a4323006e1c49011373a64e1091b9a5081a3a6f50dd7e5e2c87a0378980d2bccaa2528b054aa6d00e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h685317be1f3754692041a4d7130a6b7cc52d5204fea00b5947a65e30cada8d40a9cd6f544d0a4f7bb677cf91a3b8366fada74cca717bc749f450e53fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c2a5b1bee3f6278da43a19cdc0c1b837eef8ef5ca03f7c0e7736ff634c02dcbbb45ec0083de401104725260f26cef5200918f91c54680ea81bda8ac9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82ce8a32a72bfb44a998dd88c357382d1c118f548ee09a79ba82e2b6f6cbdf9c8dd6f31b298be8ccd060004eb0d32537580e4c2719a7fe74d8ce2dec6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644776cea2ffc8d0b3ca98d5fb8df52c99cebdac9845118dd542987e516bb2b73ce9633f0a07b9c6fd66a08b14bdded2452d962a687e8653ee661c63f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he446ec61569b6205b1c96297aa6e2f824d5c85854221acb59edc225bc1774d530a6bf1266ce4eabcb6cebedbf2f7b1866500c1f7340b5f97cd565bd5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h715a3f8196b5be7f76d8f319b05395e0331aaee3b0a81df6c56c9991ac96df23d305993173320e92724aaf7210a0ece3a2ca2bddb5f5e7b03fc119fc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28159e1b1ae29023ee31fe06b0987a7f99a11d009e9c362c088a67eb101ff55a664bf1884dd04e0e8f556d999fd3fbc885eb210bb70491bc31db4cc28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc51641077b7b20b81e1a90834b5081c4adb4ba9189045308c8bca0eb5ada63a05ca794d6ff9d7e8fe058aed8060ef4f882b30591e761e953784343a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h669f355e5e9d9ef3ba9e34c1420372ba5566fa21305f5e74d861f285a3a447b8e3dea6f4b7a623b63ac1003408c3367a546c8d7a0b734bf299a03954b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57addb65d872a7e2bb4f66a934eb9ba84269444f990fed987f4c1dbb90c98c7c4e24374b1f973c93907734158b0076d31c51a9a899bed42b7a1b2955e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fd461f44a2f34df3b8dac140f4246cf043b1da5809291b22580b09a51609fde3da1592e455d0160559180f536cf460459b3f48b45ea2749d1bdb1936;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h765e25e15aa53a2e49e25e710c2f9200ecfc0948ffeae3dd2c090d7995d3d55f508000ce1338cb8db622cb796499fa9b78b452e7dcd8f7cecfcb558ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h253dc1bde0994fb906e3fdb0f585798140d8fb57c5f858dde568926758d8f93d2a55ca7b1cb76baf92a54fc148df3134ae2a2e912ed311fba24cc94a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h822abf012ae6c24f9c86f157d89f45c4dc6014323f1e50d3edf33336ae83ab034007f86aaf27b7c02fe007c1e9c8f2d9f90023268e173b3a02f4ff903;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7edfc25dd7a7d2e1f0c04272bd1bdc384fdfdefad70c4c9e4bde6975eb2335ad50183d41532051647c26d0ddfd5accbf14024565a732008255ac662f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h197aa02ae6dc816d4549b7deba187f35a439e8b2b9973fc92cb0b486eabc9f8974ff52f51d28c7658a913140011cbe924ae511b0c3f261dd8206be534;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c3df4c3789ccc554939d5563ea81e1cd01af43813a5868b1439ffd0660061b7c5d93ee01a3e2106375c2b457f4d94a25b455039fc66c6efabf0ee4d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56e28ec8f6e393349604409d30f7c8b4d13e541b6c3168d094945a150fb8e285017ab6c63d60f6d8586218d1b6ba8703e88709156f5b9c4d34de57dc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f48dbb7e9218e40bb5d21d45ab4eb93ed602f624a2cafc5985ac674b49764915a0045ab12918f3b0134b179e73a99cb6987068d22f954c9b083b12ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd4446efbcacaff05899317ef1ef68d7ac3a51563b16d06547e6ca0a45e9389b7733b7a06c9d26d074830ac9fbb18b149c65c59917b44f5bd916187b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25bed09ddb241f4178c80b3a3bd9d8c814fb9088ec07d117539f260205a518890e6c3f216a499f6469ada73346c20f27f6308b843feb12b9b3950a528;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9df97c4da9810acda82db5f4eaf40baa65fdee841bfdaf31efc0b0b2436abb9a33ebd9925c0d09d0555180cef16c3b488194bdd20bb06dd384bf7517;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc6f077b489e68c33cbe87a32982b490bf4c3373415aa549346355eb87b62ddaf272655349bc29a0323c5ba3ba9ecbb28321f8941bc7ddd1dc1d8eb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb66a74be4f4e5d282934bc395e525f52353094f9c121c71c04ad4dda31905fa1bf0bb953d10b35d7a5b49b68e67bfa2894c512dda790ad6efbd375c03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h313cdd9b3d6f3cb45fdd60bfd3625fa8161096b4b60936a8d7440b47a34d24883d981a89156540a565a4f45d892988d32a3782aa1cd5af850efa77d49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda83b804b23b21c9b463023a48637d5b0135e830ab04442bd69542ed715669424400b485e55e5949669f2ee37a923ae1b171953ed82628d7e4a5d6f2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d630966fb0c70ac7f0192584cba34244bd4199963aa5ed1ef1d1402f2f02686dc8d92cd3edc4cd87ae5e92f962c6be32c6cff20d77209795dcf161fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1244cc0ed9a720f7631ea7a02cbf9403697985d6d96adb43eddbd0d5d534550a762b839cb1784e2840d3ba596178ed59fe47a8ef93edcfac619081e64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e5e5636d44777454d554bdda13c0ba69ca150af01533ce302ff3867a4c60f33f3588adfd65f98a7eb769be0ad7e8849c2967c59501c7603085b2d92e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd78545b76d5d2b483b1376b725e572c61e0c6f2709d44991fe71a14da58ec4d479a99532d224c033d7a2fe031debf0e86bde3a76cef829d93206c4d9d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9992d1808f70782f51c2221dc02637a95eae00f3aa390a068ec0692bc5af84a10208638d8b99c3d4709f163ec3608dce215700e9411547fd930409677;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83cc5da177fa2a39c7b0d2ca392bf04d9685ab1e4b3e7533fcfc8afd6d96c35b0a403e60ed1f7bdf4a85aa416eb9397425ed5d7ab888f138022432ee1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h767044ed11c8cdbd799cb528df72405c05c05128a52ab40ca8088bb1e12308b3e4f2a3e2e0873d1c5db7d83b4f1d0a9d22661cf779f261d4d0941b328;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0f11936eb010cef5f4d697bb256fb8a2bd228f1c975b7d630b6013f94cc630957ad122dbf6b4907a048c181a21bf211013e4c1cf516d8802b34b1733;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd02f258a2d6977ed3feefb95dee87e7f7745190cb4e2ec6743fb4853497a034f65a8a9ea31a7e5c07b6e0d82e55d1848c5dec11f2a440671e68ed0588;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a4eaf5c0282af632b7e8ae2484990128bba1e7d1d8610c8dda4f987324b12e94f4dbb9d649a49c37b40c5ea19f816cbcccbd72e45e630c2b36e46f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd17c21ed47d693798ca507e665ae80c78860f5846778457b80306e94bd64e520d65c3ae9bea875aac016dfd505a638b9f467cd928100a66f6f065f433;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha89a09b96cddb01ea488b234df4859f1db135e1e994094de830f0d4da2ccc790d7f035954a4daf92d337513ec62cdbcb4d06e107e134627828b208e66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46703cd1af673ffd7698bdc92f1627d3ddbc017e1a692c2e38c366c31c93340c84f1596b71e3e8b87af8be6282cb0d09a3cc6c00f152975aa8f4b8e93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0532698abeba74feb27e6f563d17713d805d2f8d6166a1afec3589d3c04c39b855383c2df7476ec13f691439f67903332c5273d9e680f0c47eef9979;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30070c5e7c72fd78e88dd139698c74c99284c1527940097ecf15a308a75a4e8dcbf150ffc124a07355ce11872943c4a3f4e11a73a5a85318213a45038;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9f80254522d14a0d7a6d642310f097182c0f0bbb4ef592eb7b910d02fb4ebefd029939555ef3db693fae8989e8652b0d30c71495ca17e6d74f53a80c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he433c8200ec16aaaeac2a5a2e0a5972d4e2fd56c3b7ca1167f50663151b23d7ce37e6a7de30bac5bcb32628dac60157ebd8019ec95d4be9a5755ae73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h703112aa97fbce06c0fd6b7b462db241636d1367ce8dd9274ed98bb9c0bb110c827f2bcce8572ebfd8acb33149fede587b1bf7cbb9fbe86ef5436752;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62d48bffb527693059d6ce67c01c05e6c627769e64858e791844fb52199e1ae37ac2a130ba5b43547375086033b15c6296694b6b79090c0bdcf1d18f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52eea4e1489c58ed49654a0bea9596ee59949918f91be4bdee14408e23faae3f793240adc3eec37c07869d38537c025715901f4f196fc026ccfc79ecd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19eb4b79cb02a92a1eec3585eddbe8af2550b183fe8580ca9915d2c83c057455e20de56b1de3c9997462e0db1bb320033c2fdae4c108773e55bb895f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ade2e46a6d72eadeeb2520d5184a23727325f264dc4ca18b35cd9e00993d49fd04b9e8aeb6c46a9744e558efc7e3284ed72ce2eb52c2dcf4faee8620;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37d94ba76dae29e0a484e51a1d470637dbea8f488218c90ead24295b2f31bc8ae443459caf74670fa7254940efafb388e015418f3dbba535294ee9624;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce4d069aa85391497c2b31ab85a7edf4b65dd84ddc7cae5f2902551b528bd98bedf8fed48d2b941cb2ab5e0662238668b114b0d37a2e9b20596483ed4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea546e897e2326939ead7fe728ee4b50df38e55d39f6c3be51fda04f404aa216630f91a119a21d11869010e678929d667a457972bd6e53e6ac1d93482;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4f1a0d6814f5cf2d7cb939e30b900e7bb83836fcf695bd9a19629ff037fd55138ae8375f96f74b957e210fab9aafffb02b4265980fd471efdb59c0c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aefe1e81db523b8c0ad78e16be432f5cc5fa7d438b8499f08c0c1e871eb34f52913dd6a5dc180c36b0c236858f73a454549702eb0a033dc00a21ca14;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7da49af098a72aa9c1187d2570683d72b04f12bf0550ddbec6d751922d01d972cf92977ab7f9946c8373e34a7bee1ba44a73041db8c1b88a535b50767;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h830a263a8b6552e301a19b26e6968e75a7b79fabe02ca2865a81685266f6f1068d34ec123c3e1815767eace3a2415f765676c1ba9b60c31a58df51d75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcce8794abe5e7469a004e3e806fe58fa3b3d24885962953d2cbf01ed430e9c4ce1f3bd896c19c35a4c2e728fe0fd5a50d6eb1501138a39dcb9fbeadcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h618116a07cd47996e1b1de1f7b3147006c7a4b6f31992d70f160053ca6cac46b8d4297af37e929ef8419f9c2ca9add9fce912d0dcebddc35d441d769f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h883580155c5a6eccbfba6e4e00a03dfe7707c0c6e7ec97d0560d72639d0008a55e3efddf0eed18b5127a338c94bcea2d54e42984c879f4ddb7a98f27;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd30f4e6133d8d9c9435350f61fe825625a9fb7af8629b8b8d7134a3d7aab56fb183c7077c25dc1f786f04596987cc84ab9303bdcd69cd4da1c0720ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14fb67f1ffb4a23c36cc937ecc0720d59c4771f84d52716a87a04849b22f9213bdfeba2f464841a18eb7470062f8728c282940c98a1d4c49554deac79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h344284e88752da16245550ea69134c02604a70324bbb7465af05d908008b3a1bef336f8f7ad533f61b0aefa76c2021e606e3e603c7cc9c0901a3d6309;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5ba8301f4ae7bc1c9a50048bad190fa2fb8accc46982ef3b2679e9bfa3968be9bc5460a7aaf3c12f01c733fa4baaa2ead0b48bd34c2844fdcdf3b9de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24ddcff25152d6c5b3ab1e7bffed8962f61798f48fe720ec210b01f1a93554719d3b70a38b9ebe2c7610617dd2499c9021b0a3ef32cc0dc211d10860e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2054b9b3b3e7d585eb731b068efbf7652562289e874407d3b9bbb97b9bb97d6b2a3a3d068eb9faf86bc51295d301f2675d6447feaa958a2dc50e488eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8bec439267949cb57410527f1b8aa3260c4c8a8fe0c938750fb1f9931df2c2f1e816344bf1b17b9f51ce180d6ad26f191d824ef6e80590b3381e651a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha77f5e67e4e1ab856de06f74ee50924c4a25284f5f4c651e90d520802d6d98dd074d8d3c10642ce75ee4771093f6e59f7173409fd6050e2bcdd5ab4b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3181cc78c154c5c08570ed709106f2756c7c52a98e85bc35e2d00673fdf81db511a6e55b72f5e885418fe37e46d61361cdb0d1a9beb772865bc84311f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h456f1a7dcb69b0774b834bb98b924f485f3fddad069926c36e1b6acf84b204a3a9a67c1c5513d7b0fd69ad3626add2f1e67beaffbd9899ffb0446569b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf87dd0a43a1f3658bc0fe03094ed9e882baad507f8810b59f3941525a653607afa88ef3f148eb95393e23433c1081d201362c241d261adf9fd483d79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4193b5864ca56cf586cc5e253efea3b9071e6c8e8834f7be608d6eda1f34f0216f479627e149b500d021c6b6e0ee5540da5e96634914119e24bfd6f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a85381c73b5bab66e35a6b7fc75af9bfbd7f86f083cc8da0dbe744befa876c156040422c6db6b76bd1a91a8a359e0b41f210b5ed286111da87b3c5cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h132b7723dea07adc07ce25e23167df405d033ce5494615f13cd92737b8c4644233b31cd7c85f6712e27b489ea26d1c07ee49dd7e38a52cd7818c26c09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91a5cbaaa941e68a3a8d54784e3cf864dfde87c60ab69eac2eda5f550d1b3f7fd119b806629b30944043ad5b9a74a9c2a55194db82deca9192cf3ed48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90ed3e454a2d32a1f1732bbfc320c4276bd3355f6c47a1c43a4213079b596ef454807d60bc43765598e0d8923eb0def907b3ad2e79c42755ac1690586;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h912ff8bce672c0fa8fedb69c6159ca957049791f2f14861eeffc0dc0dabd2a9f07846a903b7de4dbcd9b3eac3f8bcaa61edd41390c3bb2a2be8095c1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb376d92aeea7722384fbad9fcff556b01ede392b1746478b2c3355933f56860262bc28d869cdc9bffc9203b75bce0debe7c9de0b2185eb38571cbaa00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb975862e8f051dc72c9161a641fd7ece2354c275e08aad167465927805501993dcf7a71bfcefa35105bf538974d95208460b052bba38b239334e7abf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c52aafc758a69755d62270097e3d9922ffd2915251b07d81fdbb7871bafd3973810f8362ac683116cefe95e9eec468c70b379e34c5f28e401446a73e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4361b1675c13f1d99a3d354a05c1a855ce825564e00420c3b6084af4fa0d5a4b180b371d18ce77167fb011ab7721b2e9f35b05f5900d5bafda9e3d527;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e7b341b3bba48fda96ebe66b968c23ca88589bb14bd5e1a94666c7e2a19832106ea0bf97ee2d2751ee4ec3483782ec1bfe210eedd5d4101c3b0b1c10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89d39ea96a17c7991857b7d8e1f23283141dc791d252bd8c1751eaca98c408d9a9e273867e362d9ce6788b521ad211ca2035f7f71393dd2b1643bf641;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6787ec25d9c372645b319954bb9aede272453c4e50a993c05452496ecbd8cb80bc82f4758bc379eafc1629999389cee987629ad41e2e2799088b901b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ed613936a387d5ff69253004f4971227565c45cbedee4fb9ca71b95ddce33dbc2bc2b4f56a19b7bb534075999c4528845907761a772542496f3ecf40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ddd0e0bce22ee4dc1de936d8eed2ecee5e631019a6c6c5dbba2a36e50ad661a8439ae29ff706f73b75e93c5d04083e38bd15a22090311903f1d09a40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb1265f35fe15855a1b03cec4d0a47cbc696451f3349874d08c7516b82ba8e3b604324283da2ed995e5e9b4af871d14c344218f8156542b55f6904a2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha72560ef32f28de002e7b979de6f0adb14914f687e1407e077ab2193bacc63670a443a6f7c47d4f97edc5bdd607b3ccf776f5187007d1912f7efaf83a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a71ca1a82b3848f47faab0506a8f4781c3a8bb85ab716d1ccbe61d9667be85d424dfe0f2a47835f565aaab72c385efdf921a43fc1132dfe0239c44d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6e109c0da7b892793485e46289e73a4e3ea26a93febad89e31261fdf7385dafb06e141e3c069d387911918bda0bf0e9ca07cb9c5e4bb851491ab8ac2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82cac0d8623e497e18de3efef715683bb0ce295a0f01a536fd8f720ea63ab8699fa3a8ec6a0e34cf36316e704bee684712a79732ae82e1d381fcb8600;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bc89dba470e5bdaf0c62a0a0527ef668cc717797e2ad7a96d919cdf9d215defe8e45b923f37073b96368ec413310cd6bcc6e7dd60f8290715e8e7645;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4baff9839e4aea0f13037b57780c6c7899a5f4a2353493995966b767a579d76c1584931ecca6f0b9324df360ae9f8223fb34d83e36e67bd7f4d64b1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf39b2a8a0a28c6979e54491502eeb6ff47f2eec565692281a213b0da0278f054ed5692c469719317a576c45e08afc0189ef55690795ffadec62e73dc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h672578aa44a00684142be745a3cdd199fe0ebd9d9a2317fba7459bc172b91bb2836ed2d67e91008a302b319674ef50e645cb7bed7975a07850ba0e283;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha900ae61fe1e8b7596ba69230dfbd7df869fcee66012c579a1379c6c78b201abff0f4b2eee46f15c7472497b6cc7738fbf756feb62692c8fccf319478;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h812e6aa1804ce41375ccb10d9e0d99ac02b35b1877b23fc958bbdd20b7d6f88108b7e115e999ce7820401c9f79c918a5027ac8d5a030cb64c1170772a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4c72770c4c6da86956dd4a3d420e4c071e836461aba8cdeb56562270ed0713f1ed98edfe645e8a53c48c4569f1e285dc769c1735d6044576c640e042;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc10e5414fab19584c74c1570c3ddb3e199630333c70d1992300b6f5359818318372dbba0eb7c57b1c9bbc3e8ec62ff502cf18e379ab52330d1741918;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ea56e28041d9c6cda55454ea0d1809524498b2b931dd1deb20ca303e626ee55f04799a91d0d0277982df3f3fb794217d5f56e0704f386b6a5262c5f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb35bc97a0994f6c3332e7324b956b1d43aa0ea4705becf068a4d10400da5bf6c31820541f5f8633835f632006c678564bbe49f9e3f35e64e6d9ac7409;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20676e219467162930ee60de8d3d5dad56a31b5b57359503f5a558c77f47ad0eb7a10a1d12a5f551ab689efb3d1b147efb5b2b5d6c0baa508929af3b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbaafae93e83298a7851cf31e10cf762e8205410e0752cc37e8bf4601d23dbbc34c8ec18e694b8fea747ad39be9f187b75415e8f080fbb76c31b042016;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51234a78cf8aaf1ab55064cc43e8e97b92f03f17c294581871d1e29368d2cc11bb91acdb2232640bf447a95dcc70747e33480bad78f65d62bf15d72e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1459dc7db253b4333fab9bf9e45d96e90c1ecb81fac8af99743e1695a0e66ebbe8d5efaef809e86e097aace90dd9314a0ccd959b8b2bcaf18228fc79a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5eae35387d86115b46fe7d74e7e9f947b0167e7f172ddc2fadef3dd9dadff15d9b7e2aa89b9bf30c21cd4e9945dd76c9ce61ad8c57bb11f195dcd5d32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedd09241d225413e4e7202abfa1dceef6cf68f38ad4e694f01151e045d454a442b4ae96158d6228ea6c0d0fe93d797e7de1ad66b85fdbab83f7d2806c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb3dd9565619fd4390bb977f45b6ad6f75337ec8217db9f5065aedadbda0d7adffc89de5e2a3a8b150a739874b2f2383bb8408bbff26fe55a4f1ee8fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e6c2fa3b15434fa47558dd2ef2cb9c40b6e487355e2c80e4cc4a65ec7d151e666debf24984ede428d005755a00d3791ad3f29497382abf1e481016a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bbfa430e297c40d62e17b13f61e467dae21c176a232bc096744d992f0b182f93f98b58565a3e8d0463d8895a32d10b23734f99b2a5563259fd21e0d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7b03525e40b6c3cdebf0e8cc92c707af31d09c15cbb540a9c1ff20c66df42d21855108ef381bfff810dbbe8f505445f84e44a803f1e4677ae6dd662e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50de05e133ce6d356ea1fb9d4ba90bad4ca14e749b19199571689e2f549b05c8df918768072a4c74ca68e368c06fd5dc6b27e8d0c9df254de5c01f04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a80fbf4e80156cb63cce31d0fb7ac7b29221db95e923dbaa07545763ddafb825232383a7fef3ab4a893820090fe6897f5e003fe7a01af9a9d2bfbb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85c1ffd0c5ce187aa99b5f784d923798ac24e2d44a9fe4e07619f6e98ab65115f3db3c1626d103f3d46b796d1512bafbe21705267991da5e67d5ec91e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbea85a8632cd0f5c13256264ff416c28b05954932c046b52d200506ce8449f1803c24cec16a6b7684477dbc97bc34c34c1a58be608bef490678371b8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70b0cc9c4229828d29da755c10b832c0a80acb4bcd5fce29c97ae67ff5b721aad76a8f51bc69be0a4f6d3f71e2e03de7fda5835b7a34b76df8ea41e90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5d434b01b2040bc5c68385c33d8b4bdad672215e41fda3ea9fdcfece003a11cd468da4e34318c9987b0050a814501245f73a4f7d370bb691148cee18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf27ccc7fe6507ef8dab504f35ac5e612a8cd7c142b9e9a8c6a4e800abf3905b866a0a4d403db4a7f0a1f7629930eb77877eabd39f98b3c3b8d2fe855;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9f3c34f4602c4c6607ed3f99485d4aa97c33adf066d95531a4d0e700ca1ab16e61238b664c179f2cc6a58badcd2513ef5a51b81412c17457e762487b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e2b9350f120a6daead46557c6e2f34add4632bcd0559125310547f682171e4bca2caa6dc3b5a0438d2a67614f79667a28071e5da1ecca40b827df5e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c7a982328f76f0d61327e36c28a01b0d8e16eb853bdc3f92643ddc4f684b82200461f41e2850e0ecfc1e89b7d879d40c8c5f6e1ca900412a53a9dd5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12fc44564d4ae6c31f268dc4c17e7586bde53e5988f83c874e2501132673194a77f0e4b43ffd55c7aace8e853c82372ef7c1393d2a9ad111215b48ecf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70dcb2c2f6b899b9ce27a2bb48c87b32582ea4285a8e230b9be6c23ff37e3fcffd0ff05acc9c9f998e3a6a06f8bceebc8b1cb6880ca2548eb032e717b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55f5d1deb447cce105002a00b0932da2190e0ebb15b214f952532557ad01ba1e687fe564a84bb60b58b002210ceff1c8386126f342888c4e747197bfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60e4c0c47bedb898dcaf1caf5dca80237ad511275a5a2cadc3ef9290b2ad7574552241d9b81e57860ad24d867172d66bd544710e75c371bfa8d9350ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4fd93a33c8c7c27ae0ad7977297b6baca20ca4849b8b43fc0772bda0331169d443fa628773adb7eb04d856977c6186c236b05890e12029c0efe81b80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50963b84b5b1aa82ca5d09d25c7f414520cc230365b101e3e46c596b758e1a425ebb679d1fd14ae3d63223b70731a12750c44ec465abecb6733ce130a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b9921577af251c3a50faa38ab70ef78c58104cadf3dd13f84f36ccce102290fd64c97e1e495e12c707141e6d909496e601e304b29b0b5b19a0e14a66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6feff5b839d79383450e80f9582ca95479a61fe64da2e71b01dab8d828fa361b6181ecb8c774e882d34033562c562bf84fe5da747571e4d5f49dd7c12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a3dae0e862753edd6612bf23695f9a84588877b097f8d0718025a4b81728d05c2b6677265f97d6234abfaf9ffd6db5ddf3aea60d253a2bb8e1ef83d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb0e23205a6e99a1e1f32921cef9d5014af1e455e641de05f0ce9e9525b0e243591e7cce38a4bfe05735d355ad90c0a9de2f0425e1c01433f08c810e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4142ae4c05f4abfaf546d5488361d467a8e351d8c5269d42e8669e54f0e5b6258838c13bd77e6384f2f8a4a1df35f5cb4364430c082b2e606955bf963;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf98385b77dd6a3892accf8a940a290ea77e287bdc072203c10166037b5a1c1073e4017bbd18768b3c267748236b0beba41dc489703fa7ec3d1afc388c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24a08596ba2459d812859cb6058fe70f3b8c3616c578256fe6214866060f44db0b252d42cecfb6a00a665145cf5d15daaddf36e0d5d668bfcff520ea7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he59d991f1b9dfc5955d8601606e174e5ba23ac4c14db66100cbc04e09342d760f3573b2a50c72680b19a575e4a0da4a4ad9b8fb80eb43f9ca88325727;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6423c93dce64719a82096705960785746ef4f8f6ab268807f5ad0b3bf7737b762520efd6bbbe39698a4f13783e72a6a31d62a740f4a5549577a900a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57f8335081f8220225ddb791a9ed4f0a558ad7fbdc41978cd6384f318e1955bb71fb7d190cfad1b2efe79091a3d9979410774a650dec385a6f1ae90d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd98a1c544ed6d8f0cb9dc3731a0ef1c3e125b066160a63efdf363066bfe8d242c3c33ac80831389ec6c31c2cfea191f92d95f4fff039d99bd918cb773;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6a989812eb6d1f33a1a062aad010324e29b2c8ad03ae78150ebce32e0415fbe9ffff09c0f59642baf5f7cb2876b9c081daa8be3e2b8c9bd6f0566996;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3276ee3d6b75ce9f97a2e1de50d290a755c2471273126f4ebc6105ba712837eecd012e9b4cbc1d395e1e1a078d12143ccdd54c2aaea56263b5f9d43d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc76736cba022a540f5883fde103a35d1281b77eba55cc77e11e46be6df7d79587ccf448dad07533db32af79b016bc18c29eba3b8ea041c60a3c103d10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6792040098c65b7f32ce57011edcafd197ef3d023dc5d39a7628d1246d483f40d4119b2a30b6ea17f55f24a531536d277c9552e7d91727cb93e0802ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf54c869a235f2a7c65abf4f57022d431210c96a45f7d5014d3e87892136c6a76d127abae1225152cc98fa0526367ab052acffd10ea650044e19f9867;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f18f85bb6af29055d964cb836e0d8ebce2bf7656c059b41e9684556757e83aeb02134229598acc19e43c4458b4a75f18dba65367418c80d7e7f48501;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4ed4ebbf6652eeb633269e9f21755662829e1043db7bb8980321cc45fb4e3387cfd8a5d2e5a0dd4855619b85bdabcdf98d9b3c8f291030feb022c246;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b36fe5149866111922ed4a60c4690f187e16b31afcbbbe6502bae0cd674ea4aab632469b56dd231d6173349b2312792a1215c7daad21a88578219ae1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd93db985b2c497bd372b0f6d234db6507c0da93299e470096881c7fd50d57f08c15def16c4d0174bf97b73037978dd4fe0ff3eeb7e5575c4c836d8b9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61b8d5edf2effb48a61617114abb3582d469043eeb764abc5e0f8e46172f6622fb462df0a03132613beadfcba2a71361289a5e33ab0a43a28b28f2b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50e04228f7a26fe8aa06bb520851f0caaef084f4fbfab2d6d60baa43ab06b516ed44c12c2a84100afb5923bfddccd5a95f65bce92d4017065b465dc60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c725df5bdc0782e8e94cab035e37c365a80cbdf3ef4df1803746abbe47d1c3aaab1af0c572ca91ed69e9a23d3f28a7cb660242909ced6fb14b13fc1a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4778dfb2af2a3ea716ed342041835655f78126434f75b564020f40680ea2824456970d7aeb435cf54cdee0b70abcba34daff8a59b2e368bf0297f41cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h331eb4c7c77c65e4e0253212764dd6046632fd9a8ae4773e71cc160a608ad15144089e8557e3639295ea7afc330df8ae542c75b2573f589df94352f06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ac853f1070833140258783c44a7d94a94708904b16b695175fbf13c1f87f254634b1454e5a1db8197a87d2c984b7f7c65b0ed2127231e2ea49b4cc62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23e98fd41fadee0f1500acdf6a7da914efbdd12bff44c42039e5dbd4e4bd05c6fb303b84d97800b036eb11a6d1c3fe25506c53415503dc6c46eb45e91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c38d554a3ab7fe9e30fd9b3410643399dd0deeae66aa228d48c47c38edb1ff79ef25aff4fc2efea589d591b99cf8bfbed2dd6fb142940f7607401799;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h489797c5a21a5a0567baec0eee1702e5d2da05e663226f6a37ca521dbedb274d83dbd2f9fa5c378faaf1411d631915436a3d2d7e08f4c22f39a144db0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cd63b5dd457916d503dd72ed128ae9d890a647df1fa96b4f953a15beaf396775b075a4ad8080987cf25966ad4c16ca9a86c24b5dccf5830ca8613fb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h754fc35e20c42a5de115b67294705576feeb84dd0125d7af812af8040310caba5f1ea32a323e1749b6ca8002c7ea6efb0f82b5f5b37a5e3529ec15c45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e8ec791ba8541878ee5bac98070120ac20272e6213a3cb38ecb41cf76f8bbd0b572913c722552b76a2f336db4e59ebdcc25897854b310146c926c4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c9b34aa67f697310ab8e9f0d3b59003b12c75f25717e0ea49714814766ff37cbe4765628720b17cf2782a5e6b21abd6ca45424b83fdaccf390e1be7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47c4343ef841f3f657a75592fa0c4b7fc24bf38a8d9fee4a368996b4f6a43525bb2ef635f735d92c369dffdff7c5f0d039e2e3ef289f481b1be0ead56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4e7c6ac091dcbd5984ea2cbdb7f06bc5b41d794a70364092dd54547fa1b362a74aa87a5c89faa9e0a96f5080b37e14a7bf8815a1f508e562298ad3ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63a0a9de3765c6ed432f49e292b0094766b3e8371e5b7043f240959ee5e22d7dad043e17a0849b241c3833ecd1cd101ff2f333fc20150f192206f1cb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3d106ad6355c9fe82dffd13fe039bd78c2026a232f54623532f0c9d1c1e84beafabd10c213298fa1b2dfdb182d38653bc71ffe2f7ae6536fc4f1772d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf85caf402be9e8b5d69baaf0690600dc580155f19672c05c1545bb48b831bb6d59d766aa3338dd8591c213f6d877a92e63a4d17a39c042f44979b0747;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc79c803648cde90d614d4630947d4dbb869674aea5f55c6767daec3d4f2069b58dfa506784e76e060fd49f096d18736aceb93c257d4c832ec2ae6f9ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50dac8c561eac2df5a6329731d5a4682c85f2f0fd6d9053fd20371635ad44b2530628233d8bedb00454e9daebef0f331120007aecd26095d1a8e3a982;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44e9cb375844c80eab2ee9f017df694edd6aeef882339d7e8c683d2222809832981bdb6060854c4331f69a4606c2b3381d535599639ff4369a2dc80c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fb443fd675cd96822db0040b82100cbebd5b5c17f0f2402fd941721e269576da19e039156e34c23e9ea227cc8b80710d8dc075d5a95109db1896b1bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb31d79921096be014877d71b7998c9eeb774f5225e56a940f720a96366485945ee85501e79a41722832f94954e516833abdc73a8d35b3c96798e21b7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1147fea067e0907af704a382dd0590835bec7080108400212b2119529ef47dceed9aece0a1f876e06249a4b11eb08e0c9e91d143b40c1e1fd6a34d054;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29fadafa723c7371517573f65649f2f2b549a1b11c8d37c6af887a5244281598bfbf9f7039ecf435dfb29d50a4a5f21c282365c5f0bb354e0c9b8ccf9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31abe39fbedc312c2ca004099c827ee3f8d24430b2a392467f43907f1d9c14a48500e56d33c82a9308abf9db6d8975b49e49bd711fa001383530da6bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d52c0d1b9f5807619f19f9706a8552668f0bd129fab7c83bd4da8743489e7390f64107189e0d794f9dbeb667042f0198dcbc69a500996318fd1f9b79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97c1426b4f67c9aea75228cc96dae6fe8d458bab4b8ff71127a6d3fdf936b66e478cd2c5d937c4b6c68f9e9a88defcca1b4ffcbfcdc94f079a8c64995;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30ce74d2368ac62f1ae6e02a1dafe22720145a4a374529e6170ebf14c412834517f3a5ccd621351e7f551a6f618c0a8e7f8fb3685a337dca0760e4209;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d817cb5030259bcaa4aac4e63f30b5f2a03b9bc23f38bbd712e1ac9b8e137bc90b4d15a2826eae7ccf6db909a3cdb732bcb401b9c71a0a4b7df40955;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7937e559aa5b7e2b10fb4a3be6832b59f43b337944d2c809eb86d5e72f26ce663c403ed435215398a5a350ca0bc78d1fbeac542b37e571cb20dc54d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77fcd39c4e2680861770b0b8cc734e0a4aa6332d34e8f72f063ff1b43042cb20d407db5c04ba601847a3173266dc1853d6060eeea6227390bb08d6f12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf639eca5a1da495bb2383f1ba1e72e627aa443ece7521ebf6efffd77d0135834f84e2d6a435c2847aceaa240901fc8682e601a328f6a0a756d4896e1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0973b6d78e374037d997df48adfbb3a52f4db226a7319d6cd0bc47e71770b7df7d31c04b4aea0d9dbeb1534e22d79872c043e4605aa2965f6149f882;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d3404bc699e0965dedc1777e9f51d15486bd0209b20f48ec0878f7b01b2063640fd791a3d4c8c829502d6ab07e8534948b70d67feda3a2858fd432c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h654bc9d26a6670c0e96b64f48a13930e56b4319b98593b7d3ec5cf71dae1df362d1c460a7207a7fa1a1b3a2bda1e1f01f04af2a67c2bc611166c344d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c473cbc26d597d03a8c7b6de271a110b5f83c8ca59c90f8124a33da3b2157dddf51c810e4c860804394357245f3ca7e31f9665d1277572e231d2a429;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8510b45d6938644069febf450953461f9911d9c5b51a0a4dd0c9aa0a71fb2afe61df92debc9ffe3e9707b2191daa219e22c0685538ad41b8fdc052ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27ad0160c45900125524112c3ef08f272f68040c7b27a1317cb905b44ddb4afe8f57242f75aa0066e143b5457e83934f7d8ba4e493ebaf6cf3ea1b573;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h126521a501add295dc0b58123f377d3fdd0ef632ab3dd75a9811d506671083accc571ce71de8f10cc5da7d9e2fabd812a548c42a296714667bb8de760;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1a10f5b8cf606a4bcdc08d0902cfb4c9d5e8b2cc29a09327d89dff84dfa1702c2af2b07c0f04ef719aea629d422c5f31fe4df08844747c382c4be11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52837b1a96ca5a01096d0ace75406acfdd3abd0bc74f924a0d5aacf390fbff3a87a84248664c32e0b5a6296b387ebe072395bc5c3c7dc6b90486edd73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dad8154ef7bb20c3384706c5a22a1b0ddd2edc35e5139e919407f8c8d037ef23884201c4d8353a68c03a9b05535d821639eef19693f4e82360b55a3d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc52db351ba010b34f2afbfa3bf9bac0f21a552aa8da19638154b19ff88c6855468c8431eddc2d6f8fc7c1ad0769ac3e048aaf9c3e7a0fcf1b71c6672d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bd0bf7cc64e6ebc7fc495f4b6c54838a832e13e764e9b7ed2a8f60dcbb26e4fde958ad3d56bd1d5775936c64de7194e70e7d22caa316dfa85eb5f310;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hace38a346a35421ad4281a129bf715d254bf128b201296fd55ea11ff6fd2f17a55a4531a5d201dcb85e8f8fb85cb6b5b500796afd26c56805123747d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5f2c4305f4c65ca2c144496ba723d444ff575b17ebf30674a8218aa2680e24f52b3d47a78d24edce59db9722f877a5b007d9a00c6c3d168a6a07799a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bb544ad30450ebeabb8db221da71c9d9441b76e23070e8686e0fb0808632c111cb645c7da191b4e5d7e06b5038db4904e90ccd96af4c6760733b4fcb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2bc1542ef43679656027b370e6e5e143904082453c128c40992142d51b337b9e30e7b0adbddc983d52905edae63233b4c4c0858e6bc5f209299e366;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4920f9cc6b6ef1ddfbd7458e5fb24f8225d10faffd121f7b0b55254c5d9b2d477464b650eb72d8d27cd750930c8d3f6672a9708587e59a0a2e0543e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he60c04c6a1ee0f6bd572fcc1ef6c1fb8e970b8bf1d5c2a0f7badf284445a89b74cd99ae40533cc85d42168611cfbf684583fc544b250c964e1c45f276;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h624e072fe36f3f7d075d73b5fa9b1880252d787a5ef15dd5eb4c0387c5f8de9375e8bf8458194dcb1711162d2475931f0158e4722238d103e3e4bb880;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6aa0a063d8c5e416cfed8ab22d63a5ea399c9ecf36e7967b85097e8c78283138fcb91bb46f7b0386908b760a7432c941a82889a011c46864361578254;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h432ec0dafdb177821b4b02c3721e32b6446f9cedab3fef7d1cf1a528c3e9bd4222febb5cbf5315dbd05f3032b20df9ff967f1338726b613315ed71648;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7722d17044ec2bbe0f8f40dc153fa031c68d23e20feab89322ca28b8519f81a087016fcf16ebb6cb0def355cb81e23bfb876efa5a33aebc293898f0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h161ab0cb20cbd61b07b5b3cab3c2ad1e8e1fa53833e555d287b763a48898b0b41eb0726ff032e730f94b23d891fc54bf7b673d26e8370d45d34b62ee5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4a64d6c01176c42d7bb13f8b032b9c562b211f942e5969c5beff1e73a4cb904024aab6286d87cc0f786261279c934fa87a2e8cb1db76e143ad04c551;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8d8e8221dc4a97a60ea086f1b0787da523da3b6bb06868bb6f8ef041ac9e5fb33805e9ed70ae98a81ea417d9e7d321a61c4428ef30b97b8c91684a9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55656e1e2947bfd8583ecacda07702c7d520e81ee942d8aa44ced52b33625e66af4e1da8cb8cd539baa48732804e9dbaaaeebcf16443e619dfe29c0b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c86251f820248958f29d09a4f7f4693e864849c792a78e69dd92b868b012cc1a4211a3908e19aec20096a4590a5692f6558a35ebc470d397bb50c7a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94498bcbc3fec70127c639878d1e0c43dc53e01d649e767a3d84d637de22c4ad06705a30a2938b898c1f373249cb6eb1a94c84cc6911c2cdc8d42b85e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ea0641d99c8fd9cff25b3ddb18cb775db2798a49bd7c3dce05987b18ae173efee02e6973771a3b6d0184a7cef4acbf7c40496bccf26089704d14e14b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed19317ef9d4c0eac006a3a773ef6ae57b6f8c586f90e0f653432b6b52dde12119fff51c8708ecf48e01cb5c6a96ab56bbf4d335681a754ec97e78610;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3e0f272f3b9305b6c0628b20da48f93c99a6ba94e5122df9e0f5b01c24892602a5f35f1f1a3adf530a56ac089e70f4e13cec1dc0d5abbf058d1cd5a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h696e077f58bf048c9348bb03f43ad828c9f6a076c0f5de9a820282da8373aa74176c2f46ac2d320592de8657de86cedce8e63d9b9821ef5d53e3a13c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4df0292a9821e9febe74eda06fc8a87ac678cfc51f0b2fe848097b412d26746589372849392c6eedaa893c47dff387ced6efdbe0567aab54fb558be68;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13b06205c67cd9ff4776b5ade8415afd110685dde3bdf8b3aff1f7b96eee851698cbd52ac5c05a0eed2b623a699c3815bd906bfeea691176c7de5b735;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55477c45e7dd25c555a968bdc1b298da99cdfe94e6bb065d17eb6038dd620960d91ea3c527c6142f4db6cf99e4327b6dc9cdbe349d717e7501016d5e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58fbb1ac7e824b496be5f18e19c0e56ee80969b903e2aa3252c8b3c151d6b166786dac4db548cfeb1b92dd7893a1535efacb42b0541cdcaaed1a3c66a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h227bd3beb51d4b4137595d71c042cbbb790e03964ca0167709fd70639703db17ac2ca382fcbf72aad5cc5bd103db705f03995bcb26981d1acd9038596;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h117f70bb30d1c404897c1edf052b536df2e7f27d1668c3b1aefb8c8f30bf6920056d60e442414627966c5ff6e2202cc219a23790dd8f114ed32473365;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc6bd569710358c323e562f2b04479d042914c59b86e0153f93f115b79f4f8b8b3b2f68e68973c00a93740b7cbb03c33b3169857d348cb17f78f0b6fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e1110a23ae77290ec57b18f43f7c734c2d58d0296131388968e0710e04b5cff56a30e629fd19ec389c0db1ed61c4f66b7239c016ef68c72a35c190b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd52f6f8a84981b9abaefaf621e811733da6e69542e82892a369f9ad057bd63219596e1e920f429ed468c869c508ce811e4dab2c63f60b9ea0e93f553e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h830f7250c3e30dddacf1c8be7e731d6b3d25da964a7a5edd568c024cb6ec52706dd3435625d0426460a6134b943633062963395fce9b423fb9853db51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52029c18a60a0ca99998249ab6ca30f96a4a6fef723d2d8ce2674d82ff8d9da83b29a8bb632d624c297ce8d72864419deeb5d25467ba70b8389a42d2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h131212312259ddaed4eea4bb722ae462de7abc8499d3ccad23390a327744c71c36fb8346dab0f3445a278a0d0ab27dd9313dc2175ab2a933ba77c6620;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h982e05b4afce29bc308c382387dc98247ca90c90d7d6d11c87efb8cbf5ffdfa1d1614142fb9b2f19d2e2d2a7cd99d4efac69a31bb0597591be82bd64c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb4deecea8c565cee8eb43b2ad81df4bcfc57bbee783d3a856e213004d1d36c3458abbaa5e69305786b5dc9002893079f29a27044bb460c744d4b9522;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h664c64019ee90030c1d24d9b5bb6cd2e6ada2dbb5276b62e4b0be840c61a7c3419f0f1722809f6732e880d4f3141a978be98765ff949361e71b175dc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8641bcdcce28c88a34cb4d16c6a23dca534c66afa04fc665c280e6fa3896bd160b11f9910bd6a326afd88b49b2e2d6dd6b85022f2565e7c37602765b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66f22c025484fbdadcb61915096c655b3841c54d225071762491bed2cb2893cfd5aa6eeb7c86c9a87d1e2944ceda9e6ca3930e862553a6af807b6fda5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fd59adaa1eac6c90ee162dc9a0c00864977d001dd17480af91dbd440bfca728585043a3a23d663d89dc2298ff72f289a487464865c2b231d6218e824;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf76e7f22ce8da0bdcd5184384e4b16005aad1a0daefe33c35c02e22e8e4eaec62b563eaa65b5b830fd7aa7569b50cd132f41ce3f4bba4686bebca5341;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha387b322211f44b251acfd96ed0f851c17b4b223027ba96a0e231a103aa7bffeeef6c63e41e5b60ab63f7899e9d8278786c43a30e5b7637b128004a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9bc4dac3d12ad4359e2c83ac97614ffaf06962ce151991d44ca65676de11823f6b7deb91564df353a4aecd5c01b5c23af0b3da536f1596070aeea5b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6707c2f5020331ca268240c2a2f2b4ba33fa2bc349d0bb9618e77a1a38a43cfe464792588d15b39ba91fef53d2aaf523c6dc7bda1867fa22629375d4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4843b34b06e66f055a3d051931b895138175ddee03920cac9873d351cd06919c7bd878f532e23144b026ce699cd47472011aa5c562496cdb2d12f76a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0010d80c81630793b7e1e9e217152337fe77a40fed687e018e1e2beecf9c05047d83274c813448a0cb63d2d50d227311b966a08ea3aaf3306247aa0b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd21014bf2ae19a17235215ad3eec220fbb056378212ce171cc778ebcf932a59fde5477a5afa5d2dba763dc37429e0a073612383e4bbbb66c085e42a6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf142169d5decbda65201b8adf2aff2ca92d806b616ad1b90439d7a5583ab84f7cf7804bba9cfac01e2847ed8fcd71e70d78fa17a02c69713a6e7d61f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde9d7e55528246f4933f530d832cfc6c4d8ce35042aaa8ada5f8bc3dd69d65698426f6426e9ff6239963cc2ff40744b1b63e970307a970d8b69dbe4cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb8ddbf5d4efe5bedcf1673eed9fd123856a49afdd533daa0726374214897af5673d9c32b3d455bcf196c6daf311853d4384fbfa725b79ee24f24bc44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13fd2cd8469bb16aa473ef3d1c3f58452f73d3c53e7e7b20bbe3b17eafaca4205545e0ed5d3dc165cd3a64bd9266a2fe0c769f9ee224c9853a008ac07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44090b8f8586d6954f642a0c878f7e8e4498b486dcc2f23fd5235bd3c5ba964789007d13f6865889e4507400d7abe4d9962af9b516389b04a0ab6170b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fc33f4d9ee6cb306792a344392552f940da9b1bb44f2d78be5971d8b1b8807b7523221e0df3e2e4d76a62ef7dcf3e3748246891e3281849a7b024601;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf8d058e569c96c17e2c0c70c24be7a0d2d044c50ee85fdea41e4119efe520a6299ee250b8adba960691dcea4212a278564e567108e627288734cec89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69ef01b61b38d9f6dfada17885bfccb236a69ad44da40252038f81a114e7d3aca73f403f3cc56c3ec85cdeb2a4a409c2713bfd73c86e26eae3a3de67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14b1d3d761e2d1cef1019701e1d3d7abbf9dbf59640142f058395f7f252a9d69e943b21a479a21ac0e86f4b652f5f69618bc288dfff2df5e31b627ee7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb67ff3876b50fbafd23adc41119de4c9d090a50e9826363f8b2d67ec9885add78119ba1ccb68f82041ba2bc01064e97eed6681e60a0872b7266b8c93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80832ec3b3f393be362ed94ec4ed44a11edddb2db656483edda1f45db82fa269009765fba95e41670a7965bc1e9bb95711136e481aefe23806b02a4a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c45dee1d83ebfb57f4b48a27b4d7b81947de1e0774bba3b9ff43dc1e7732f7e74979c21d45dbe7910c7e935e639996f1d56de1def9793c21f6ed1ce2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3d352770706934e5f49e6f102bb0574c25dfbfdbe60e9e97b6c5a5e4ddf7e5d890e064a8f78d3954eb39e93278f9bfe46779367a89b708eebbd7d2b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdea44506172997d3f8987b039b3d6b11e5cef9bb35ec16ca188ab5262ab94811015e1e68063de265f56cc2ea99fbddde4c38c1347a4f605ee7c58fc0a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae6f25e2e35401be795409b74b51a60b13e173f0bf1de6a4d612ed9a8281f9c5f304adcf096ae31ee823b6042281e9da97fe1df93f0b7cd89def50eae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6943caf5cbe10692bf0e2a3d2d81d08cf237ad9e83efcd8b234d0724fc8292186544e4769ab9af214367e0c3afd0c7d3d8dbbdc3e69d7ec26b4737198;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he39290e0de5740d9278e80c98839bd7533edc537fd4fc1b2e42224c9e7fc5d640db8a200bfbf5a097b17829068a5485f42ab2f45ed3f6f3277c50027d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0b98b108a0aa93905d4b5c49502bf76c1ec50bbbdc203ffd49644350bf6cc356a5a845db86111dd1fc9a3d719bd33e592296550c50a23e67bec6a941;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1b37d126ef7b8d63ab7582261950d65ed35ba44de8039643da2b960042ebbc8f5737986b1db893b4c04fca131efdf7a06d11e4b19a4e9a0f40223d48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb603b4d3c7680c474057a5448ce95289a2a49938118a882c8c5312f2de874ace03fcf10f50de426674dade7f7c7b5a2791f7811c9664847a1169ba606;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha917bec67aba48455ea1d65e90d2164102adb703fec243392e69ca84eb13c63b208abf0abb112c2a5c288faf73308d6711167dbc6ce0641ab7380df10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4534a36be97b3bf89f153f0a35d323db52515968958f98630615ed6891a6b006f5933ab64ec06fb7d12b3949b4ef5406f44a2bd87871844e048177345;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d2278ca27a1d3452eaa57acddea21b06c16e0b6bf737cd2e6894335d522da1aac073f3f7dabcf4e6f7e5aa4c1e1500bda9673621232db2c424ac7e32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65f113d471074ea7a370aebe1b75ad403135e561a3fcf4a3889638647ee2796cf19dddba0630b73366411771aea916d066461341a52de4290a4fefb33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3639f5ea6107a44147ad2d2b3066cd301c7d15bd47ca6ef4a32a24c455c34ef29f13221881d8ca8c630b49338a6a0c513ae0c21c408ce0741e47e5390;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc531dfe6756dc496eaca660596ae5174f102630133642f2b0379e73bbe2303ae5c49144953cae0d2083c42782eec21ab272de7a59645892ac17951c23;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83504d2b6aa57e238572c26492acc4d623474e91b4a19cdff7d0a67d99e029411698fc08dd78416a7febd528a50c6475d5c4a9f7caad387b244e6c33e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b52ebc2bb1288801327f1e87ef4989f0718fae3a7866927550f95ec6e1bfa0e31471b5c5adb8d970e4f221c662d5f51ec44661f1aea477539a121df5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4278380ca7386c11ffbc791ed919ccfb2f51cc253eb515c1a7a1c603030d0b04a081aef8aa759246bff59372c404360efb0f39c910e6904dfc4569b2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f93ff052c022a115877bb02bf24e4c4130dac93926cbfc23d8917c915c8bdc177194a3ade1d0eb4752ee8e80a26279ae7f5070f96ae21faf95b751e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had962d98655ed4d74828049c0afdb344b98187893a576e6484e3da8035cb37a5b28ce711c88624f41940a58553f1bbc38de45873c8e80df5c7b93e801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5e10e5db81acb169e3c783147720d36ee5a0d682b1cd6906f141b0f3dbd2fa47c7e2d9802a300b956fda76eea3145d2a372586acdea5f2d72c23d28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1e7c82d5b808f184335cdc487462f1f724a834e82a17edd3c57fb9838cd04f5b54f8fbda7d89bcd62f722413085209f50632f5c01f299607f8788f8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26e38628b9cbee6ee0c73fcef13e460c680955ce3bef8ec55408182ebe877afcfd411a220fba9200cb7f8b6284a8926e95a642bcfc1e105a45e255b9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d4ee4c5b243f92fc39639505a7617bd5724598a72556a978b3ab0dc780ad174b21be13e324f9b5006512d103f5c59ec45db7218af9ef9e4f0f12a482;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69df0d92ca1b439f9b3589c7d0a56b0c38244891ca6026de76298c8c41d16408c9b2744e79c0c1f8a4c01c74092806bb6763a49fab3d98c8e1b54f8b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9b48523eff801d3b615e9696d2a10e61ace90ff43a339e319a5ab6560b4fba52ff32fdc6b1b413b8a2bdafc18c2d14ea17dda6f7c49dc2b53565f982;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8125bf0e75b395e62aeb45b9cecfa97b51b3655781b1c1574794e0d51d0277058bb2caab40f78638dd09c4ba8d1bb44c0c47b2580175f4342c42941bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43eb0cf8424b17cb2e92a2d92c9dbd737dad4b6405e6ba1fc57aa9aabd43fbe5a29cb599783318da9cc74948fdc052ee3215d137b61a713ed5cff3c67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd14c9f3cf6f87c63904893d4c58a21ac90bc60dc83fb51687bbeea90fc486d72760662ac8fae7e610307227f8321436124380547e435503285077a285;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a9a6280842309aead2cb560a3a8b2313d58ae356c64f21ec30b023bf767162be0528cba0ee52df883f72cf1ecfe754ea10d06df01fa8f64062b5be6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h303fe4719c22e91323c9a38bfe5ff500fa8df6390bd8806a0f8233c20e0072471b38653d9a4c057bbab5762376b166640a447b8c31879098a03d5a460;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3776abce0543084f8fcf597b2e1ad66de42da525592e63de17ab123eb70f22010c960d638af1a29ba50aad97485cc8eb65473553e9a892a0230a9c610;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d63f9defc425481567a9984893f040eb396b8bee1d8c11a5510756c49846ba6163b46125e4e60318a3fa6ec12f78a7641e479a0d824fde7d2fab6c2a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8248878784d65eac74e63b909ca000eb168d58c86fbe5e27e072f098e547a6d17ccb2e8f0dba96372e2853fbf0ddb88d4403216a287394692ea821ba1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64627288bd57c8198d9a4c8cc513fab4542e2f60852f036095652e63bde78a5d5a63644abbb77eeb459dc10c1477cbebc86a4d32fa98e0338d70a801a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9fdcf8fda5f93e3dbe644b3729fbeeebb497a99cafb138e25ed503d106b6efffc470fdb31dd4201a0ed45dd55480cb4db41d544f40200479d2e71b43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8db494e9bf74a1bf894bfd6d87e2a176ba4cf68a0bfe159273cfeb6892d92182c1dbda903ba77f8ef9392930225afab75186ccf2ac0596ad5986afcc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafc264e71b2bc38fbbac3cc4cf982fc62cf4d590be64ee0391fe888e30ae8856198ec6c3f3dc8654bc06f7a37019c99eccc082c646c9178cff154741;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1b45a13101ef8b9202bbd1ebed8479bacacc222a080a7e7db3ae39a1bcbf1a9e32f4f8e26b9fa4d10afd087285cb3173abb4aa803c8db961af35a740;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had96638cd5bb78fbd29527017ab1378cdeae313085eb297d605a1c78ce47b0a6e1c7cabd4287c2086a6a63a970080fff28836075c9a7d233d94c1a130;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha36a896beb3a77a706a22410b2e5bf09946a12b709838f0dc1a746b66e4a372507e5abe2461fadf4044863f18d3763785d81564981012eba713e1b650;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48b489331458b6da1490c8c2f2c56bddf33ecd295acf40bb4c6882b40c2a33db6f458f31c21aa65e10106aa879e63acc993e554f2785c462b2000b371;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf78eefa9a05aad7e137baf2b49f146db427a30fb00865401c55a53b43c3e00b3e07b7304c861763630f41678151151bf4d066383ccb7486f1936caa3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf425069dc293511f7d9df2a4edb81b8ad1d46fd1c58cf525ad21d3deaf9a0fdae462b3b8085873c59e2482bb465830ebf2e5d56a2607be2e46e8f35da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc587c88a937e25927f7c79bd64d421053cf6325f02387f28ac690d7dd254662425ef25d9e20c9766e1c8589bf1a9a4822eccc34083a1cb7326650f397;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3945f9a248cd121d822b5d6541c37de285a247638d286bff99e577bf20ade3ace0ea624074acdc2c0935e72e2927fa3bcea84958ac94832dacd208753;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb33023f9c2c1ea57494ce5a605922cda14e3b466b571880af6e29fb053357159a53f9ccf67c0e87c67041dcaad6022ae5b4813b97376f90e82aeb5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3530a7d18801ac49a8f884ba1aa81db7d863bd864580ad7cb83b4d124d905656d8ce564bfe2a07adebd114474a594d86911b567a41b4fb484a04ab49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd82b50be79e6f5d36f2eb8cac5898eb1115b69b05c583755df87aa732f441c1aead9c2f3c7a6d219adc6f23fbd7d52d950cd3e76ac7c2bb8f423534b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ab1b142893446f09874077ea1277ef1fa5be9c11c285dccd76aff6b0ceada7a9adcf25578f88c7520fbbc67572c35ac8297a30628f8d25562d10bb49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98fc5cb535889ade160d670a3a9c1ca5254e668bf4d7605c5aa3bcdad1d3bc673719906e7de2198206e4f1db4db3f85e2415104bd7a71b49006042602;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14a2fa8606cb190ddd62f13e01bc4c13996142fe6846c1fcb8c3387eb667f256361893597842e41087b7d2034b2a3171382e27eac1f70273553ef41a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde04fe35a81c48445f4e159e0f08bcb21d9b4492df0d44aed374465aa3171e5b43683dc26f241dffa0c69506de68bf4dec7606a4f6a2a10a5c770b451;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha39d48266c45e4e2f0a3d4cdc83d1f3dc2b256ec897eae87219dddaec4b7cd7fdf2fedd2daf628b602358590e3b2d1994448b289d9d2067e57a58fad4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha82be420463efddd10a4b604ba0b40b906b85a04c11356cdb1dbdf4e5d250d05b765ab0b55db974cabee45bfce3eebd9cb3aa84f4b0410eb5f087212e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf520399b8b28fc0f0de77152d592d596b528d49d8f0cb0356bb9ab1b087840068cb822d3c9c180645e7dd1db2ae976c92ec3e49ea8c54455cff090c22;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haeaa1e1d58aba7df843247c558a0283facda98b87ab2b4f4e84e312f4b718f7dd730036283f3b6df3972dce5341806146d103b7d5888bd9b3cc6e4196;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43f497ba516492899b5a941ba78987d4fe5d969ffcb999b2bf275f0e7f46fd8a7aa42b39e21e502a704ae5e319c63523691bf7136f5d66ee4d9e5e567;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebd259c39c927ba0a0b3e39f61eb0b77fc9ef879ed0dbc821d4f48aeabe2f73c7deadea260e1c1eb5733207ef36eecc2902c692a4a883e435b87592a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb54b5ad697af4ac256d4019011d31c762441c6b43cddd847c85a0d395179ae08a385fbf19efc79347ffa4da7b749400b1f53f45e556220277fcb7cb96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3d32b483256bdec4a42a4f0c8e76ddd1b87a826247b9e3b4baf771e9f6e43f2862c2092fcd5610f5998f5876a009a214beb0d2b2da5d339723f4459;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2570e126d99d9b9b105c133596581076aeb585a286353a5279a76334a22968ae975d73fc858557593a6c545f5666d3b0d7ff5a75a256dd0b67782503;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha07089ed39703ca380232ddea6d1697fbca71b909b97ec0bac264a2d38a859dc517f896589738df1082fbae77efa729c29415eca651433a4f341de825;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2970a2dcf4fd28cb5230179f0a090f6c45d4ecc2ea07008ed88ad5c4a1e316e15bfa2ab38dd95bf886344e92f123a72ff204af0338a8f25408f1a08a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9743e71afbc9828d4022c04d72d34854cbf04abb55685c44cdb343288df01bbeeb107a1235d299233508861a64c450c94502597459969466886c7776;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1574f1a1206c0375ea5d460fc8961afd9215655e0033b2878a5c661e8c51112dbfb14fa56615d03f337ddf275033fb3caae8dafa0f50f12d1193b1e63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h240aab75e4500afebf0ff1f0c12a8699dce4d44e13fc28c94b506296c1306e2b6f4f0bb0b2be6f68cd216c65c53b8fe4877ca0fa58fff4d4e53093a2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c427e4cca1881ae06a4e2a2bc1e3785b0ac12fa9a9b2edd8c7ab7e4341316c8b0869ad6d03371196a57ef13c208c5558eb6a31ddbb7d3edfb96ad7d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecf3e4d9ab8d9fc9c833b1938156b25f88bb388aba45aa5c5d9988a4b2aeb9f082963120cd8f48388b8fc3d8269b9b4348508a143281163fb77a1e3b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h458b22020c3641621492d9250d422f874d1260b0be0bc80fc4d6f7e3311f07c801a161a8d036b41750554d76aeb3b9c397ae7de48694ae2360d7620bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81bd9c49da34ec3336d85a0f182556c8940bdc0c14d2bb4d4c4697d22ff031f3195cb00328dd83f128f33a2b2557ce2d70962e920552a13a257aeb7dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5b1c5399589ebdba494b1c77c162ba55799921ac263e43ad641e79ab7194a5153b7d69fcd0006470d4c9c4fa64d657d43991f1287585fb39195b8fc6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f0929148115dee620882590af89ee557df5e60950d1180de22b5c084ac6d3e14f96e7206ea36aac7af227806b7bb692fc8c31e8794e978accc00c9e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc45ef64ce2e6f17cc7a8ad02b7d6862b149f515a5673f77c72a6798c4c602a5af3370a250eb0625849f2a2fa6d133149a1b988e057199e859609333b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a5b28bca4c367c4e4f4099597511f76da7e4d5605635f42167d343162939349f44edd5aab1d8c159dc7ddfd74481955da3a13ae6f24ecc817b381552;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2894dfb7161f51a3ffde289b61f82c13cb574e1b16640435382c7b7d02589704fdb0930fe6b41edc66225c06e1832b5b8be53c43402b6b22bd2287eb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb72cb12fa691a7bfc5cc6a07d8ef8f0a52366adc031230ac3e57ec91f9682eab88fd3285e05c99a85d64d5507ade1aa08cffd8df8e5f18c09b6a89d0b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8144abf1e27080ade9d7535bffe4dd3dc647145ca23e32e179501ecba0852354e464e8269a5bd4dd509797dbd64d02475cec02f29715ec0b928e7782;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29411a10c50a80de268eaec529a35438ca2a243e5ef948090eba3136a9409624748443b4d556a86769dde47cc4d4e2663f49b44b1f1ba474a6567860;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a32ccd1d218a9ba2191afe8548a2191e68209125c8f51ce4e97ae14ecfc9d79c16947c896a117a19788c3faff2ce299801cb808807e8756291b00336;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefda33e4f30eda0bddbda6e9cad8eb7e0bb8963caebeeb4fa5ddc231c7d8c4681f40681820ad5a66ba8b1ef8676982ad1a35673e2a479a3eaa952f5f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69aa4dddf8d882f6749ee18652d2aa6be3e018089cf031a2970bf9953d47e925f5fbaa223ae1975589a35e819cdd9212bebf1bd8ff0eaf808952dc733;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4ec60153106c55c3263a08743e38826702e3c301e83c5df3b3b45d1fad3860479c2a5ec12379ca950fd25209455a13e8c7c0c99048a45f6fdc29ced0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41e4e7c881eafad79d0a0ca4b39005df6f0356b950b2e43324ffe3d6bcd1adf76a90136eaf88267a301acd82d57eed652134da814a2255202e9d939df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a22c566126a25a0bf1d11d42ca892cf6a3720be612a0cbc2f1f43ffef8ce46686411909498345ec34e04be4d86022c4fc518e02135624e9f4d8fe48b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h429cb80f74ca855642eb0cf10971f154d2dd66d137e7fa03d7a0a246627858919cab7956b845df5f6d0847c3fb0da578eb0afe6e0e2186dfe400f86b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha942ba8e1fa8120d63cb5c49f2b1f160342ab9ff70b6f34c8b69f9c329e2fd2d511485a66b0a66dc9644abb32803711d14a2104ee48ed61ef0637b33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd3585b6287baac9a86fbc220b26879998fa89d36f569aa386f3fe42fc1b09c757a2081a6b7e46a33e21cb879ad3360011d8d183a99daccfad205b782;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h710147218d97b9ba6cebb00f6cc73564ed24e9962efa0eddd51768e0874ae8d4d36895ae65d738d4ae8ff3b3e2356eeea77c968684b37d5553fc7e3a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98f7b1f9524c5639f41c542d58030084fb06d5793b80ba38973d073f5d8528e45f1cc1959e97d311e45944aa7a36267d9ffa90594cde68911645bb1eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a981781224a6e8aff4b606e62b155a0cb072a25925eb75950c129858762e9a0953adf468fc392d3f04ace2c89276c4e38252d12e384797a370b2051c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84eeb0ee52fd2e529eac97e0e82a3559b08ce6793ca3c976d6456456d9097aea3ef2f3bafa3d6d023fd85c3db14d33591b057acf22c8d2c7886a687f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b7dd5d37150dd4629f173b8399186370170c597761994dea7f55cfb1b28f2e46c949bcdcb96fc1d845088ae2c5d1a5f5f311d055fa9a6897be70b8d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc99fdb17e3a66684e227c0b57bca14dd9d2eb5ebd873f9cfa8856dd27014fa7f9700159e3d86c83a2deb36d9f8c83c0840f31f904835226a7974d2c83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfb08bbd37295bc0eb3c4a052f151746bde3f1f0d2a6fdfb9040fafd5f8c9f1da4dde134e6b27d10e702ab39b2626025cf84c29058723377a58320269;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had013b4d670d18ddf0712f57b3249a272cc3c38a1a5c045e940a93835104927e637fabfb0a997d4378c0003773248bfda4d8ec7de9eabdd0ce00e9844;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3479c74ad54df7cac7e8fa36559a129f4d2b4cce8a907374bf2f0ea7277d188074609a7a64afa4f3321069517d142c28f903caa21e4b149d644c66824;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc04861fe534f60e8f270760711be85c1b9bd19473564630fadb05a1bfd5c30ceb855ee1e62b3a09bff5160fc5431ca13d0bc6ef9236a8a90f9c7c2799;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20d8833932100db21114575393e2282a1232beda151e96eae893a9f4dcadc69703d403f6dc3e5a83a0502779afd65a9a06fff65d6930c49a5710c58e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fd5f6bd978ef8ebc97dc20227d932642b87e1e71a1653fff638762a7b2054b576805930872fbc97875ad9961f664fe6ad43ccc7c6210873845dab414;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcfc674f87d10d79d448bd51aae1ef68f88e3c36211ac27fa3f62b5ef5b26dd3a30ef650cca6e65623d3a29af367c58f005ef1a1915b17372a62ce5fe;
        #1
        $finish();
    end
endmodule
