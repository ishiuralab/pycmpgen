module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    compressor_CLA32_32 compressor_CLA32_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
        src16 <= 32'h0;
        src17 <= 32'h0;
        src18 <= 32'h0;
        src19 <= 32'h0;
        src20 <= 32'h0;
        src21 <= 32'h0;
        src22 <= 32'h0;
        src23 <= 32'h0;
        src24 <= 32'h0;
        src25 <= 32'h0;
        src26 <= 32'h0;
        src27 <= 32'h0;
        src28 <= 32'h0;
        src29 <= 32'h0;
        src30 <= 32'h0;
        src31 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA32_32(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    input [31:0]src16,
    input [31:0]src17,
    input [31:0]src18,
    input [31:0]src19,
    input [31:0]src20,
    input [31:0]src21,
    input [31:0]src22,
    input [31:0]src23,
    input [31:0]src24,
    input [31:0]src25,
    input [31:0]src26,
    input [31:0]src27,
    input [31:0]src28,
    input [31:0]src29,
    input [31:0]src30,
    input [31:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [0:0] comp_out33;
    wire [0:0] comp_out34;
    wire [0:0] comp_out35;
    wire [1:0] comp_out36;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[1], 1'h0, 1'h0, 1'h0, comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [0:0] dst33,
      output wire [0:0] dst34,
      output wire [0:0] dst35,
      output wire [1:0] dst36);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [31:0] stage0_16;
   wire [31:0] stage0_17;
   wire [31:0] stage0_18;
   wire [31:0] stage0_19;
   wire [31:0] stage0_20;
   wire [31:0] stage0_21;
   wire [31:0] stage0_22;
   wire [31:0] stage0_23;
   wire [31:0] stage0_24;
   wire [31:0] stage0_25;
   wire [31:0] stage0_26;
   wire [31:0] stage0_27;
   wire [31:0] stage0_28;
   wire [31:0] stage0_29;
   wire [31:0] stage0_30;
   wire [31:0] stage0_31;
   wire [10:0] stage1_0;
   wire [14:0] stage1_1;
   wire [11:0] stage1_2;
   wire [12:0] stage1_3;
   wire [18:0] stage1_4;
   wire [11:0] stage1_5;
   wire [12:0] stage1_6;
   wire [20:0] stage1_7;
   wire [11:0] stage1_8;
   wire [17:0] stage1_9;
   wire [11:0] stage1_10;
   wire [15:0] stage1_11;
   wire [12:0] stage1_12;
   wire [14:0] stage1_13;
   wire [12:0] stage1_14;
   wire [17:0] stage1_15;
   wire [12:0] stage1_16;
   wire [18:0] stage1_17;
   wire [16:0] stage1_18;
   wire [11:0] stage1_19;
   wire [12:0] stage1_20;
   wire [14:0] stage1_21;
   wire [11:0] stage1_22;
   wire [13:0] stage1_23;
   wire [22:0] stage1_24;
   wire [14:0] stage1_25;
   wire [11:0] stage1_26;
   wire [15:0] stage1_27;
   wire [16:0] stage1_28;
   wire [13:0] stage1_29;
   wire [22:0] stage1_30;
   wire [9:0] stage1_31;
   wire [7:0] stage1_32;
   wire [4:0] stage1_33;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [3:0] stage2_2;
   wire [4:0] stage2_3;
   wire [10:0] stage2_4;
   wire [5:0] stage2_5;
   wire [3:0] stage2_6;
   wire [5:0] stage2_7;
   wire [7:0] stage2_8;
   wire [12:0] stage2_9;
   wire [3:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [9:0] stage2_14;
   wire [5:0] stage2_15;
   wire [7:0] stage2_16;
   wire [5:0] stage2_17;
   wire [5:0] stage2_18;
   wire [10:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [5:0] stage2_22;
   wire [3:0] stage2_23;
   wire [8:0] stage2_24;
   wire [7:0] stage2_25;
   wire [5:0] stage2_26;
   wire [8:0] stage2_27;
   wire [7:0] stage2_28;
   wire [5:0] stage2_29;
   wire [5:0] stage2_30;
   wire [6:0] stage2_31;
   wire [6:0] stage2_32;
   wire [2:0] stage2_33;
   wire [1:0] stage2_34;
   wire [0:0] stage2_35;
   wire [1:0] stage3_0;
   wire [0:0] stage3_1;
   wire [1:0] stage3_2;
   wire [3:0] stage3_3;
   wire [6:0] stage3_4;
   wire [1:0] stage3_5;
   wire [5:0] stage3_6;
   wire [0:0] stage3_7;
   wire [6:0] stage3_8;
   wire [4:0] stage3_9;
   wire [2:0] stage3_10;
   wire [1:0] stage3_11;
   wire [6:0] stage3_12;
   wire [5:0] stage3_13;
   wire [1:0] stage3_14;
   wire [5:0] stage3_15;
   wire [2:0] stage3_16;
   wire [5:0] stage3_17;
   wire [1:0] stage3_18;
   wire [2:0] stage3_19;
   wire [5:0] stage3_20;
   wire [3:0] stage3_21;
   wire [2:0] stage3_22;
   wire [3:0] stage3_23;
   wire [5:0] stage3_24;
   wire [2:0] stage3_25;
   wire [1:0] stage3_26;
   wire [4:0] stage3_27;
   wire [5:0] stage3_28;
   wire [6:0] stage3_29;
   wire [0:0] stage3_30;
   wire [1:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [2:0] stage3_34;
   wire [0:0] stage3_35;
   wire [0:0] stage3_36;
   wire [1:0] stage4_0;
   wire [0:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [0:0] stage4_35;
   wire [1:0] stage4_36;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;

   gpc1406_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[4]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[5]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[6]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9]},
      {stage1_5[0],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc615_5 gpc7 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[7],stage1_3[7],stage1_2[7]}
   );
   gpc615_5 gpc8 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage0_3[11]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[2],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[3],stage1_4[9],stage1_3[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[4],stage1_4[10],stage1_3[10]}
   );
   gpc615_5 gpc11 (
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[5],stage1_4[11],stage1_3[11]}
   );
   gpc615_5 gpc12 (
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage0_4[15]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[5],stage1_5[6],stage1_4[12],stage1_3[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[4],stage1_6[6],stage1_5[7],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[5],stage1_6[7],stage1_5[8],stage1_4[14]}
   );
   gpc606_5 gpc15 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[2],stage1_7[6],stage1_6[8],stage1_5[9]}
   );
   gpc135_4 gpc16 (
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16]},
      {stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage0_8[0]},
      {stage1_9[1],stage1_8[3],stage1_7[7],stage1_6[9]}
   );
   gpc135_4 gpc17 (
      {stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21]},
      {stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage0_8[1]},
      {stage1_9[2],stage1_8[4],stage1_7[8],stage1_6[10]}
   );
   gpc135_4 gpc18 (
      {stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage0_8[2]},
      {stage1_9[3],stage1_8[5],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc19 (
      {stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30], stage0_6[31]},
      {stage0_7[15]},
      {stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8]},
      {stage1_10[0],stage1_9[4],stage1_8[6],stage1_7[10],stage1_6[12]}
   );
   gpc1343_5 gpc20 (
      {stage0_7[16], stage0_7[17], stage0_7[18]},
      {stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[7],stage1_7[11]}
   );
   gpc615_5 gpc21 (
      {stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage0_8[13]},
      {stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[8],stage1_7[12]}
   );
   gpc606_5 gpc22 (
      {stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[0],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[9]}
   );
   gpc606_5 gpc23 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[1],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[10]}
   );
   gpc606_5 gpc24 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[2],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[11]}
   );
   gpc606_5 gpc25 (
      {stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[3],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc606_5 gpc26 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[4],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc606_5 gpc27 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[5],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc606_5 gpc28 (
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[6],stage1_11[8],stage1_10[9]}
   );
   gpc606_5 gpc29 (
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[7],stage1_11[9],stage1_10[10]}
   );
   gpc615_5 gpc30 (
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[5],stage1_12[8],stage1_11[10]}
   );
   gpc615_5 gpc31 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[6],stage1_12[9],stage1_11[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[2],stage1_14[4],stage1_13[7],stage1_12[10]}
   );
   gpc606_5 gpc33 (
      {stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[3],stage1_14[5],stage1_13[8],stage1_12[11]}
   );
   gpc606_5 gpc34 (
      {stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[4],stage1_14[6],stage1_13[9],stage1_12[12]}
   );
   gpc606_5 gpc35 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[5],stage1_14[7],stage1_13[10]}
   );
   gpc606_5 gpc36 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[6],stage1_14[8],stage1_13[11]}
   );
   gpc606_5 gpc37 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[5],stage1_15[7],stage1_14[9],stage1_13[12]}
   );
   gpc615_5 gpc38 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22]},
      {stage0_15[18]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[6],stage1_15[8],stage1_14[10]}
   );
   gpc615_5 gpc39 (
      {stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage0_15[19]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[7],stage1_15[9],stage1_14[11]}
   );
   gpc615_5 gpc40 (
      {stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31], 1'b0},
      {stage0_15[20]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[5],stage1_16[8],stage1_15[10],stage1_14[12]}
   );
   gpc615_5 gpc41 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[6],stage1_16[9],stage1_15[11]}
   );
   gpc606_5 gpc42 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[1],stage1_18[4],stage1_17[7],stage1_16[10]}
   );
   gpc606_5 gpc43 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[2],stage1_18[5],stage1_17[8],stage1_16[11]}
   );
   gpc615_5 gpc44 (
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10]},
      {stage0_18[12]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[2],stage1_19[3],stage1_18[6],stage1_17[9]}
   );
   gpc615_5 gpc45 (
      {stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_18[13]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[3],stage1_19[4],stage1_18[7],stage1_17[10]}
   );
   gpc615_5 gpc46 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage0_18[14]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[4],stage1_19[5],stage1_18[8],stage1_17[11]}
   );
   gpc615_5 gpc47 (
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25]},
      {stage0_18[15]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[5],stage1_19[6],stage1_18[9],stage1_17[12]}
   );
   gpc606_5 gpc48 (
      {stage0_18[16], stage0_18[17], stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[4],stage1_20[6],stage1_19[7],stage1_18[10]}
   );
   gpc615_5 gpc49 (
      {stage0_18[22], stage0_18[23], stage0_18[24], stage0_18[25], stage0_18[26]},
      {stage0_19[24]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[5],stage1_20[7],stage1_19[8],stage1_18[11]}
   );
   gpc615_5 gpc50 (
      {stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[6],stage1_20[8],stage1_19[9]}
   );
   gpc615_5 gpc51 (
      {stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage0_21[6]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[1],stage1_22[3],stage1_21[7],stage1_20[9]}
   );
   gpc615_5 gpc52 (
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22]},
      {stage0_21[7]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[2],stage1_22[4],stage1_21[8],stage1_20[10]}
   );
   gpc615_5 gpc53 (
      {stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_21[8]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[3],stage1_22[5],stage1_21[9],stage1_20[11]}
   );
   gpc615_5 gpc54 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], 1'b0},
      {stage0_21[9]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[4],stage1_22[6],stage1_21[10],stage1_20[12]}
   );
   gpc606_5 gpc55 (
      {stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[4],stage1_23[5],stage1_22[7],stage1_21[11]}
   );
   gpc606_5 gpc56 (
      {stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[5],stage1_23[6],stage1_22[8],stage1_21[12]}
   );
   gpc615_5 gpc57 (
      {stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_22[24]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[6],stage1_23[7],stage1_22[9],stage1_21[13]}
   );
   gpc615_5 gpc58 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage0_22[25]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[7],stage1_23[8],stage1_22[10],stage1_21[14]}
   );
   gpc606_5 gpc59 (
      {stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[4],stage1_24[8],stage1_23[9],stage1_22[11]}
   );
   gpc615_5 gpc60 (
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28]},
      {stage0_24[6]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[5],stage1_24[9],stage1_23[10]}
   );
   gpc615_5 gpc61 (
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_25[6]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[6],stage1_24[10]}
   );
   gpc615_5 gpc62 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16]},
      {stage0_25[7]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[7],stage1_24[11]}
   );
   gpc615_5 gpc63 (
      {stage0_24[17], stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21]},
      {stage0_25[8]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[8],stage1_24[12]}
   );
   gpc606_5 gpc64 (
      {stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13], stage0_25[14]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[3],stage1_27[4],stage1_26[5],stage1_25[9]}
   );
   gpc615_5 gpc65 (
      {stage0_25[15], stage0_25[16], stage0_25[17], stage0_25[18], stage0_25[19]},
      {stage0_26[18]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[4],stage1_27[5],stage1_26[6],stage1_25[10]}
   );
   gpc615_5 gpc66 (
      {stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23], stage0_25[24]},
      {stage0_26[19]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[5],stage1_27[6],stage1_26[7],stage1_25[11]}
   );
   gpc615_5 gpc67 (
      {stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_26[20]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[6],stage1_27[7],stage1_26[8],stage1_25[12]}
   );
   gpc615_5 gpc68 (
      {stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24], stage0_26[25]},
      {stage0_27[24]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[4],stage1_28[7],stage1_27[8],stage1_26[9]}
   );
   gpc615_5 gpc69 (
      {stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29], stage0_26[30]},
      {stage0_27[25]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[5],stage1_28[8],stage1_27[9],stage1_26[10]}
   );
   gpc615_5 gpc70 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16]},
      {stage0_29[0]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[0],stage1_30[2],stage1_29[6],stage1_28[9]}
   );
   gpc615_5 gpc71 (
      {stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage0_29[1]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[1],stage1_30[3],stage1_29[7],stage1_28[10]}
   );
   gpc615_5 gpc72 (
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26]},
      {stage0_29[2]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[2],stage1_30[4],stage1_29[8],stage1_28[11]}
   );
   gpc606_5 gpc73 (
      {stage0_29[3], stage0_29[4], stage0_29[5], stage0_29[6], stage0_29[7], stage0_29[8]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[3],stage1_30[5],stage1_29[9]}
   );
   gpc606_5 gpc74 (
      {stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13], stage0_29[14]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[4],stage1_30[6],stage1_29[10]}
   );
   gpc606_5 gpc75 (
      {stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19], stage0_29[20]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[5],stage1_30[7],stage1_29[11]}
   );
   gpc606_5 gpc76 (
      {stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[6],stage1_30[8],stage1_29[12]}
   );
   gpc615_5 gpc77 (
      {stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_30[18]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[7],stage1_31[7],stage1_30[9],stage1_29[13]}
   );
   gpc1_1 gpc78 (
      {stage0_0[27]},
      {stage1_0[6]}
   );
   gpc1_1 gpc79 (
      {stage0_0[28]},
      {stage1_0[7]}
   );
   gpc1_1 gpc80 (
      {stage0_0[29]},
      {stage1_0[8]}
   );
   gpc1_1 gpc81 (
      {stage0_0[30]},
      {stage1_0[9]}
   );
   gpc1_1 gpc82 (
      {stage0_0[31]},
      {stage1_0[10]}
   );
   gpc1_1 gpc83 (
      {stage0_1[24]},
      {stage1_1[7]}
   );
   gpc1_1 gpc84 (
      {stage0_1[25]},
      {stage1_1[8]}
   );
   gpc1_1 gpc85 (
      {stage0_1[26]},
      {stage1_1[9]}
   );
   gpc1_1 gpc86 (
      {stage0_1[27]},
      {stage1_1[10]}
   );
   gpc1_1 gpc87 (
      {stage0_1[28]},
      {stage1_1[11]}
   );
   gpc1_1 gpc88 (
      {stage0_1[29]},
      {stage1_1[12]}
   );
   gpc1_1 gpc89 (
      {stage0_1[30]},
      {stage1_1[13]}
   );
   gpc1_1 gpc90 (
      {stage0_1[31]},
      {stage1_1[14]}
   );
   gpc1_1 gpc91 (
      {stage0_2[29]},
      {stage1_2[9]}
   );
   gpc1_1 gpc92 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc93 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc94 (
      {stage0_4[28]},
      {stage1_4[15]}
   );
   gpc1_1 gpc95 (
      {stage0_4[29]},
      {stage1_4[16]}
   );
   gpc1_1 gpc96 (
      {stage0_4[30]},
      {stage1_4[17]}
   );
   gpc1_1 gpc97 (
      {stage0_4[31]},
      {stage1_4[18]}
   );
   gpc1_1 gpc98 (
      {stage0_5[30]},
      {stage1_5[10]}
   );
   gpc1_1 gpc99 (
      {stage0_5[31]},
      {stage1_5[11]}
   );
   gpc1_1 gpc100 (
      {stage0_7[24]},
      {stage1_7[13]}
   );
   gpc1_1 gpc101 (
      {stage0_7[25]},
      {stage1_7[14]}
   );
   gpc1_1 gpc102 (
      {stage0_7[26]},
      {stage1_7[15]}
   );
   gpc1_1 gpc103 (
      {stage0_7[27]},
      {stage1_7[16]}
   );
   gpc1_1 gpc104 (
      {stage0_7[28]},
      {stage1_7[17]}
   );
   gpc1_1 gpc105 (
      {stage0_7[29]},
      {stage1_7[18]}
   );
   gpc1_1 gpc106 (
      {stage0_7[30]},
      {stage1_7[19]}
   );
   gpc1_1 gpc107 (
      {stage0_7[31]},
      {stage1_7[20]}
   );
   gpc1_1 gpc108 (
      {stage0_9[27]},
      {stage1_9[13]}
   );
   gpc1_1 gpc109 (
      {stage0_9[28]},
      {stage1_9[14]}
   );
   gpc1_1 gpc110 (
      {stage0_9[29]},
      {stage1_9[15]}
   );
   gpc1_1 gpc111 (
      {stage0_9[30]},
      {stage1_9[16]}
   );
   gpc1_1 gpc112 (
      {stage0_9[31]},
      {stage1_9[17]}
   );
   gpc1_1 gpc113 (
      {stage0_10[31]},
      {stage1_10[11]}
   );
   gpc1_1 gpc114 (
      {stage0_11[28]},
      {stage1_11[12]}
   );
   gpc1_1 gpc115 (
      {stage0_11[29]},
      {stage1_11[13]}
   );
   gpc1_1 gpc116 (
      {stage0_11[30]},
      {stage1_11[14]}
   );
   gpc1_1 gpc117 (
      {stage0_11[31]},
      {stage1_11[15]}
   );
   gpc1_1 gpc118 (
      {stage0_13[30]},
      {stage1_13[13]}
   );
   gpc1_1 gpc119 (
      {stage0_13[31]},
      {stage1_13[14]}
   );
   gpc1_1 gpc120 (
      {stage0_15[26]},
      {stage1_15[12]}
   );
   gpc1_1 gpc121 (
      {stage0_15[27]},
      {stage1_15[13]}
   );
   gpc1_1 gpc122 (
      {stage0_15[28]},
      {stage1_15[14]}
   );
   gpc1_1 gpc123 (
      {stage0_15[29]},
      {stage1_15[15]}
   );
   gpc1_1 gpc124 (
      {stage0_15[30]},
      {stage1_15[16]}
   );
   gpc1_1 gpc125 (
      {stage0_15[31]},
      {stage1_15[17]}
   );
   gpc1_1 gpc126 (
      {stage0_16[31]},
      {stage1_16[12]}
   );
   gpc1_1 gpc127 (
      {stage0_17[26]},
      {stage1_17[13]}
   );
   gpc1_1 gpc128 (
      {stage0_17[27]},
      {stage1_17[14]}
   );
   gpc1_1 gpc129 (
      {stage0_17[28]},
      {stage1_17[15]}
   );
   gpc1_1 gpc130 (
      {stage0_17[29]},
      {stage1_17[16]}
   );
   gpc1_1 gpc131 (
      {stage0_17[30]},
      {stage1_17[17]}
   );
   gpc1_1 gpc132 (
      {stage0_17[31]},
      {stage1_17[18]}
   );
   gpc1_1 gpc133 (
      {stage0_18[27]},
      {stage1_18[12]}
   );
   gpc1_1 gpc134 (
      {stage0_18[28]},
      {stage1_18[13]}
   );
   gpc1_1 gpc135 (
      {stage0_18[29]},
      {stage1_18[14]}
   );
   gpc1_1 gpc136 (
      {stage0_18[30]},
      {stage1_18[15]}
   );
   gpc1_1 gpc137 (
      {stage0_18[31]},
      {stage1_18[16]}
   );
   gpc1_1 gpc138 (
      {stage0_19[30]},
      {stage1_19[10]}
   );
   gpc1_1 gpc139 (
      {stage0_19[31]},
      {stage1_19[11]}
   );
   gpc1_1 gpc140 (
      {stage0_23[29]},
      {stage1_23[11]}
   );
   gpc1_1 gpc141 (
      {stage0_23[30]},
      {stage1_23[12]}
   );
   gpc1_1 gpc142 (
      {stage0_23[31]},
      {stage1_23[13]}
   );
   gpc1_1 gpc143 (
      {stage0_24[22]},
      {stage1_24[13]}
   );
   gpc1_1 gpc144 (
      {stage0_24[23]},
      {stage1_24[14]}
   );
   gpc1_1 gpc145 (
      {stage0_24[24]},
      {stage1_24[15]}
   );
   gpc1_1 gpc146 (
      {stage0_24[25]},
      {stage1_24[16]}
   );
   gpc1_1 gpc147 (
      {stage0_24[26]},
      {stage1_24[17]}
   );
   gpc1_1 gpc148 (
      {stage0_24[27]},
      {stage1_24[18]}
   );
   gpc1_1 gpc149 (
      {stage0_24[28]},
      {stage1_24[19]}
   );
   gpc1_1 gpc150 (
      {stage0_24[29]},
      {stage1_24[20]}
   );
   gpc1_1 gpc151 (
      {stage0_24[30]},
      {stage1_24[21]}
   );
   gpc1_1 gpc152 (
      {stage0_24[31]},
      {stage1_24[22]}
   );
   gpc1_1 gpc153 (
      {stage0_25[30]},
      {stage1_25[13]}
   );
   gpc1_1 gpc154 (
      {stage0_25[31]},
      {stage1_25[14]}
   );
   gpc1_1 gpc155 (
      {stage0_26[31]},
      {stage1_26[11]}
   );
   gpc1_1 gpc156 (
      {stage0_27[26]},
      {stage1_27[10]}
   );
   gpc1_1 gpc157 (
      {stage0_27[27]},
      {stage1_27[11]}
   );
   gpc1_1 gpc158 (
      {stage0_27[28]},
      {stage1_27[12]}
   );
   gpc1_1 gpc159 (
      {stage0_27[29]},
      {stage1_27[13]}
   );
   gpc1_1 gpc160 (
      {stage0_27[30]},
      {stage1_27[14]}
   );
   gpc1_1 gpc161 (
      {stage0_27[31]},
      {stage1_27[15]}
   );
   gpc1_1 gpc162 (
      {stage0_28[27]},
      {stage1_28[12]}
   );
   gpc1_1 gpc163 (
      {stage0_28[28]},
      {stage1_28[13]}
   );
   gpc1_1 gpc164 (
      {stage0_28[29]},
      {stage1_28[14]}
   );
   gpc1_1 gpc165 (
      {stage0_28[30]},
      {stage1_28[15]}
   );
   gpc1_1 gpc166 (
      {stage0_28[31]},
      {stage1_28[16]}
   );
   gpc1_1 gpc167 (
      {stage0_30[19]},
      {stage1_30[10]}
   );
   gpc1_1 gpc168 (
      {stage0_30[20]},
      {stage1_30[11]}
   );
   gpc1_1 gpc169 (
      {stage0_30[21]},
      {stage1_30[12]}
   );
   gpc1_1 gpc170 (
      {stage0_30[22]},
      {stage1_30[13]}
   );
   gpc1_1 gpc171 (
      {stage0_30[23]},
      {stage1_30[14]}
   );
   gpc1_1 gpc172 (
      {stage0_30[24]},
      {stage1_30[15]}
   );
   gpc1_1 gpc173 (
      {stage0_30[25]},
      {stage1_30[16]}
   );
   gpc1_1 gpc174 (
      {stage0_30[26]},
      {stage1_30[17]}
   );
   gpc1_1 gpc175 (
      {stage0_30[27]},
      {stage1_30[18]}
   );
   gpc1_1 gpc176 (
      {stage0_30[28]},
      {stage1_30[19]}
   );
   gpc1_1 gpc177 (
      {stage0_30[29]},
      {stage1_30[20]}
   );
   gpc1_1 gpc178 (
      {stage0_30[30]},
      {stage1_30[21]}
   );
   gpc1_1 gpc179 (
      {stage0_30[31]},
      {stage1_30[22]}
   );
   gpc1_1 gpc180 (
      {stage0_31[30]},
      {stage1_31[8]}
   );
   gpc1_1 gpc181 (
      {stage0_31[31]},
      {stage1_31[9]}
   );
   gpc606_5 gpc182 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc183 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], 1'b0},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc184 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc185 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1163_5 gpc186 (
      {stage1_4[0], stage1_4[1], stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc187 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc188 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc189 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[3],stage2_7[3],stage2_6[3],stage2_5[5]}
   );
   gpc7_3 gpc190 (
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[4],stage2_7[4]}
   );
   gpc7_3 gpc191 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20]},
      {stage2_9[2],stage2_8[5],stage2_7[5]}
   );
   gpc606_5 gpc192 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[3],stage2_8[6]}
   );
   gpc606_5 gpc193 (
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[4],stage2_8[7]}
   );
   gpc606_5 gpc194 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[2],stage2_9[5]}
   );
   gpc606_5 gpc195 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[3],stage2_9[6]}
   );
   gpc615_5 gpc196 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], 1'b0},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[4]}
   );
   gpc2135_5 gpc197 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage1_14[0]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc198 (
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc199 (
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[5]}
   );
   gpc615_5 gpc200 (
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[3],stage2_15[4]}
   );
   gpc615_5 gpc201 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[4],stage2_15[5]}
   );
   gpc615_5 gpc202 (
      {stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[12]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[3],stage2_16[5]}
   );
   gpc615_5 gpc203 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage1_17[13]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[3],stage2_18[3],stage2_17[4],stage2_16[6]}
   );
   gpc615_5 gpc204 (
      {stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_18[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[4],stage2_18[4],stage2_17[5]}
   );
   gpc615_5 gpc205 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], 1'b0},
      {stage1_19[6]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[5],stage2_18[5]}
   );
   gpc606_5 gpc206 (
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[2]}
   );
   gpc2135_5 gpc207 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4]},
      {stage1_23[6], stage1_23[7], stage1_23[8]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1]},
      {stage2_26[0],stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2]}
   );
   gpc615_5 gpc208 (
      {stage1_22[5], stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9]},
      {stage1_23[9]},
      {stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage2_26[1],stage2_25[2],stage2_24[2],stage2_23[2],stage2_22[3]}
   );
   gpc615_5 gpc209 (
      {stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13], 1'b0},
      {stage1_24[7]},
      {stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[3],stage2_23[3]}
   );
   gpc606_5 gpc210 (
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[4]}
   );
   gpc606_5 gpc211 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[5]}
   );
   gpc606_5 gpc212 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[3],stage2_26[5],stage2_25[6]}
   );
   gpc606_5 gpc213 (
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[1],stage2_28[3],stage2_27[4]}
   );
   gpc606_5 gpc214 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[1],stage2_29[2],stage2_28[4]}
   );
   gpc615_5 gpc215 (
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10]},
      {stage1_29[6]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[2],stage2_30[2],stage2_29[3],stage2_28[5]}
   );
   gpc615_5 gpc216 (
      {stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15]},
      {stage1_29[7]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[3],stage2_30[3],stage2_29[4],stage2_28[6]}
   );
   gpc606_5 gpc217 (
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[3],stage2_31[4],stage2_30[4],stage2_29[5]}
   );
   gpc606_5 gpc218 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], 1'b0},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[4],stage2_31[5],stage2_30[5]}
   );
   gpc615_5 gpc219 (
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], 1'b0},
      {stage1_32[6]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], 1'b0},
      {stage2_35[0],stage2_34[1],stage2_33[2],stage2_32[5],stage2_31[6]}
   );
   gpc1_1 gpc220 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc221 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc222 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc223 (
      {stage1_3[12]},
      {stage2_3[4]}
   );
   gpc1_1 gpc224 (
      {stage1_4[15]},
      {stage2_4[7]}
   );
   gpc1_1 gpc225 (
      {stage1_4[16]},
      {stage2_4[8]}
   );
   gpc1_1 gpc226 (
      {stage1_4[17]},
      {stage2_4[9]}
   );
   gpc1_1 gpc227 (
      {stage1_4[18]},
      {stage2_4[10]}
   );
   gpc1_1 gpc228 (
      {stage1_9[12]},
      {stage2_9[7]}
   );
   gpc1_1 gpc229 (
      {stage1_9[13]},
      {stage2_9[8]}
   );
   gpc1_1 gpc230 (
      {stage1_9[14]},
      {stage2_9[9]}
   );
   gpc1_1 gpc231 (
      {stage1_9[15]},
      {stage2_9[10]}
   );
   gpc1_1 gpc232 (
      {stage1_9[16]},
      {stage2_9[11]}
   );
   gpc1_1 gpc233 (
      {stage1_9[17]},
      {stage2_9[12]}
   );
   gpc1_1 gpc234 (
      {stage1_12[12]},
      {stage2_12[7]}
   );
   gpc1_1 gpc235 (
      {stage1_14[7]},
      {stage2_14[4]}
   );
   gpc1_1 gpc236 (
      {stage1_14[8]},
      {stage2_14[5]}
   );
   gpc1_1 gpc237 (
      {stage1_14[9]},
      {stage2_14[6]}
   );
   gpc1_1 gpc238 (
      {stage1_14[10]},
      {stage2_14[7]}
   );
   gpc1_1 gpc239 (
      {stage1_14[11]},
      {stage2_14[8]}
   );
   gpc1_1 gpc240 (
      {stage1_14[12]},
      {stage2_14[9]}
   );
   gpc1_1 gpc241 (
      {stage1_16[12]},
      {stage2_16[7]}
   );
   gpc1_1 gpc242 (
      {stage1_19[7]},
      {stage2_19[6]}
   );
   gpc1_1 gpc243 (
      {stage1_19[8]},
      {stage2_19[7]}
   );
   gpc1_1 gpc244 (
      {stage1_19[9]},
      {stage2_19[8]}
   );
   gpc1_1 gpc245 (
      {stage1_19[10]},
      {stage2_19[9]}
   );
   gpc1_1 gpc246 (
      {stage1_19[11]},
      {stage2_19[10]}
   );
   gpc1_1 gpc247 (
      {stage1_20[6]},
      {stage2_20[4]}
   );
   gpc1_1 gpc248 (
      {stage1_20[7]},
      {stage2_20[5]}
   );
   gpc1_1 gpc249 (
      {stage1_20[8]},
      {stage2_20[6]}
   );
   gpc1_1 gpc250 (
      {stage1_20[9]},
      {stage2_20[7]}
   );
   gpc1_1 gpc251 (
      {stage1_20[10]},
      {stage2_20[8]}
   );
   gpc1_1 gpc252 (
      {stage1_20[11]},
      {stage2_20[9]}
   );
   gpc1_1 gpc253 (
      {stage1_20[12]},
      {stage2_20[10]}
   );
   gpc1_1 gpc254 (
      {stage1_21[6]},
      {stage2_21[3]}
   );
   gpc1_1 gpc255 (
      {stage1_21[7]},
      {stage2_21[4]}
   );
   gpc1_1 gpc256 (
      {stage1_21[8]},
      {stage2_21[5]}
   );
   gpc1_1 gpc257 (
      {stage1_21[9]},
      {stage2_21[6]}
   );
   gpc1_1 gpc258 (
      {stage1_21[10]},
      {stage2_21[7]}
   );
   gpc1_1 gpc259 (
      {stage1_21[11]},
      {stage2_21[8]}
   );
   gpc1_1 gpc260 (
      {stage1_21[12]},
      {stage2_21[9]}
   );
   gpc1_1 gpc261 (
      {stage1_21[13]},
      {stage2_21[10]}
   );
   gpc1_1 gpc262 (
      {stage1_21[14]},
      {stage2_21[11]}
   );
   gpc1_1 gpc263 (
      {stage1_22[10]},
      {stage2_22[4]}
   );
   gpc1_1 gpc264 (
      {stage1_22[11]},
      {stage2_22[5]}
   );
   gpc1_1 gpc265 (
      {stage1_24[20]},
      {stage2_24[6]}
   );
   gpc1_1 gpc266 (
      {stage1_24[21]},
      {stage2_24[7]}
   );
   gpc1_1 gpc267 (
      {stage1_24[22]},
      {stage2_24[8]}
   );
   gpc1_1 gpc268 (
      {stage1_25[14]},
      {stage2_25[7]}
   );
   gpc1_1 gpc269 (
      {stage1_27[12]},
      {stage2_27[5]}
   );
   gpc1_1 gpc270 (
      {stage1_27[13]},
      {stage2_27[6]}
   );
   gpc1_1 gpc271 (
      {stage1_27[14]},
      {stage2_27[7]}
   );
   gpc1_1 gpc272 (
      {stage1_27[15]},
      {stage2_27[8]}
   );
   gpc1_1 gpc273 (
      {stage1_28[16]},
      {stage2_28[7]}
   );
   gpc1_1 gpc274 (
      {stage1_32[7]},
      {stage2_32[6]}
   );
   gpc207_4 gpc275 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc276 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], 1'b0},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc277 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc23_3 gpc278 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[1],stage3_8[1]}
   );
   gpc2135_5 gpc279 (
      {stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[2]}
   );
   gpc1415_5 gpc280 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage2_10[3]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[2]},
      {stage3_13[1],stage3_12[1],stage3_11[1],stage3_10[2],stage3_9[3]}
   );
   gpc1163_5 gpc281 (
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_15[0]},
      {stage2_16[0]},
      {stage3_17[0],stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2]}
   );
   gpc615_5 gpc282 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], 1'b0},
      {stage2_15[1]},
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage3_18[0],stage3_17[1],stage3_16[1],stage3_15[1],stage3_14[1]}
   );
   gpc1163_5 gpc283 (
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage2_19[0]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[1],stage3_17[2]}
   );
   gpc615_5 gpc284 (
      {stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[1]}
   );
   gpc615_5 gpc285 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10]},
      {stage2_20[2]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[1],stage3_21[2],stage3_20[2],stage3_19[2]}
   );
   gpc606_5 gpc286 (
      {stage2_20[3], stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[2],stage3_21[3],stage3_20[3]}
   );
   gpc615_5 gpc287 (
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], 1'b0},
      {stage2_24[0]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1],stage3_23[3]}
   );
   gpc615_5 gpc288 (
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage2_25[6]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[2]}
   );
   gpc7_3 gpc289 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage3_29[0],stage3_28[1],stage3_27[2]}
   );
   gpc615_5 gpc290 (
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4]},
      {stage2_29[0]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[0],stage3_29[1],stage3_28[2]}
   );
   gpc117_4 gpc291 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5], stage2_31[6]},
      {stage2_32[0]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[1]}
   );
   gpc2135_5 gpc292 (
      {stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage2_33[1], stage2_33[2], 1'b0},
      {stage2_34[0]},
      {stage2_35[0], 1'b0},
      {stage3_36[0],stage3_35[0],stage3_34[1],stage3_33[1],stage3_32[2]}
   );
   gpc1_1 gpc293 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc294 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc295 (
      {stage2_3[3]},
      {stage3_3[2]}
   );
   gpc1_1 gpc296 (
      {stage2_3[4]},
      {stage3_3[3]}
   );
   gpc1_1 gpc297 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc298 (
      {stage2_4[7]},
      {stage3_4[3]}
   );
   gpc1_1 gpc299 (
      {stage2_4[8]},
      {stage3_4[4]}
   );
   gpc1_1 gpc300 (
      {stage2_4[9]},
      {stage3_4[5]}
   );
   gpc1_1 gpc301 (
      {stage2_4[10]},
      {stage3_4[6]}
   );
   gpc1_1 gpc302 (
      {stage2_6[0]},
      {stage3_6[2]}
   );
   gpc1_1 gpc303 (
      {stage2_6[1]},
      {stage3_6[3]}
   );
   gpc1_1 gpc304 (
      {stage2_6[2]},
      {stage3_6[4]}
   );
   gpc1_1 gpc305 (
      {stage2_6[3]},
      {stage3_6[5]}
   );
   gpc1_1 gpc306 (
      {stage2_8[3]},
      {stage3_8[2]}
   );
   gpc1_1 gpc307 (
      {stage2_8[4]},
      {stage3_8[3]}
   );
   gpc1_1 gpc308 (
      {stage2_8[5]},
      {stage3_8[4]}
   );
   gpc1_1 gpc309 (
      {stage2_8[6]},
      {stage3_8[5]}
   );
   gpc1_1 gpc310 (
      {stage2_8[7]},
      {stage3_8[6]}
   );
   gpc1_1 gpc311 (
      {stage2_9[12]},
      {stage3_9[4]}
   );
   gpc1_1 gpc312 (
      {stage2_12[3]},
      {stage3_12[2]}
   );
   gpc1_1 gpc313 (
      {stage2_12[4]},
      {stage3_12[3]}
   );
   gpc1_1 gpc314 (
      {stage2_12[5]},
      {stage3_12[4]}
   );
   gpc1_1 gpc315 (
      {stage2_12[6]},
      {stage3_12[5]}
   );
   gpc1_1 gpc316 (
      {stage2_12[7]},
      {stage3_12[6]}
   );
   gpc1_1 gpc317 (
      {stage2_13[3]},
      {stage3_13[3]}
   );
   gpc1_1 gpc318 (
      {stage2_13[4]},
      {stage3_13[4]}
   );
   gpc1_1 gpc319 (
      {stage2_13[5]},
      {stage3_13[5]}
   );
   gpc1_1 gpc320 (
      {stage2_15[2]},
      {stage3_15[2]}
   );
   gpc1_1 gpc321 (
      {stage2_15[3]},
      {stage3_15[3]}
   );
   gpc1_1 gpc322 (
      {stage2_15[4]},
      {stage3_15[4]}
   );
   gpc1_1 gpc323 (
      {stage2_15[5]},
      {stage3_15[5]}
   );
   gpc1_1 gpc324 (
      {stage2_16[7]},
      {stage3_16[2]}
   );
   gpc1_1 gpc325 (
      {stage2_17[3]},
      {stage3_17[3]}
   );
   gpc1_1 gpc326 (
      {stage2_17[4]},
      {stage3_17[4]}
   );
   gpc1_1 gpc327 (
      {stage2_17[5]},
      {stage3_17[5]}
   );
   gpc1_1 gpc328 (
      {stage2_20[9]},
      {stage3_20[4]}
   );
   gpc1_1 gpc329 (
      {stage2_20[10]},
      {stage3_20[5]}
   );
   gpc1_1 gpc330 (
      {stage2_24[6]},
      {stage3_24[3]}
   );
   gpc1_1 gpc331 (
      {stage2_24[7]},
      {stage3_24[4]}
   );
   gpc1_1 gpc332 (
      {stage2_24[8]},
      {stage3_24[5]}
   );
   gpc1_1 gpc333 (
      {stage2_25[7]},
      {stage3_25[2]}
   );
   gpc1_1 gpc334 (
      {stage2_27[7]},
      {stage3_27[3]}
   );
   gpc1_1 gpc335 (
      {stage2_27[8]},
      {stage3_27[4]}
   );
   gpc1_1 gpc336 (
      {stage2_28[5]},
      {stage3_28[3]}
   );
   gpc1_1 gpc337 (
      {stage2_28[6]},
      {stage3_28[4]}
   );
   gpc1_1 gpc338 (
      {stage2_28[7]},
      {stage3_28[5]}
   );
   gpc1_1 gpc339 (
      {stage2_29[1]},
      {stage3_29[2]}
   );
   gpc1_1 gpc340 (
      {stage2_29[2]},
      {stage3_29[3]}
   );
   gpc1_1 gpc341 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc342 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc343 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc344 (
      {stage2_32[6]},
      {stage3_32[3]}
   );
   gpc1_1 gpc345 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1163_5 gpc346 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc347 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1]}
   );
   gpc135_4 gpc348 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0], stage3_10[1], stage3_10[2]},
      {stage3_11[0]},
      {stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc207_4 gpc349 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc606_5 gpc350 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[1]}
   );
   gpc1163_5 gpc351 (
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[1]}
   );
   gpc1163_5 gpc352 (
      {stage3_19[1], stage3_19[2], 1'b0},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage3_21[0]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc1423_5 gpc353 (
      {stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[1], stage3_22[2]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3]},
      {stage3_24[0]},
      {stage4_25[0],stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1]}
   );
   gpc135_4 gpc354 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage4_27[0],stage4_26[0],stage4_25[1],stage4_24[1]}
   );
   gpc615_5 gpc355 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4]},
      {stage3_28[0]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc2116_5 gpc356 (
      {stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5], 1'b0},
      {stage3_29[6]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[1],stage4_28[1]}
   );
   gpc1325_5 gpc357 (
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], 1'b0},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[1]}
   );
   gpc1_1 gpc358 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc359 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc360 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc361 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc362 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc363 (
      {stage3_3[3]},
      {stage4_3[1]}
   );
   gpc1_1 gpc364 (
      {stage3_4[6]},
      {stage4_4[1]}
   );
   gpc1_1 gpc365 (
      {stage3_5[1]},
      {stage4_5[1]}
   );
   gpc1_1 gpc366 (
      {stage3_8[6]},
      {stage4_8[1]}
   );
   gpc1_1 gpc367 (
      {stage3_11[1]},
      {stage4_11[1]}
   );
   gpc1_1 gpc368 (
      {stage3_18[1]},
      {stage4_18[1]}
   );
   gpc1_1 gpc369 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
   gpc1_1 gpc370 (
      {stage3_36[0]},
      {stage4_36[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor_CLA32_32 compressor_CLA32_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdb1cf9d234d5d7201f8d862dc04dfe031c9e76b8f02bcc931a849bdd67d3f592fc5e81080b73de6846d8dc4c6200ac4cbbd424b4154b962db2a108e6bd4db79e7a11e0e8b86dfb58d44b31448c38580f69431ee67c4c8f7a6907310c535cf033b3ef5e26c2b04075909a014c384b6a901e6dddca5228a2fe36e605b87739adb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7ce7819968f461184c262c5dc2697bf3917c839f6b3664a1785285fa33a581a452d5c9eddf7643ecf4cd63499d7370449f6f3ddfb678b5e00e7d2e7798ba01ca918fbf135c57d61c5e7cb38f37f7a1b492a7284dc260e57ccaa3976e01f37dc4458ff02c6dccb17acad381b97923b3cf88527e688b6b96cf355cd7b68b67318;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80138dfff8b47ce04dfd08a691f42bc525837266bf5c7c7df42b80032c7dd642684e42f57de46f1eb5bc1396111a207fd0b34c765677c1e34bf55043f79ddd9f472f6ab410727ab697922312707b8b44ea8d7654320b67829211a0d33355925a5aae00455987ca962b01edb5db8b93cd192ac635a10b1cf637164b85a558cf41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98437f6315b358d246d8230d929cc4adb37e8c1f772c91468a6e0b817f015733977efef3383f676add0ff56d61ddc49bab61c27d425ea16ad0982284d4b159f55aa4e3f3d0a65d8c855c7cab8088d9aaf4384674b94fd9f58b239c8f96a8edbb68febb0d16390dbc5453a6608c2691a126ca8a73460394d2654823360d702d03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97e2fc23ab8e3f692d3ca588cbdf7458859567367284973f4fb54ce922a4b85bb5cdfd7dbe4cbcba87aab4ae3e673e13c7ca9519c44f9fb44a098ee82480aefdac506919fb86a5fbfd1556fbd7021be7058d49041be447fe2fa3b9b2457ed1d08e14f56ab8b00283d1132fae31ac412634e8acbaf183716f431adf46c7ed9994;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1d961f077593e9bf5e650582590b69d8099719d206edc8d074c04c25702859eaee88d1f2be38a457506bc5268a9a04859263a3c773d4ccaa501245b1259f4fc7e28fb1fb52999e602fe0f6e0b9526807274f407c4f6dc89628853ca5ff5bcf6c04591bdad6525ab68a607babc854093e87062fbea3261d34c885454f7b42a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb7f3c3b52174dcc9c4bf32b9e8ba72ad06274ac4387b07ee9869e86bf04ba6d7efbad7fb345d075fc7cf8e16b56a29cff40c1605102464c1d8e5d07878810657b1697fb50b5e3a7957a51208228a4259c2a34e3ae100fec019859d413aad0950f72fd52b5c61c66653d5f2a68ec9628d8a388e2b683e8ac305d7ab604ba4bc3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee0b8711c68ed5f5b4e86952c8ef1f4b9ceb533a1cd1dadecf2e0a7867c0fbf9ed171b8432de9f1f80c2f79347f8a23e7b883c81be023d1c0844912ad128dfea01de9900f6530b86a19cc5988f61096a6d520924ea7811ed79f9b22045d39135a39bf8917ed65d12bedb9a0b66e47801dd79291c0376fe6117b85ae9986004cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heccf3264fb1fa2f384ea874005749d3885e406af47069c25179f3419b2cdcb52864a092f234ed2146d43a19b858597865fd55dead4ad61208e51c0c176ee0f733820e6ec1e768ac5f6bdf66a2e745eb5b3686aa1c7c6a78b537aab7afe3deb64bf8faa108babfe3ba082237274995888aadf3610e4f913978ea781d9a2d24226;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h303a79a5344d784ad4637e1cc0eaf4845e30bb39f8da5ec737a0e3990ad87249d383cc13df1253a35a88a279acfffd24ee4cc544c2859af1d80d3aed70704bf107865d6550ace0e94132e4e941482470b301a99b7b9a5d0751ad39e53ecae040a05340b7ba3ed097c00fc17aab2f603f82c2958f6c462f2f7662dcb1d13f8d65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h235beede310ba33b5b246a16a6704ec8910babec2423fe440666dbcbaf103614a3c34036ccc2fd06c9229e5f12c389466a38557d07109965d818751cb7436f36339c4b349ce1e4f973dca0613aa8fa3ec1eab33069abba76206bccec4afd782fd5d850fb64742fad64808e529e2f098c16e6791301673e7a662c0804d9fbd72d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e06cc12552d6e32a4072a9949c75169e3fbe8e08b0fd4978b42b891a248036838fa517d1070f2a8a88a477d3f68d4fb0ceadeadce8b3cf6d476aa5286ad295206f472c7e9d775f231b88fb815bb24e037110b5ffc0699646071cb907a863f42c5c70b6fbc2d311fc51b0ca58459f8e894860c80f6bd8b161fcad4df8803ad4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6fed0137e0a7b7b3f9afe204d4556c55ca0e9bfae7156d55028f6fd4db37f40de0e65086e60af1ac515246b2377a00127b5d7fd5a29ab8c32e8461b5f8035033137ea4a6e60ff82c4b3e12d36cd4da8b357554ab9cdb3f05bf4fa71675ebf972aea5b4f8ed9fc3181e8c89389b4cbfb8b403879bdc55170b75519347c586e8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6149e18042ff32cce5e7460ab2f924e71d21e8f64e8dd7d65a4d86e1c64e0d55c4e2a386811af65da01c898ddad1acfe1cfa64b3b966f93983fe56020eab20ce1450477f6067c9de458f8dd0e3e836ad95d556490b65911aa655731c71e10325ed9ca00fd0b5d30b724402b0f47fa8324a945a0c0481d5ea1568cdcca78ca7fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf876095e5d3138bf21ee61e6f87d51c67aa3b119989674f20352c5dc0e08828115c03beea6c1d7bf47df51c1dfc0dae4196bb37d2920d3ac84efb36e810b3b8a21b78ce2b66c15c669a4b08e44fb1c30529bdbf053806b645c01913637b080da8207352e488846f79dcd1461bd204aab47178a28f23774e9c8195aa9298fd26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ef591f9f27593bb71877fd6f7ba824779987ea98b30e6bd590da01d17140bcf0d0eeed93c4ecf8b301f99a2fb2b55977855603df9cccbe5edd8987a0c6eb015b41f25eb29208858e6c149e319ba3dd4fb34b47cc0f900018898cd613618d2e57c6269302f554d353a0506f0fd01acd26a2c858cde754cb87e34a9a1dbc962d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb47d645a1ecb329084cfa02547e1175c325cfa7fa3e8586ea46fb1855bb13791453536104269fd931fbf59e5cd6b87436c6cea285f636d1f9976af92593d1aed631026c3c4a539a50adea6e01249c325c348fe4272a2ca2fa6832a09b2ff2e5f54558d7ab87d258960fc38bb822c50a280cc69555e42dc04271c6464ed32239b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fc6f98c390edd856e28276303d08b7fd10ecf18b141204b4507e6ba3f84e0eedf6677a2225518b0ed9d513229e478db40a975a4463c5b46b368022a91f641a0fb6806b6de1c7cb233ecff6eaf8e20e2e7f0594255ead11e32b6c1163e7bf346aee91c39a39164abc6d80e2b67f5a42e885903f265cdb2e6d5c1ea5c2678c3c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3544ec2c345616839508170d75f4c6794588deb27ec7d607516dafdb10d3b55cf1f44190e6f7f63b9ce2692b2aa0c1e159b979677d2b26f5a582cd3c5fc3bdf19b7bde407aae78f5a175d05cd345cec528e4864ce939888da23f8c2f55b7c5f44dd95c31c6ee4f5694d2475a58a5aeed8d113032c80c4d8350de742b28007cd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha14d5cff612bddca7e78809d3498d6b2fa30e7f1dffcfdba540b6b1d6d5cc1ccd641aa9ca703b5fcfef46e1cf5aa8984b8a996930889bb8a95423948801b7f90622f0891c3ebafb1c1dac3c1471d6a24feeeb364d1edef2e0a60b73807554e1eefea8abbb759a41c51e335b7e9c86a635c856e17cf008dd413a0cf4e0ed17251;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ecd034cc73d57d950556c6f3e64791887305f0d41040059548ab21aa638da8b1aef0d5960e9037bcba3701cebab7efa14a7905a7a1f94431434bf1a27474655b52c60b987aacd16f4edca3a596fa60586bb6b333e8d7eee659654748bb95c442e513f21aa068566bd37abb7c2d4a2daa19343a8da7de669baae556e4e354ae3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30358d9083011a1ae8327e17b9a24d520174f44c4c496ac644781260f61158132a3d70a50bde8223048a6522e9dbd87f77597677ada6202c71f0228759c9cceab6d8ffde060aae403fd03ec89d479fba7133be43e052b7a6818830fdb0405ec9b365600346417e76c5a7e2c941e19e43f75624172ca799b77d53200287a24359;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc9f8e9f32cc5397e6aede0b14de0bf21469f45198361be4414ca52584dcb145212d7a07949d864bfe4e7ad6f94b05db13257f435d30dfc20c52bde86993b474b2c0f19146b558f08d0cc55f9e86cf4d5bb22f4224740ba169638d51fd7c9f4abb56ebdff837288a38534aad1e7eb72ebd83b638d5dde37dc8c1e014815c39ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h463e9fe4dd427643b32ea6088d2a09cf58383f8257887d9bd0dabd050b65bc6898ef65199d00e7361ade7958b41f0d36f3e5c72a0ef505056a35ae2042a079e377f2008a83157f947a9ff1c827cf9ed72747003e369efe864d44f73655218909a48e842b8188b75fce702b38fd2d5f270c99729aa4721ac5864cf2452546fa96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb2a0a82a71cb0ea25588a5adcc4a922d85057f10f8e0d7d20a4fc104bcbc36e3babae9701599079ebb7a97ee2312b2e80856b46e6ee16cee1a04fdfd476bed1dbf28f307ca297ab6e2e43596191551492a356ac37377848a61c01b154be61614ff6b621ff5721423397b3d8a90d7e48ea2aeb488284e3577df126a25824fa80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habddecd56189461d856a52ae512c323f6df2c3eb7644555c3e4a00f5d6dcc2ee5bf3fd4d411558205cba0ffd1ff1b3143a9f83319d61c42a6aa54187d9159edeb068ec9be4e87553bb686ac8556972961309991e94b6aa8cca9a574b6b4920de390e96e55ada510b1e0fe6d71a3dcdffe7c65053b7290e68957ba83ea5aa8db4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf60df9d7787e264130206b0ab597391ac78445ebf21bf6060c9fe2fd5ffe02e3d6456545e9a392bb64e17a6666358e13712e75bd210ae8c7b4cf1929f4667efdaa57a2feb81bdbc95c3e127634b3c637efa28c3a21cadff8b8de6729cd872c5445d7d780d794bef93f034ba7f21f70876c9af2a991b23210432e75675ff0de5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5cb781fe54b99bd10ad1402bbda408833b46f7da8a5bdcb20cf635d6a06bddc029b7b4a62ca69847c1c5d3231987ff6df14a6a9833d8a00fef611a6699108302b65eb727e37e69a7340fd5103bd263fced2c2b71940f129b7c7e61192af4b18b7b7fa030c4a10533df74a00a39a5c5cc9b7eca66a73016cf1332de18e1a524c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6ebb8e998e689954a88fdf117439d86dde2fbc799e632fbe2f9068dd49ecb9f1c3283b957ab2d8a23dbf7041554d4b26a0217a83716c86c186fd89fa82549be1800be536e5b1643ae03922bf5e61a863e69277c0e7a3b2a0ecd3b9f084943a948d208e7fe7074b4beb9a5a660d63f87348c6a65948a51fe07b213d76e0ad379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c655465372a9282f9e0575782b482e96f2830a44aeaf31e70a115a1a45445a945955fbbedb3507313f887d688aed525071484b7321bfbb2ff44971c8159b044bd610c6810f8652671caf9321c403e5708bd3861c67db025ca120ff3f72572bba19c12f3aef7968c2fb2782c338adbc73cc6bd1e13c262e859694f0ce380e112;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b0572a30f166ee235de86005e624d267a646aaf6ccd4f34faf16ecd7d6e844d073169443fe776e320f35b38ad62ec831cd4bbb5016a3127097e11a6ebab389971275120f055f30d05b588ebd4af0c00b04d90e925abc933b65a9c8710cc2c83fc3650d62fe4d007e00eef612392638fca75990972d495c5bedcca04beb1f18e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8582b85f69b57392d236c9d7b5bcbc8b515adf8aa1cacb0fb428a350cded398da238e3f103771402847946f0918286c41632898bbc3a3461ef9af5b5f2839dace8416042218cef47ebd906f615d18de6d98dfa648962489e5f6f5ac074f482fbe1d30b9bb46a6b1ab88a64d6850ef7438a36b9016e167a0eed2827e0a07c0e0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc389d5ceecbce261beaf3b53987b093e574948229bbb454f1c254c1d49b3ad99ae0bf05e104b09c1486dff8dcf31b58c82c380d2140070c5f648943db0b39a6f4ef0de89198942bf7d0fdc913fdf2eb6e6fb9a25339d9fb7d2d3f0f86b2ae5fb3ccbaf5ae32ba8326de8d15dbf7ea0833164103b94480e0f9e20bca8f212c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1f746a8b4e7615b5f1aaae4bfd19adcbdced7d992c82bdff27e0f5c75709a9a3e0e4c3a66ec693b1b7c5af72878811862b77bf4a918b62fd0df003b058d7e43f0c26d7256e94b1295b35c08377baa932e9c826c79d128beb16a6654dd19f2a24ca7aa791f6d41435c66f1c69377ce51e21ffc245f98db654b8823437d224819;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h870ab333658cdeb6d91cf6bf5dc7630bf4e58cc73a25e286930ef59f703c2fd82aad286f2d3e6ce4e1f558674368df7797837c4cfba408f986c13c92550a00c282e257c3415c018ffd273ad8e0bc5d6a8bdd1d6f62d8970fe24488f08d5dfd2361ccc1a205fb5a04df52980cae722e9f5e68302ac2e259060962898d1dd04652;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha904a5982b86159cb765b66b54fb00d03cb53ffceefa850e40598cc7c9d80fe740418e48bd4f52e57d0567b88b3acd1653a80e200c9fc2070ce5b1a4835b83da156c1be76cb2544fe46dca5658e46a11aa923d84e78d7e39546f5ae9adf43c46ca21b46708b4fb24646b348e1fb1d6d640d91d818aa42d974c3a64373872e6c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h844c1a7c93b849168690d0d26c2a76bada6b3dffe5c955bc6b0a64eab0ee9c678c7a93c1b6e0a4cf60bab5113134356fb05c6a736e036cc1b7cfe539c0ba25935e1b593d5c50a8c2ce4158d07a098fe9eb1ce4a3dacbf3ca2ff94add48aa5aa1c1d82e919a34fcb2825588f04a9471e94d821020dc9513ea6fdd0468fe73dab6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb80c6d202b8f099a550e3299c1456e89c248f649816065bdd37d3c38c391544ddffae649fbd0b06f439f39602bdac2b45b358e153eb9e7820a328967266dc5da6e54fb572731c7a2503555d3e44eaa9e3a75dc46ccc582d041b18548a54fa0ac111666e0b6f409653fe085927ad2a1131f626d0f4dafd5ec37c65016173f6e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb64ec0e88fd1ade6e2fcc0194d8b25bf2977c7bb1a2dba639c7b2f59d3493bfef491d1f6b34432eb41b5f50fc8f381c251c4bc19662ad1cbfc0ae51cd585a4cdcee4fa5335da761e75c065e46f8c4a5a2fbc6657e6d03eba4f127b9148a58499baa7535453eb1c3d712621ac302364fe21208d93554c47f29bf6083f5db9a9e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0e3871b9abc9b6bd353304fd771f979f7b493c32626dc199b49357e148850eed5f59cd2330eaba1f2b4b1b1384afd9429ec06ccf15991af3f4eabf7739cc938794e1aa02d277cf3724ceb282b0cb00f8947343cb345c27744af158f5b08d2c095186b8866eff23c52b1382514a73c6204d8bf935fe68961ab859bdc8a4a2433;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd69e0cd769ad92b8370b861723562feee472232cb8827faea4ea2728337a85d570ded2f5d689559243e7e835e6f8e450a70981620129c3db53e773b1ddf3a345bab60f0a5ecd148519e49d5a545a912d636defc931af892fa6afdcebcd2097a3d1b12dcb710608931b1750e2a6148a242e470008780e327591b7947259a31e24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fe69ab02729e7a4b27adf84765520f8a9a6dbe602038b91c07584cb77e54703e43eb6f2cf0c15fc130f876164aaa2651274fda871e1e103812c663f6e2952a4765b673d24ce4446a0436d2c96c911d3c464c75f0e808db492343f4b9b041e7e432a10968a3e000a244ade289867d7784dfede8785aeaa7a16c8a7401371b4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81a5e8e6070d5d1eeb838af783064654cbe81f0e092c399e0c242e7b6ca0113eee21ac0c67fff34e17b1b402ca4a4db961633309c4a5cf9205969325126c09f095a7a326eb06c82266f21517d76f76daaf1af3e36fad5a3383c396fa482854b04bdab65ff781eab5aba79b6422f4b6d3f79091ea6824fa02fa2e3711e00b1164;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf0b7e802e495a9861bb6b17d6379ec257e5ba083826e2110c5cc836c2e9801b85ece24b64549fb5f325b9ac38bc2d08824d1f403427c178461bacc9b359808ee0815e5630e99b7d0cf2c21cb679c0c3b27b7c23dbd7b953b81b8ab32c0c9e518987229511d532b0a36577551d160f931e63452a13dbe21a83518324712ae741;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h120f672f6aafd93eca5574afa22243e80fdd0f630094524055cb36492edc4934b6d498957e6da3aba4a4eaa87650d409f665678b4454ad5a5032b881eab5d7af60aa906a3760638064005aa6f51bc5fd75aa67fbb353778c138f9479c7c3194b4b412eadfdd7a9b06316f465350a97439f3616f43103160f1ea0e85d359e128d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ba153b562fc301418b80a3542b31e9c109d24e0c23b63e7bc610ae5e849e18986d8ebffb3c85fe6a97063ad3273fc127d1b3d3bfa6dadcd6d81fecc87a16e89e848b38156f70007c6d48618c3917244d225f68133ca432cf77875019d440e483e635e115f3f648f3e3a80b34d57db24cffa85cb0958c78768cdfd985814f33a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h472149214231d3eb0a3027de6367f9ad608eacf010e4e70a9a7bdcadfbc44dff1fb02ab6be7fcb0d4b53012008d01d0569e22bc31b1445e59d8dfec8ee9585451d3546c378bd087da47c3b728deceac306e0f181fea152c07fedfefa682a6104309baefe612420c1b3f8cd211adfce8e67aec2be9657d8cda353ea3f8fca5c7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd761c364032fe3446de814c684280c465e1730df930c5a2b75613de52a9c4efa59cb325d34263a9026c922451b1338ca04555f32dc33ba9dd3c7675318583d72d4d4017daa856c6cbe8a1cb620c29b472d55a6d3f209a9d1b71f0eb3b6ecac802e41e95ba2a9ac96f16ae6f417f0f22f896834499c71a5da288816e3f49fd994;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadab6212bc908e14ad62b5ff5fab9c07ad50521dd36fee2262fde0b99d1a101b97a58e0b36bbcebfab49dd523a94621aaebfba26d2c01c6fee8b4edbd24e48bcd90ac3e15f91f77bc040edf737e0ad59e16d3340078e7fa00769de142d881827eb15cdce55053fb5eae8f3381772eda8f439c3b14d84401077dc7bc61be39530;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59bee8c20ff68f868ae10e69ba0bc65ee5de79052584563703b2e0236b565c6a2bf87257a9c8a05d9d05b1e40f65ce983deb899d2664dcfa1543d250ef4d6b9c9fd0d4c6dbe795f2fae782e57d48077d28799727590fef037d337cb8ba4d0abb26969b7ee990a407062f42204e5c7f1f9d144c41cc0bf28f96a20c69fc1a91e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd376525da00ab77e84dbdd43bf597c90b2e09ee9a5bef33d4f90e8cf8542fdac79b5d6b766375367ee435621eb411e0a18702472a0354ebfc575d7f582786255fe4a8ecd5cf08af69650b2360329231703b6efa2d7e2c22b832e699bdd9f4da5c016e2de5fa0ee6253bce5f17e04ea366e64bba22a7c760ec9e09259b858500f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h512f64bda42d9bed0e24744a5e4e588e764919459489ae33d3958b265e6ccdc05fd981f4ee0774f049e1e9630805ac8d72b3ec13504defbf2701fde5ec5624080fe11dc5319200506e6ba3c50d91e985a1aa1aac9a139bdcf188a926eed1ac7e5d0078b3770985650ed35bfc9771ae894fc92f390943514d526ca5df03dc77c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6c8449bb984c1f16223b329cadc3b25608ed2c98b20f9eb410e6346d14acd3028b1ce97bc4e73f455f850b7ec28210fde98be9041401e6e91b4e77505959cd917a7d268fe954afe95f3fc597c9e2f977154c76ce3a518509cf3ee23be17819365e506aedb525a886335dad5de54c0da76335ca188baf6145e89386359e8ce93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he60d4490ba281623935943e86363a6440ed45481af52f8f4870c8a486da154dcd2e602070169229e0260db60a6d59fe9e65f71cf090f0d34a45b519bc51a779e9cb792a7b18755bfa91440c4d936ccef4fa59236d2fef8e104aa604e895550436e9833bee2f3b93fc44090cd89c311cb4e0266d4e3459c76262af90529c83443;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h512f8d20f3d0204887ab4b9cf895095db16d26e84dc3b0d15b015fa178a6aeb6c84cbebbdd7a55ff28549d1120b3a08a8e2813304361a2653f2b6a7fb32955d6b4e730431ee04c9338aca2dfdbd3436c6e6d824f4cb76ac071d3889e8324bd146a3008c10efcd20fa1dfc9747735c7523121958b15f2544be2c930ede42baa87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5626e1e548b8bf18738d5e9eaec7557eba52fbced54bb6b2aeed510b8c7f5b9021569d4877db81f5508b49847282ba4c6319b9674fd0faae0077305527937e49679821dd335bc7323b0e419275199adade3d825b8f7d823bfdada987f5c0f5987d19a14c880f26a9de5ae8794c10b707657164f7dc102a15ca30833a736acf7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h403c2720652c91e5f69e7980923562860412f9125636440ba0ff046096046a0ad2e670a36cd5a5cde54574a0d58228b15b4d0d1f5b89a28aa3484b2c69520463eba28b06bdf3f451e8282ee39079ba72a0832154adf2fffeb08bb0a014b4ad20e231f504fb6a7ccae1053c6b317d38cc1d7625356554f4a173e10d9dc36bf750;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf92dcc7d63ac4ed9a178602a6a348d1ed41193bff97af250229aebbf1294053ba20ba3be66ab14438e02119a37a01838889169a4b0461193f0da0a2f25aa85a3c723255bc3d5cef39de5a86fcb27808570ef1388f83b012d5373285cf48da98ab9af86abc70f26bc83fbb33a517b95eef524da9b9cd272fe7e1e23896805623;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h990d7a2cb687cf5468b0294b5c632e013fa1c6c71c1ff1ecb0c604a273a183d4db98a59ec48a1818bd2254d61bf176d989fe46223271c5d07695734bc7f9466e897d2be15910ca121115b6457a8cd5e50538e08c634d2c856a0090203eed04f6008d54be83e6006ebb8c884f6c691802ac72736e045bddef38bdd652ec9e9a9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h252fd1c95330f0edab6dcbb0a3af52bbc6a4e9b1f3e4524bea261486b35c188d06a9459c3a6bc4f711a4d44c9263152b3a2c0c754cee841d1a36e037f354cb5c23592d223ba0b7efc699fef56bb1e7ec093be68b2e8c22af8197a8d3c86bbd6f39722c938a2704ac011ff6c9f8700c6abc5999d0e2b93e83c86f2783a72e5366;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2ff83ec5be5a4ad35ca2a0afeb19dc2493a7644d1a4f6c80eef29b85fc8148428fdc47e112b137e0ea1170e3d99c2e3ccb619cfc463851916ef705991293830cf8c54cb4b49e6c184d7fd6c8c7d9a862ef463e262135104971af82a206aff4c9b862a03a2fe8623f267a423a2ab2c2abfb42ee421dcbf12b895cafa2a9dace5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe1e1865fb176458db1e93526770ffa7e143b006a5fcde965b61bf6adc28f85a3f298a27471e7a2449b7b1e97c030f6b97a58f42fabfc3713eff7877216c15aa8898fc8a380993bb60d8db00828174f7cb1abcb2ce3991ad17549a1d32dd10a6ac281b5ac77a84ce5796c9556710917363e7e01de1193d4da2b13b2e3533355d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7959767a7900740b56e312c22cbb3ccc0dbaa929c8df006b5a6bc2a3bf78aa15879c4681a4d9c2339fe01a21389ae7b8fe30a4ad068fd23409137af26c460d300c4f3dac5ac875ce657546f5f8e61fc4ce2a5d84eef894cca67171e61751025956032a3be5b39a88fbbc2251ba779526f988d3432396bb2233495fc814f95198;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e56cae4b5b6774a23793718e7902fb200056dbfd1a99a8ea695ec94314a00d4475830bf2299f2cd34d2143035a2de165179f78945b44eb69c4080a174df4d91de07117ece69e06ef458002775732483abfd25b74f22063e72ac5afb6015e796f22eb591d9a5b5d22cb515c9d722cc4e5fc88daf9eee66ef1c7ee65f6a2faec1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9705f3d4c6aa0096835e033bb95709a4474b318b8f19690007d6066d4447d375f00f1f4996d19cbcfa2b759310b5cfc2159116380b5655d0eb17854467e17dace8b88373815ca620fdb228ece66f37372f78187f107707fe1a9a9b95a5ecb64907cde431ca03777ee55ce34ac3dc08b0048b2cdd5f3f08219a1419447befd29b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7293731952cd5c31fcabf23dc2fcf635599b58e06f60adc54def99878ba0193b29b6ea849d766a0c3418d8be54224e59c3b8043b148d721c42ac51e0705b5e3ad50bd1fb70b7f6506469305c2d0f842dc3592a3f41096d54b3f2c8cdc8d9ea8335bed70f135e4bc390be0f2ffeefe187b05d0a03ad2c683253fda5046e85f2e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c20997a149826d115e7728365ffcab59204e9c778c3259a7546e3021927c9d02aafb9fc3cc1663243642ccbc3d423626145e2179007343b03364328d67f1c5a01ca4c72584ab0b7d279fb6c6086ac4d264b3637e9c068b510895baf3f9a8fd8c763d41fd85204bdb554bda9c4fc662ca69d4d1cd68b97e103ba03b673e45708;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fab827a78579f8c86538249072220c559610011c36c320b263fbeddd0816598eb85663e4819df44c39ccc1ad2996c21db1f88b4845fda788def3766e16a7a22ee303826172adc421ee4019494a5d2359c96b63e9654f9efbb4378bfa125e73bc14348e0bbc0becd6085b93bb6a8b0ba920ab359a2f70562db1116bb18fc1d2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bb1a555c35f884a62ee39e5675cf8e85662d1b8ce72671a75199ba96ae708aab8cda7ce521f90f09522b053c5935a4a62b54edbb9037e6669911e76ff3d2631454544242c8a5668c8dfbbd9d1b7effd5515c269d1ad547c2ce13015cfb3c8c95837bdbe2d43c2dd6acd07bb0da9c581e06e92ec7307238851da4ce1a464b7b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bb4b2cb0d8b7a6c81971770628849a9e472a00bebf0b7ff6710ecce62bef755ac46cccaaf330900abd29350ebffa43f04d7987c5baae5b9a8d73695c0f514c6cd8c56474676360301e6d74a5aec6a52aea7af2708cf429d81ed99c76bd34cb11f9173ed58ce43018a68c694276ac7ba3836c32ec01013b68f881d6894a4aa71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70a9a3a31d7b43c110438becb5f99123ca87743050886a3ecde7592dc1c9e0d5c4ca66bcf550853cd8b8400943448f255ac1942830b6d68753f80d7a9bd1b223811d5c6bd8d43a15a9257058f18f39d283cbe0197bc732c03e21eda7a1c6b84e38f891173867abce6bd8e5623b6d136c7c0e3fa483a275e8e3fe285523b9cced;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e035960db7d20323119d761b252ac626e033ec8d1256b0684dee952bbfbd593f45c7ea39aa651654ffa402fbe22c2a338f8ce7b2c24ae15ebb66d93c9dd8ad00711a27894b0f01a6c34d7b95d64dc887dbf139c87a90763a2a476721351b32be2490f10d19bb9c678eb6dd8e3d2d2512c1778cc60d15139001bd7fdc5c3cc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba82a39c8c09f694a90bfbf21ea3512340292cc2f9e66bf706a3198d1037bd0254a7e9589a98d0264b13b541105f0f120f2b74740ea6e4284df440959bfc52e858acd79aeb7d1026c901a38fb9691dd8c2d935d37b5a9a1f057edbb6a9bb163bd5a58f7cd29678a77ac09fe0ca4b46ff58483cdbb6d9db04a7bb6a11cff84c70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h695785cd5783da9935f140bc5bc6f9cdf8b16a0d724799db8803baf7bcaf108d7004d117baabc208faced270f5409e6279392a658f3f2b78ea768be2f7bd5157fd69f04bf1646952955cfb9bcce4f09291d6a96008134f766349b96ecef30d8fb6626b2731a772219f09468587e680cb2725a43da75e34f72ee41cd172fa9ced;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7c69686664193d3d6f40f8e0a11f423d3581659f14a470e19780ca0c1ab6e675e1e6ed490e3eb0ca177ad10cfc09be8794635b0aeaa5339d57bc269f9466b768b5fad159af84448cc832ed0bd527b6c4442cf8a69dd3fae83def405888c9d48d01290b19163920c75a2eb363e327455a74a78166d42869960fbf0226b896ea0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a1b73c93b92e830f11876268bbd105f1499a1acd3a325e9f555da5f7269ba36f8bedcd25c67fde668b017b452cce96f1e05912a041225e8d12383a35ed2e13eb90c7075529484cd226e5bd690a3c29c177e501dc70f43181fd3e36c7d9461cb88c87600228b28ebd69af5d0035e93f148560f5d8e148c6460ce7aa0b44fc80e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae0331400f412dd69d10f5d65d065007863e91c056188b77fa43f01b2cf0a7c5579fc7059ccadc365ff4a23df28e9f65a64f8cb164097201bb51118222dff26d8ac819b303ab0b4b8ff717ae74960cc2987017119c90ba51102b1fe5cd1fbb923a5016b5ed5f5867b61cd2637f88c0cbc890d4e25c970be7834bc15cf92e7d67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7141e93768b905d6fa0c9f890cb14be1db14a14beda770e4faf151d914a4fd363e815639a072334dde29bae7e1ae0a6d1d37b9c6267d9e51d18b6d6756c14618d29cfb1e61c8755ad4e0ceeecf21d9077e9385c0b7f3c2f7cbb583fc5a2b3c1b1ac7d8b9f6018eab70e1716bbcbf111bad63c565a19ecc9ebd2ee1028fd4f680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94e570f74e504d123e460cb5bc25f9248a35e165e225c8dc179c60c593f953b5e5650ec914377db0d1230e402d0511ded03477b637069926ff937fc69c359ffb6cf5fb2de7231c9ee9257dffeed4f13ab16d187d7f73600f6205dd5c310adaf0726b2447ee631f6ec1e3815f3e97da4da5f34e492a748a33d743a5610a921910;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27df036eaf0afb36fb086bac80fd1dccb01aa56fd1d7171df0db1e7768cc82d809034e037e9a80948728a26c0051f8cc6bd462c7baab42994ab997dd1f7049e556791c0cce31e899fd02d8e81d43cd33fc470313209a1e18d1619e2f39869204a7760432249ee1e8fea59a8789da8589d5eca70ea73a2c43cf8fcb856f19ae20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h680f74bbec86aab780b3908837ab3c7a212f3c4b7e1b2ea8affb6ebf50df69243017658f99b75ac05307ee8608d08507f98608a25d38078bd513b49410ef7b0687d3d8c905e81fe9e363c38bbac9a92391a3674d09dc292b6fd8dc9d1b80b6d26479bacf0efea10b9532427303a3974a9dd3002fd7621f9e4d7323d67eb826d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9739ca23cd9ff1eeb039a7d0536a3bae75f2a988e8300dbaedcdb1fa362ad84b2245631d53b2ac69f60968e2c63dc2ede0e193c598c5484fdcc45ac7e65c21b85e71c0ba87d36e1a7bcd34ef08480a4e8943967b280e1164f7ffc170f56df1a0838e8c09e37d5e039cc3f2b6214bb8a1f498ac23052d01304433da9162b859aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'head1d91b353c2c8148925838389f4122cdbeac8fbe0f23e518ad4e2a9a50aa8e422de2121bf537815705bfc59325c5640d3add816fb49f4381734787b002d61fc86fcceccc0f9b27dad09c98a08a98bfc61b8a6c651cc38bbe86f806a9e4621d5195c79406c8e528e7a39b653e699e509fa7ff39c6d4e727b2de4f20f367f00f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d06099e38f934ad0724ea6cb42a08c9c446e9081334bc41a3fdfc4f6f4b5426fa7c46de61a606d131a5c89c26ee56b042c33aec51c7f2e8d27be106acdbb4ba7de851188842f0f4602e81a91c544cd15d9ff51a9679ba78850e816549aaa4545aa3f874a40f59c3705151c98b0da655c1304286115f08a339d63e59705d55e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d4c875a6c9221f4c29727ae99decd09291f2c8f90e796d4979387815ae239ace63581e10bd9331970e032756a756cd178ef809c6019c1c59563ed90f3d303fe567808c4409b6ab7d822d2e604a3a0f23e2906af2d6df34b2366fa139ec99c3c304ced98446766782ae30b53da4568222b3a2aefee8aaa155613cab232b8483e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4a12237b2fa814c114bb0a33c8c37fb7ebe015777b47b1c19fe4ad2051cfb1e7104057cc95867b1666791f4c4eb0074d78dae9dbbc57a1d4025c55f04864037bb85e02ea0ae8882cfa44b84964c6449843e6a021a455429f2dc012f7d8f5fe666629742c9cd80e05ccc9d33087451c093f8b9dd3f6229b94b3b214cc538e684;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47de870c8e5879abd9d7924874d9df4b95ae9c794d480c3734db14416d2c4db2d8a88b8d96712f2e999094d25297b08ef20cdc67a558a86f3cea1be5a4e137cb9df07c9ae3863767b04debe04312efdd466fed5b05837136f93e9eeca9ea6564d5b2d5ba1c4b436605a3931191b72f9bcbe7a212b9ecaa39670b900e8fb0793b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5d6922b6534d4eec5ba41f64e4be7f8f714ccb70293dd1977f654132ece64d5a5137fa8c93d2db282a0da62e45a13f6f48826db595f32be6f59223b770a98547541a234f48346e6c537584f5890d20da74a91d8306a4d6df90e845ef9038fe948985c0e8df0a33bf508ccaadb8320e1760885ed85cb78ebc677f3f7b34c44e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e52209657a741eb41a4d77dc4d2121ea6ca73518b9e605de8246bc33c4c93c9b0ca48d61f53e43825eb997d65f5370c26d09d6816fd2d81034c394e53a00ebcb07806b4984ca4d7b61ecd49300696e7553b671513b124fc86d4ff10d8e2d7d22c438a7c4d29705d95df2ff9e252debda1032201dc449ece36952e5b2a61164e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a3db5209c9d7cfbdd10809fdd910c2301c6f53ff03820ff8a1255bc02d8ef07458a409927de9d9b94963631852313500c93fc86005edfc0f623d9ec9112e1df8144734ac712357b375fb646a7b21826be35762b31b6dc16f7666ff9a46f653729bb337e24d88f7a0bbababf2c643b461024008126d48e147a4be05bec6676d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h747c0927dc315dd0d48534fad2250e4a0f424f2db7f098faa1ef5f009ee04e285aae2b327b64ff71d9c8a2bccfc9958866547cfe579e7e4024f76b8ab59ba226f2af20c95fc09571e7d69e5acd42d99a81ae7d9b1bd18f0e96ff557fa82da1c3486a929469654e3aa4f0081e7d020417f85ed18ea8b2cf552d778a90cca4c4f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ea96a1efceff22fff68d6fea1094bd0663360baf22d22dd9accbf38ddcd6c8e5851bced39ffbc0f59dcd280c9c4f428b50ab396eda650cf373c54a38039945eebfd565d067e303daab73c5c36af6db92b57d66673360dfe211d815aecb49950a43fb6cb8474f0f195d17d3b53fc493e18758f9eae9532c2411506650c50d205;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h553f48e94acf4693788b25200b55f3e532b62bca14958293e7d72a402e49968694d7e50ec495b94c9d06f8a7a0d991d8d824d73e9fe6a1538d5bcbb7699d3cd4e481cf31f2b2a2a33b80bd02c0e794bb4876f3884e814c14bf1f011c92d07c7c3544e475e72bc8b584e7f6179e67f7c85efb2d4cafc0ced40ac64046775f9443;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b69b0bb7adccbb2d5e7f0518e3580827e20675df9ef857fa32aa03dc5470f0a44cb17cf76f41b1c67cbfde38e571b3cecf4a3083a01f9097bfac34a3954930524f99f959a10de988351bcc1d3a3ca5c7e0aae9d4298a7ea2e0d44f0b41d4919478f7bdb50b5a1d16051b46bd545c70a3f1b9a869df570f6c0add2ddbe855c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38d1152f4880fa3ade578ae2e83ebee304370cfd5b18f2ba866cf6b38e1168299a9b29bd44481a3bed239ff88b332bbb90f79ebba1e58e77cb280512c47888280bb65aaa4e6711575f904fa547127a91be8f192c531a4925fbf0b6b339b51f5b515025356bb6f3d6266ec963751cd6343cde75bfc7c723ed55df40442ca0f570;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71b9181b9fb9ec817b25eb565ecc0bb2bf8497d163996ac52c4454834c44eee46e38cdf4a8eb172a18c92ab039a49f09093ca276aefdf846f5840306a5c0dd8a1e4220c650cad8d4c8c7e675bbf5b0a8eaf4ffc10f0800bedf87658240115179c48b5798a13bb3a6787d47bac45523237c1d2530ba10f4f60ed31292f47a045;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfab0cf20bc87952a9d959cfbecb8b17d7b82ffb8e98eb2a87bcf5791c229d8aa68e1a31850738f52cbed6337161d39da6e23b37017fe6e3eac66f1088136a564a9a80be22bb1c0bef7868602ffe4797e25e4185a7d297aebaf4ed3666ca3aeadf4eca9f709d08fdce5f8fcdd44d1465db57b47a3994cea664fd4a734b450ad1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h314830922e53cdf4a3cf34328f1562767a41cd7ef2ccc2122b6c1753286377743a291c5cad21746a033a9e5701a632d9581bdd4f38bd0eb09b0a10e7f8aaf9f546518fcdcbd72dc0e3da8999b3d5c7254a580c1b3585e30c1cd12078c03fe07e4fb0aaddc95df9eb2c6e43d24d6143e5a65b8c4dc765c1a47764bb7960e6933c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57c94aac1213dc86b7068d4100b1611114f4016fd6a11dc4813bd37ae31cc5a8e2d619fcf88ead569b8b9ff65117f183f2fb3474d919d68d42b69b3f32cf045a7b6c55fe7fba2a08b5bbe6f69c96cfde0889c5051bb61c9141fa23fab479c0c5d636bf845714d9bd11d250ad08b378d437776da30a37ba871c49260f0ecacc64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcb7ca7fbab3dea8f94b06e13adff4c08771adb18dab44fe46b22269bcc7987a759a9d2dd68e8773384a40ad76b19c69dc2405a31bfe9728a22e46b814997044b2ef1ec6aaa799a30c89828a920c08d3177fe6339cd8fcc197e6420f777aebea2757f557b706a4156528f7ec502b4d4300764a00adcfea145d360093bcdac9b6;
        #1
        $finish();
    end
endmodule
