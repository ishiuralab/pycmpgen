module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [7:0] src9;
    reg [6:0] src10;
    reg [5:0] src11;
    reg [4:0] src12;
    reg [3:0] src13;
    reg [2:0] src14;
    reg [1:0] src15;
    reg [0:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3])<<13) + ((src14[0] + src14[1] + src14[2])<<14) + ((src15[0] + src15[1])<<15) + ((src16[0])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14eac8823b0f8e7927039;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e7d931e8f13fe4ed42a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b10b9194764a86ba0059;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1622a8084a78c8d1e3266;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d782b1036e2ba60a07c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82d6a2ac3d8bb1a8c76c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc34ff8a213fd1895606;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34b2eac42a3fc94f5665;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1341ae0b0474df29d5cee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1359c29f855d5e2bf8b83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8acb55b2b9917f3cbfcf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58c1cc8ac0a76e817d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h46a0c357d4eb00fe1741;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1732e4121b36d0cd2e233;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e86af72d70ea3b6a396;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e614f546f8f166ccaa0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1773bf41caa6fa5195d6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144cf4ea8b53abaf5eeae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f95c2a415509e24b778;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1672eb712fb2ba171dd87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8989a43b2393dfef73f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb68e2c5a28e15ff69a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a38f2e091d142f7abaab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f6e786981609a104bcb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e4c7987df92bd8fa32a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a66a24775381fb561fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5c5d7a11cfd1f910873;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12021aceedc4b401897ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha361a69348e3f94f7b0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a7abd871b27c69a1910;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167a1cbbb9d64a2033b7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1b6c9ec2df5a3bd9af5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6379531490fdfbe43766;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79ea7b4b10539c16f728;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26563eb799be14a859bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5922b67eeeaef0421884;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118f8f5a1d949a18ad914;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dd7a0e4f21c2626f6c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heef8683ec3b1b3db147c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdd71afb9dd816d2071a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f717505bc0c00135718;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc25cb09291af9ed3b90b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1a3d2131a94c4ecd5b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c99ab37fa2d3613d78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7420bc14c0fbdda92cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e130763fbb4260a12480;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b8f1aeadaa6ef158940a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8e2efe45d50977113d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f873b37de59667b1c0ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he24dd93080661302be56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h293781c47bf9339ed85b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1123a52722f6b1bbddf7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92d679b95e1c7bff600d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1e54fbeaf67527607d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h195de195c3c5d38f3b4d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1046d7a8d223b6d4ab855;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4204ba4dbad18e26508;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4a301e83c2ac9296aa6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h153d970d83d6d550dc6ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d138ef6875aec55223b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128beebfdafb7c52ec672;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17987d4251199b851df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he98774727a0c21717be2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd329891ce142bdc798df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135369f5900d84113efe4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbaf1c5beacc276ffb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1581bd637a5dbd06c7ad6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d9e5060709156a35f4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89ba71d4ea4ec7b3f2bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26b38e5604fc9b538dec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92bfb52d547fda010233;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e70af1fa052104abf626;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ced1a0811c4bea004c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135688bfa47c4d2f403bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150f090edcca1f9478e96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115b5e75768ad7feb1b1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he46bfaa4802a882f9892;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he097a3ed4a23ffb68cf1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a038fae21e6c080325bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0d628e7b471fd486c44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ab26957cd6e3594d373;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h315e165d7eabc7860cf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hace45d76f9696d2180f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8edee40e4cf00c28abd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151e50cc7f980ebbd0b9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe16c8bb815f695ad87a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ac34ef3925116382b45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1346db6e444a703230011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eaba8ca34b3ec0603a7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab6122adf6e00f1f8d72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104e424ff3eb7baa11adc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5f1e2553ee9b6c15f2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2672247c4dc49fb3f509;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3c1aea3991f02a1fe75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc22c03ed5f0692ebece1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113c67adcb548ae711c67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c355cc5c7b56efb1fb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haed3623573c9a9932d2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h327dad24c393369a6ad0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfbf8f688d925f286c75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hebc1c7fe69520ab049d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cb079f3dda49e8d3f7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a665e825d14cd2b7840;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h77d07935674adf648d49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a70c70dfea7abc0fd10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf6d863676d20dd9af34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ffd373c8a039c36191b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f6dcaa77df04e86a995;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a14cda72e247dc827945;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba738b19e29d913f7d4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc39c50d0802c17fe50c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e32ac60b24b87740351;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e44265061b16d4f2439;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdefade26313c2b3dece;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b49a352a633b99cc784a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190636ca21f8c1c70eea4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4df56d8dc0f26f8b2c62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1446f1996f9063f7a4689;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d7f65ade2ba6b12826b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15194029141b43a79f0b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ea47a58b5277255752;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1beb2e5b5a0c5221e0987;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71e3994636829f87bfc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2e00235379e74389d54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97dca7fad9d0c03c38da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a361ab26906440649745;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121e20db56f7225468758;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae2484407ccadd0d53e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95589d6b92dea1bb4f74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h357f67d73b51889a4652;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf965060a24e72a75996;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16624abfa1ae8959eac4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f18a62105a28c0f45083;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199fe87a55158e1d481b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8bc22b22f13d53f32ba8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc04b7bc1443ee42eeeed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1978af4b9d6f2d678;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b30ca673cfaede4d7af8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7be60dd37ac2f43bc1fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10791989b89564b515b5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1acb84b32f55b47921e0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17497e942c0a3d71ced9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108e0ea466e8ee37685f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1f0a3bac45e7ef70394;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc08453a208d61cd9aa0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b003d0567f79cbaae76e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92aeb3b99c5a3ccbbacd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd023dd74dbab3d9e3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h523d7d3da98708c8d06b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6c8f2e08c5f1507da3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9a76e3ef42a24530644;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113055ec6cddd38561a62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178e6e6a848f73abfa899;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec04a6bb610b49addbd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d795745db1a3036ac47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2364f31922576a844644;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha56e9ca9e90333e73e75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3f0bf49327bc1e2137e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3c78572129e7b1e5d1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51179e4e7dd5dbe8b36f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h816d9b7dae7f537d484a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e70fa5791788d057a486;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1639726c210a0a1f81cd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e72b48e8e4252f4c2f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af8710a0190899e116b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1540aeb94da1749c8409d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf81473a25f743ed040d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9c9bb611923c870988c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7e961b07f40d1cf73ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6119fb30ba20db3c0f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11439428ad44f2d8fae82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fac0303aec80e5ff1a8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e9d2a80bf38261d8a44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab8f04baffe4e55093d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106c8a77b49ec07c12917;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb436cd47936bacaf598e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf591411a43325075f105;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2769b716f8795c6a35f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f5d7a9803ddc9edc82c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcec8f0115f61f966fbc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h243cb997cd8ed249bc64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ba7eccac1f61b8c4a20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dce883fcdbfb33c9d225;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b6edf6e03a8afcb7692;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5880c37d7599c33ae4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab4728d7d40cb5fd4692;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1342bdc45fb27a298a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fb6691f16bd1fc1ef94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1708b378ce8deb4386a12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff27cd746096b2cb320f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b9d0135c27cbaac8024;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19be4aef5f913b2c51905;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1f51e03c43ba9e30bb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b82c6461afd53cc41ef7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1128669b00572360b71c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd97c372ffc6e8faa3ee5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2009d2d9bdc29c3f0a51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8baa4102aa7f13b8b9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10dbd9d412f71be1daea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd5587de8a11d137cd97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2de07ccba3be0ae1508;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc1d7d11dacb5bb148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7309333dec952b934fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17784d392f171576e49e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d410dbbe6e597049ac61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8bb42ba5062567c49c16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182c85ec0a7a1b5bdc5a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fda954f3d0a8ec1a96e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca5aeec3659280d48126;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c51c28deb410e130caf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h648b6cf49721b6eb1077;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c42816af45aa18ae31c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1797901d01e2b57151918;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde0727a59e6d4fe19f6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191db0722fb6a2205ba13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a36d8b9023070b445476;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f79b6029e5a58b664a74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30087c150068d70bf63b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heff774943051f6c0d6c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bf8aa8522bae1500aec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce0297ac704b8af6efb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b870964d0fcfbde0c26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c916f32fb98f332c246;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1075b954f7f9420b83237;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e49b29947d2044a246;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e2f07e856f954bc653;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139363e439a67b90a27e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4ed83c8f1750d1b0989;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a975ee569d385d320f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7054d7ef8e1326a23b1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h879cf108128461db122d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7174e22771fcf8259a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f8abbee247d4518677c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9b2509bb87e16e6322b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8b2e12bf8a480fef54e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5acd9d579f72316f30fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a01400dab7a9217a142a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62c4ff0dbf736df4e351;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33b6a8098933cf72550b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa7fb53e9fb6040efab5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12420889b4f571fdd49ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c2136f605ca45a8d8c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de4708f5058a83b4060c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h253b98e4f5968f477e83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h591293227446178e62f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66afe8f6bf9479fe1929;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6165c8638d532d5a5166;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he31d780a937de66be65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc42ff136189ca59d6576;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58969fe88a3bfd280baf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e9cad8fac55cfb13c29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbddcb85e71391930b7a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7b4206f3fe568abbd62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h243107412e393661c6a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3cc746257fbe82887c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eba24f58a92456cae6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10904b85ecfb5771ecf66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ccb19c1378aafde4f7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdceba9e3b4a00971b380;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b44911a9756f08234fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60fb76c14f44c53a273a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1057779932ba07f219dd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h29f71c492d8f544b85ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7262bd429132c25978e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2713492ddc01fbecd8e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb62d09879dc991b9c2fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c16bf11f91f4d951bab0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbd2613165cfc720bef1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1567516dc6e3482b1829e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f7b8de74203bca362f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e4d80d5268b56b373c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb09c4ad8e0fc9c0fc1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2e7d83c57ce189b793a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156b8b50860e252375640;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h551d62ad8615707021c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90b433e79e4e6560cbc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c76f94caaaf10d8f589;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17809678cc88754a88790;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdf4cf2e7d4ac75b479b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3bdde11aa4cf15fd926;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d45b661f5732c630c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17dba1e56393b1f828c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89d0e3e34a577f1aa5b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bd9b98bd113f9e28a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189b50fe60b60866fce4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177fb614f8c63a7db996e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf17186f42e217fd3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h597e93dab58a0299344c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbcad0438c64d6f5971c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1515dda13b735b56d90e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a18c7cd64f8ca015e9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124eea414796f717342be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147b4aa4468a4ab347db1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11689549bfc71e2eac715;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb979b5b6df388e6e5a1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8ca4e07b7bd49ccbbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd421d908e2ad6056def;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0aa5c379cbad39f2798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20f5f2d71d255276f4bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f172952665395089fd99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h828aca059c8760f5058a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d571c47e7ffc629b14d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaef4487be54f0f7b7bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178f6eacf35e6a98f0208;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36fdf9556f6b25473d2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33430547d7534c44712a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h955cf2019985c5fe2fb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he99e769cb62c46b230f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb3f5338dc6fd569d9aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e056e66a61de02c1b095;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1800630ffa305759ec690;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aedaf5de97eefa9f889e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf88d3ed4d6d1c45fafd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c771e62c10d9eb582f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38f7f1261b0ce832369d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120c22eb297c0e642aa1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19eaf232d053d6fbf89f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac15fdd66c456a27237d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe4a30fd9cb747991379;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51785d6617064618648b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf74e921d5edfc205261a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd5664ecbeaa7185a436;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2effcc2ab21517a0bb20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f65d291148f58e323ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h915636ce42da9251744e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d22144f06b56b52f9a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159863b7e7fa24dedb5d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac834f5342dfc53c938b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha31dcdcf539c12f07539;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8f4c78bf943d41141ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13bfe9bdef4cb132857e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56c6ed79b17f00fcad39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9738a0b9bcce0671ed7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c9536ca8840452ab88f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107a25d5300612f9b1bd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b91d0e4448738d0b266;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1929b4da8cdcd4e17c26d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e732883ac3d88a33d507;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1067037b42c0634854841;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1639a42878e8f1c80624f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6f2717e7b73b7b0b43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b1c397f22436e460a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbaad2d9d0939f10697b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c4943952d9cf2af4843;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af955dc61fd40b1392a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e772519d4edb8d9b7f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11028f373de3abe130888;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e97b1fb70cef1ecaf25e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28978e5b69622183b487;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c953e0dddbac768185e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110b093edfb3629154cdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b84fc7c07864baf55d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128ed857282c2b9533dbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189def2d1f71ddc9347c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83152dd7b3105a5d8ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103dfe8627cc681f16770;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8ab5c7b35fa9f68c33b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161d40b6c5c95d21ba874;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111255f2521867555dde8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18555dcab27a2602cb253;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e108bd617287d146ce2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe39754c30e6b77a23b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1448ef4a1f5e2a80e327a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c52ba3ff5fbd2d5dc04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb14f8397d49d42ec50b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92b97346c997965ab41c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae1f8b1fc6c2f61c6986;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dafa999771aa46ba212d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12aa7f98d2a7010039d3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd4fe687e4c978f6295c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h690a0a709f14798d16bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cb0fac6ac49eaf150b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha62c8831321ec0da640b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdca4267738ea9b1ace2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34d5af0cfd7eeee55233;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15239c50cdcf77f5d9826;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5091f556a5f1c6df83b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d07bbb448805103dab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7d011512c85c6f430a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26c0496a19f0712f00f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e87c592ad1cbc3fd40bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14de42a64b8b82c3b0807;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c9a117a34b8131d34fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150dc28c3dbeb3234e5dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107251424c5765deb0066;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fbef13cda0f4aada74d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8c3285028c89f22d0f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60fea34873928c660740;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d61fbab5241c587f651;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e93a9d1c5015c333d3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e5b6efc393d672638e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb4ae3daa8feb1ae5826;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha411ebef01ae4b6e7437;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6afbe43e7e280aad75bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c915a06af872d889f80b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c0b443337b9bba26925;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a55fb0234780c83d3657;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3af7115ab7070e60243b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a555ee3a554c1c6c10a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb79284120b6f470920d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23e7a647480ea22767fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b7bb62912a4ef3fbcf1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187757294bf6cfcbacc3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1e09bbccc1df322b23a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19db4ad26baf9e595637a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1120d4662231b687d06fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b688b7e19dd971170a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1820826b6c7b174ac40e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17c3923e551ac194d36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d7c2a7b6c2b519974bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bada3cd51be7c968dd1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f046f0391329d809de85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b48f31a188f5228b6f99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175d4af6c9ec78fd80ce7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec521e3ae270a679a7a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0a82991d5d126c46490;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1907f6c630d395eaff019;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h913e09c8ba9d5d13ab5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c53cc6fc304e784c342;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1879c5c43d355e534c5a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8119576487e986ec88a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f36051a798e55e0ad672;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d6fb5d10cebb80f0464;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a14d2e9a49733686f0a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6c18c2c0b2b77b16a38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc18730d3feaa80a4a52c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b87bcbab0a01887c68a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88ccee4bb3a3d55150a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6d3c9b93f9d989d5d5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1830acecf2103da4f3ba6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33258bb740ae289bcf66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10250b47f81c0c991bba8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e1a863603cc52104aff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd591680b20e84491640e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1369bff0d64e0ccedff6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bc690cb322198fc4ef5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d88a29f4d651f666f4b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc2619d21cfd0874624;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1a46fbf2688b3b9753f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e88c2a6e84cdc9663e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b67bbbd6d9f4e40ef895;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d49780645eb021fb7d8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183e32569cf99351baa27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113529ac71f8af163e937;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4206b5bcf3991f644622;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2bf919ab8d487ee76546;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cdca19a5ce79f200a42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefde70cb29af1de98ef5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7451600a85ce05c416ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c1b6e4734cf453957b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cdaf9d8009c123d2b85c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f06f3d95d46ab4bae400;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ec1fa03621fc6408a3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f50e2915884ddd41f587;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1716ce7a790e1b25544da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h335365f3b0826fb5f22c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19abb097c2dc579340175;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9fc2e29aace2aa3afca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c81953024eda05001009;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140e3de3d1b011aa066fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53442efe62a85a01c542;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c573e10097ec71ef3e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b5bba576a6f686085c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143f3c2b47a2f2e7e1f24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3aeae18648239d59f41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fdeabde8cfe8eba3a6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd031857245f593273;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb37afcc10fa67aefc893;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he924ad54627336c2f8c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b421ee407fb41adc082;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3e3e29c8e90b23c24bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94152fcf82b8189c1338;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cae9183a32c6686927ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cd40ffb46857cfced81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc792dd0f12cd8502dc30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h420e4e98ea2ef3decfab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddf8f7b3d86f2a130ec7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117a215f0b87fb87e4ee6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6d54086d29bae332780;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12124d40fa44ab9915391;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cc917be52c707240ac5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1851fc475a69278bd3f4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41d91f6a30761ce98181;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a83d1e2a7a7db6b0cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hebc00df74934f18d4c7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd35e5de77604574a232b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151271ed83eb66212bb7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c2b9d7166b8b3179567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5679e607137a52e4b05c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12832c5e8fc8c96b4184d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9287fa3948df625dc12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186fc15ba8da14db8eec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d4bd55f37024ca23cc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8fd47b20473de58a33d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1873084459ca08b7a73d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f73666cc9546eed2674;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20d3b5b531ee0be402c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114275f49cdd329b96d45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c3428ec207bde924324;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6b1862f42270c2d6e42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32279451b895263c933e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149cf9fc54e8997d1521b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce634b90ca59608bb9d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159c233412c40d3324a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c517bff8850ddd88041;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cebc2ae14f4f8294b06a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1512bb1fe885c720fd89c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d1c0d93946d5c413dbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3b9deef4a7644f00f07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e41b8769075fc57608e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ea497f4258f5c4b3567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140aed346dae52cd72f87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a122b848198913e8de8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21440e52f3694cbee988;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d5b5df0e8ca582f8cdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94d3127cd3c23f403be8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ceedea47a199d6dad736;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eca50c712c2afb2fabd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee071b775483747a8586;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f5479dbdd3cf6ae0fb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef95b591330951137db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6ca003157513484ab24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2d9fb6c15af0e4509fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39601950d292fd036134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb86d089fc74f882d2a60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e551305075b4bf18e81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2d5402e1f537b869ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1660d146ef5943b0b83a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174f0312d4b878c3c29d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c761aa70c00245df2b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de2e729cb9dee07eafe3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8af74ddcd5e751088cdd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6b8fa7d57c11f02bb26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5666321d9cc8893199;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1240a0bf8615db4df4d2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he577de59739186e3ffb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e4a6206ae2e16738b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc20fe395620926113cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d49de5397ab85162f85e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ded0462957f56f9320e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12492b2c1949790603f0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18804192c2478e723dbd3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b5dd90a7f399f62d3f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cdebaf89ec5153f4a24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71bc7501eab0c2908d3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9ebd2e6d0b7ca2f574a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2cde3a7db8aadd5b472;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb40adc3b6ebca931e99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10515bdd53fdd20c78343;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h861ae011e9875bde3391;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6e81219507e81d79cba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130ef2b3fdde03c24dc28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d114e96833252d790b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf17a3bfaa3a212063db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182fbb9dcfa59418dd5d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172405d41a33088f2aa11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9b51563dd333565ecd0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9e011fa61a94d9f9a88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cff3fd1c477f12bf2cce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89bcc525b4874b537dc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb060ce612a593e14940;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176a6e77471499c8a3ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a39406912fef620c71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1109c72469f1b20f4c944;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ff440d4a0adefc6d181;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2014ac282720e2603e39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1595325659c5c20434e79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda3acd51b940652dd218;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a64f928d8e4249b17ce8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2b1e6c32697590ad49c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde15b571ce5c3e0ec36b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2aad149dee6882f13202;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179c263ecb956657789a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0a998fa0f3bfd876d1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140eb987c86ae733d12f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd907b1b6cc4a7e3af5d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4a217f1e39e16409a36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a73ee342efc8d1f08ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14870d73db532fc542cfc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7d59c05e0f1094dde58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdddb1acc561219a8fea0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af071aa84fad0d9b2670;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1abe35de2b03f3687274b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e79fef9d9cfa8ba2245;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4928390308cf7d338fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7d1e9cff7538ac571b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2dafbc1f347d340c6812;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1c4a3dae2a2f495f885;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75e70f72389c01d9352;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd442d2aa26e5894e84a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59afa11ccc155d86be7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1554f7d3d9df9251e66c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb02c468c54ea53376d53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5232dfc947ab45cb31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1352fdc561a339852066;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188d97437bf8f1a1d2bb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139ddfc2745b3b2052cfc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e892ac147f99cc7088d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h539cde72cc7c27908a89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8db85c1227b23c3e0f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148876dd10287e346b206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd3451d487f3176e4e68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172abfd75918a040c9fb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c5de9d952e2534ada1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8bb2bd138279a8021ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2256b50668b2b5043fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18215534799072e42d8f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf2227957af6e8c47953;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1535fe191591ad1d0ebb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd6683d0946049dd1fef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16685cf1c8fcf422d512e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129769950dc749ce4afbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6f5e284ddafcc2e011a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16257d7cb239c5dd553c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17290b12d02a022a7c8c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67e64df9a38eeceae08c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a011797ef3581ba235ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a0c024051f3d4533922;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a291c80964aa59aed19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h277ce7b90ffed99f1fb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf53118655b136e591c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb93e7592a6b2ad0a4564;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af329d409611fd160fcf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be91bd824ce8e82bf74d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125a8376f34c07d9a2671;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7bdf006275d669564f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd14991f89234b50580d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9aefc886716997c4a8f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c568247f54a3f4678df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h727311447eae3bc3fc37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe78800f1864fb3b462e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffefa1e44509fd7af95e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h916b7fe9ac091a119289;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3c1b64f1b22f15ff0cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1621a09107cdb816db0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e7d47d597ee3f970fb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8c3176b6f37322b48c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h697be21198956d8114fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e309c909936e11477bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f9a2924ad02c8e86181;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131ae4835d07432f0e24b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5d1b1d7b3a19ecf3a1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab5025e216804b7c477d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165eb8add6e65bfd98b41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa031492dd7277da24f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ccd165403770fd8d39f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a07683978b85de6450b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e9f08d0aae67d995ca6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb421a6285780a130f14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbb27aed8ffa0c9ad5c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9d2b8741de8b555c19d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148496296484a2e7a7963;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef7555e18501266ee114;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec9aeae3e49fad749b89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a95dce7d4784395b8c70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1bef22b7a738714d798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af69f8f7a283551a702d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8f87d9cd1b1f04530d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h91502d6dfb5e105a7964;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d904a1cba5e2cf62409d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1062d2ccf8666c9176816;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bfc180e28b8a2573587;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4743246e46c11db1bc23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h306c83d4ebd1d1755650;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d869673bdc7aaabbb31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf42af2389de7267ae6fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13270a363ef876c9c918c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dd09edd18171eba9810;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf43139827a44e7343a48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134301964364196ca31af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf64a2b4edc2715680130;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd22dfeeb769fbaf82cc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1abb990874408b8f58215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af6d357468912f680b40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h601a67d947b7f87bde86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa11674e358347f2358f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f6f63582de9cd6e871;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154bc8e81de84cd5a5255;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50aff7d3fa141e0a3fa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139358ed6b4ed248e64f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe11d32118721eac5c47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d71964a0d5f3645008cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6713389fc64863cfc32f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f85a404bfaa4b12840eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d43c6a978d8755984771;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6258552fd0eaabee4f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb76b20cfd27f7d93dec5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158669f26494c52ccdc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc423bd97f9e733101f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139c081c5e70d5fcb7ec2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0c7b467753471fabc15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e192af7a56b9a4d6fe8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85a49565d94b40763ef1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c095941bb11498b5115;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a7ceca07afd3ceef901;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1999024c44c9057abde16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138bdd26bd670b4bed993;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1603ee40b2324a808d148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8445cf34dc4f245b7bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c66869fc85b6cecd5071;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7bf2ce990d9669554cad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafc065231ddd0c5a643c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5078bfc3672c1c91d99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc947e687599cd5add46d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73d0539a50dc772ffc14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57f94b37d503c069221c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44c58a5400823becf4f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2b3d7ebd584768f0628;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d76dd9dd7d7c7fae24c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9eff740d5f14eef27a99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f8fbd16fa5b55129852;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd1f949efc8e0590a655;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a021d5f14adee547d7d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf748c032a4a3f3aff6a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4d9035796a899bc1a6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5688b89ab00fbdea88a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150061d6c9118953306d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b84b1d5857e7a8ba1fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14354841f4418dd13d4b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17bc2aa430cb2470ca2ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4ace99e9b2a4ce66c23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128791d4dc2d2400ff08c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he40c136b854423691b75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db9bcbea525b0a920cc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha16d72b2aea86426fc01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24e627dfb157e90f844a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c63f75c893e224d890;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100291bf6c7e1d208456d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db0778298ee7d6d4b4f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d2635813efa292ccf4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c340b084364fb163f3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116a8e6c6778dad07de47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd50e7760703fe6a42c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dba49bf3cc6887f5d733;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130853ec81cf1d55d71af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d8463384dda1b7cfa4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h63f4454244ae9c644e21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b11de2cea1972457fd4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf52429963cd9ba8d89be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9ec55f6b8b0a0dc4419;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e27569c19d81368ec7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14722a3db0ab379fc7a6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b17b168a9ca74bd2ddc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76c43bd25d81c05cd14f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3afb834b5d77ffd7fd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb9dbddd53c4da49830f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11317207c24e3d0c4d669;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca9ed4d10417f83e948e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141ac9e86f2ec84d4fc08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac2f149037f7f9a0bd80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1120a10229a720f6a7b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55aa1b487382a4e51943;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f5770a7f5fe6e7c1417;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afa04aa4609c81ce8d8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbf96853037c6a094144;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ad2837f78130a024ebf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1496635c71ca24a1a6403;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h875b5637849fbf92119a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb473d6650aec1876f50a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ffbb008132cf5f6777;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152baa4324b01f8491590;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec8c60b3dd6381b26e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7539a70f361b75d2d148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7d5fb65fd7daf0d6a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1904e3f2cc6d85ca4fcf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19798e0fe242c1921bd8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155f3ef9ade7ebee68eae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d70568ebcd68de5ddb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a16b6f40db983442f33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c6f66b21a6a77efe0bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150a0a3d4130ce0aba8da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5ec3f4f3336458825ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148162ba84498b7e0b48f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a1393cd5fbc6bb0e60a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c1efc0acfe6bd7dfba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1657b6a09bed40d61bb66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1255ad4f76ac10faf619;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdcbb29bd89facff8673;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3ad81668ef09f36c18d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b6af8e73817e68bd102;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115ca2ee0b0c31a3cb10e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148747082b9a8e5dfeed9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f8ecf14bea46fa4e8d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c3e2743ebdfb1318266;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2228a8d6677ac2c7831b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3138afbe5cd6e7899c3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d051c98e43b4f59e5fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a844b5a6ee1052aa55ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4426cdd3e0078477dbf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc327a9bd2c17ea607a4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16db79f4f9238f7ee55a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c67ec0e22130be2ae6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1411c0d4129beb8c28e31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e80ee975037993a7245;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16615f179299b55f61972;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30b65ae2cfc8bf6ec24c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ad589276df7ac58f025;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha553853835c29f173f90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141803138057f92d096a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4e1de7a410a31e174cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b71119d64fd20b2d1e3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ab26a185557651d0100;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd50d3423057473be2ff9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb73e328bd109fef4def;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ae43a81ea58c950c89e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ddfe4af38b636437f8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185b6cdc915120f584d06;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186c167c6122cf846504;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e6bf3a55032874c88b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14cb3b07173cb721cd2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123888a6a7d0237a69afc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd39625f934ce89050d33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0952a10550edc2a80ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a627e2ff5094de9e25c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bf2461e71786155978d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173f9abc72140270843ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51129f7468d8788dfe8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14bca876ed34474d7babb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44ad80c524fb211deffe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fbea40604d95340c9a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c189e22075fa136a4ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1821a99265a7943ae02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1993f505c8922af477623;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b105efcef6261f6e34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a7c3c1afee3a9254331;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea679458bac7ae7804e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107ebb261bce9e5b08e5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c0fcd51b3d878253760;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h895f202bf348f8f29a2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h563ab75d6a96ea1de544;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1e95b7500676ff3d805;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb343c8cd1f1c0ea0d4e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4ee5ce88c65286c752a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25eb245ee9132fe45226;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12746cae37d9c11376f8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h524b850752f6e69c3aee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d576a0832e2556e5654;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aee4d1c4084903cf6ae3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fb1d34726f59d9037a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15dcc215e3bb0bdd68f64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9c261b36ef6d67eac55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbee67aa37b6d42b96ba8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8b9e6c1997afa75ad32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b14fc97ad3cbcd7419d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31ef218c9b0e5a426a6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148402d35fa614b6a19fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7e992f112ad96ae6baa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e32fb9fbd044ca0946ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he60939bb70af1f80a4f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a489c80fb69c2ff4d080;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13bf4fc47b928b9b2f59f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7607b7804f99663faa8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e146590204b1e9dadcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14142a95dea70293fe3e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd14b0763e6bba0b9dbf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1874a532dac357fdd2fee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heabe25134faecf5893dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb50f28744c9597bcb8fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175aec741dd02bdf72857;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f3eb97bd1bdcafec940;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffb0588914d5ede44268;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98dccba1ec7faaf18b6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16276a396db709ed36c79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b13ccbe8de77d2b0805;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1677da3333cafd000b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4457a6665922c77df775;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1567a75f19aa380bf00bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2a6a090fba6fdd9400b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c15daff2f66b5cedb34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc69e6c1e83a009cb7f2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118a8e88c0b57733d88fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1222a23cac9cec88cd06f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11671d9fc50a14f3d793;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e13fa612aa3d40d80264;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c726080a3098e4046615;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1b70e12d210000b633f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e28a7ca1bb2c457dd3ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20af506bad01247b5a45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dfae0f9de1873c32efb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188ebcb5ee295576ef0d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2924732c1264b5f4274;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e032c90aca718937962;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107b9782efd1f95d8b06e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2234876d4c54134bf6eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe7ad269b1f02e399967;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196ee6fc85d86b02f5daa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18343271bdbed8e8be57e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7e289621afde4edc7ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ee6953fece2b95d40ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6e959d1ceace9c7de40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ee0d872d5c8bed914ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e9175bd7183e8c1488;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d646d2bf075f92711e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1063ac5607195674d20e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1804159d3382892075a8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54caf10ca427d22c4061;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6955a0e52f0637af6acc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c2689c9badb43ac5b05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170f471cadaada6d90877;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196b2b831fd316598a64d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc03a9c775b0b738fa1b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0d7641e4bfdb6a5d813;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h581026ef5a42308ec04c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99910c129acac352f844;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b50dd3aa1e5e86c96c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121f216e91a51627c083a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e61c2fd47aa09f8f955;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1169ac212db675d0ba311;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b40f931e7a86215b230;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d7aebad73a4491ce519;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c19bb043d442d8bfdaa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fcd8aa85306f2c6234b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75017279bbd516ae00a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1147201dd68b5a64decd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20a72f9dcb616bfea321;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12373782bec76e4ac5ad3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c7c8208518ce802a113;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6beb14b9a3bb0bd6b4a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d982941e3f248059ca0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97da88b2e03cb2d64451;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1705524377f0d35bad0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4b1f111306fb10e7b42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1188b83ce594215053bbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13be5b402512d69165f17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6e081a87ca201c59e8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188d0e00d600170aede3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3e641f7a75f11b7cee0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f28302fb045c20425375;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h954e4c70b4b5254b52f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf78cb20110d8cb075eb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7d9c8ca85752bd6d8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14cff89d3d1324c8e8c9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a341c5b4e853b6b8bc28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa7ffd31751a889bed74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h240e4c8d7a808a69fca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25449e860e8c3be71433;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h753e4c8eb60c083e1e6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3e2aa7d1f230960a4b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d4abe207a986876909d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb15ec520e6bd6ad69e02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa7a87aa5d967903a546;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1a046328149455f2cc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfee18c008df7f23f22a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ee9cb60cb314ecca20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1226e30fea56d66eae1e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e8cd5bdcf3b073431db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11796700b8b379f4e3a46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f34f44d644d6adb647c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1759113cca0df25150c35;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1782c072ef75ebbd91418;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62825a3e8324d2418370;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha72e76f4baf0034b2643;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aaab4ad776295bed5471;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db90110cb540633aa878;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38084bf476c8ce4d3b3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10feed14a9f880220f807;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55b738deaece3d2ccb1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ffef28b76500738915e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ba5483e13d1a544ffb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34825cb0b65078941667;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1692556c1ef4cc40f1ed1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h504bfc6901890b971850;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e7271700e76b9cc6571;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d40a6bfb1102e8ec332;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8dc590d901c8a6cfa71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a18e5a7667356ac09dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc33aaebc3ea668168879;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf013a0a2daaa2122f631;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120b07d056db0752026a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha304af7d7b599bbc6125;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1654b3746503cbbe0ef51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ee56ce7de87b3830033;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd44a61aa0e40de31a78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0f279cc8af62ce8f3c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb52c0740a0ed98f0b68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66d5b29645665a8d541;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ba74b9ee5c514a67e71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f2a97fb379a478d8148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118683c267e3faba7ab07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c11883d5aef5ee525c77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc880500d6555041036e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f64933383c4915d63f83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101c654987f5be69f629e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae013098081bffd0461b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha38711a365775e4b0487;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114f3c8d307f30abf4f6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbeddb70be44c1ad6b78b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11492cfa983fc8249bc98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19809fec58017e498468c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150603787379450124168;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17fd72dfc5145400e1b60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ba48c8b3426ea233103;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7712819012856652590;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd1c73c9216a2bbf4dfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c64ef0c81c1ebf542f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dda364910e4ceafa6c39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7967076e6738b5641e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3322ce9a41f9197140b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e75ee7de6561ccfd3b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11bf8cf0edc5d63e9265c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163c56e47552b5568205c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165c71ca7334239fa5cde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f6c9d5985e635316a3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ea6c9ca72a00be59cc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158cb41a6ff6768d0ddd5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe58e84056d79c3b9418;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h336117169f95a58f5427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd492eb4edaf896ab270f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce1802bea5b0ffdcf1d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfbc33c8e50cfb2b03eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf046e908774eae9f7473;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42c2ec2fe789260d2c78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1820c322f888ba5218e86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h997a20b200802bf2964e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1484e4bdef02587220d2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc06cd077d95c9ddc0b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1044196f211da906821;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h839421d8054f2bacb189;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h400b91430cb0caddbce6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1278bef7b678adb679fe4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc273e253c19e0481971;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac071402cfce8064beb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100857cb7e0649a46120;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d98ad293ebd7e1c1aa1f;
        #1
        $finish();
    end
endmodule
