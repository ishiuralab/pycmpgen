module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [17:0] src19;
    reg [16:0] src20;
    reg [15:0] src21;
    reg [14:0] src22;
    reg [13:0] src23;
    reg [12:0] src24;
    reg [11:0] src25;
    reg [10:0] src26;
    reg [9:0] src27;
    reg [8:0] src28;
    reg [7:0] src29;
    reg [6:0] src30;
    reg [5:0] src31;
    reg [4:0] src32;
    reg [3:0] src33;
    reg [2:0] src34;
    reg [1:0] src35;
    reg [0:0] src36;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3])<<33) + ((src34[0] + src34[1] + src34[2])<<34) + ((src35[0] + src35[1])<<35) + ((src36[0])<<36);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf90e358009df81b4af16caa83ce4e8f22f03092524fa99c8adfbdd58b73e9fabfc7eec8b58ac7355931247e17e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31ac603fa373d0a2ea201163852bf130b0f9671d345df062f66b9bcc52cf888627c6e99f9e9b42064268f2bf7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e69dd82071b05b75241efd23ad7a1933da2f2e4453bc38b03f8e1b828d57221513cb1d29269550660d8f86cfdc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4caa749b00bd5e8a2eba1b6a215e8f05f570b143070222a472e4f6f65e1b77f4739dffd71a0201a56f13408e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e88343f9577f486aa24cbd267c4ab5ea9d5e96026d677e336a77abd740a9513612827e477540f632cbf4110dd3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1706c4428dc9a47a4ae241a79be99cfea7fe4785ae8d8fd62852c35022c13178c4a7690cfda99a6d91835d5bb6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e9f147a318228d6faa55c04ba5793a5c93ff007980b19f87cbbd755a0373d51420d0539c8da33bbd80bd8e7fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11806b4d1633c743149a086d7406e5c32aac6567ee7c82cf0b0c82b905d5f5080823dd37d82c158846d7e3bd52f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90d31bd607a53d240e1d3145eea3440bca9baf2c1b85a0b5b51bc1c75b5369f895c29377e1cbf7b1c29d856652;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf01b538302996156546eec289a36c4d35b7df7b0e7ea4a0307f0737db8f5d5a91576b3a364f334d3ef2279a664;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2ebb6dd4a9cfcffb1b9bf70038313eaa927907562c8ca1fdfe306edfb7c09489ec7dbda8e608dcf16aeb863fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76e05ff956654be1aa509ef561cf95729ae4415e84b3d417d349039398a410b00ec54b9b690c5c7d11918eafba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38af504b5feb793c8496d0ba28dd69cf7eca666715d11ecbe9f58914443775836a23ce293df440a1e0b174f7df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff4f99534af4755e38c3565b81b6bff24babf07ef63bd035a16cfc87db7ac4211a2ca9ecaa6194323d2d31c162;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h600e3ab9850176a4eb6674a59b9969037ba8d41d2890dd5b65071a520c2c1aa245aad6343e335f96e3debf13da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189c52735148ae2dc02f60c219478229b97a10e5429ffaad5a4aba525ec6a58baebd9baed75f48cc09fe8fe92c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a3b0894deb4d9222ba48611ab3485dc757a8234283d0d5e99751da3ea73a5e5aa3f0402f4ab1b7b6f5f6d5376;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154be38aa135482d540c77821b6576e4e2c9f2cdac3a80d7d3639f11073c2a373d17b5224e0a36955d8048c29a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e059b29a95335c57a4118c8047d4dff30955d448a456131c455c516d9389f8721309e02c9d1eec367ca06b5f50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9cbf7e25d2772ac9b35a57b4182e455683ddfb259d1303d51e9e1512d76c7d292970eb125f16eed621470dba43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9be4272a02533deb87ef9b4bef42c6b9f594b2f8caeda169b2adc482c3df8f9ceb3e3f4513a8b49c25fd6c5d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc87b532a971650611cb6cb47c848f2d4fffa4ca2765ad11b72146d87835c2d41e6ffe8bbeb9e831c3d2ece37db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42c8a5bc1e6ffc5797dc8699301983b957ac606a9617897393d6162953f74bc82b8825e4614b07be3223d251b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1217e72378d5c4eb24ead870972760b5e6a373a284426c2517fa9a257b378f5d9de3c813e1ec1def90dae171610;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cac227d4ea3d52e18d72da8f28694068e20c6fddf976f2e57deca7f5de63ebd459cc68f66a1ff2a1dbdc17cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc730d7c43943bde8b00922ed4c082b79405319d375c8bb5b6ac22f4289e377e37c43d0fd1a5e371a418ebf27ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eae4ccc4a848e2fbacccabfff37585fe6079537e3322e3d400faead6a08c990137da6d552fb45b6b1ffd5644e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41e0c4b5e0d0ca44dd205530921c291dd6bb662aeb29f91e9ae13e240e102c0c7679eb472853c645f7368e3bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14222bb3903c437ba6270469fad520a1912c5d44e1fc96ce15fbd4a8b4b26e1388641dcfcb2f71a68ea480a8754;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea8ab9f4183b210c5125c14f32b86f87faaf2538692795335271c3079c0c692e6ede11091fc4297399b2dff699;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dd90e95c5194cfa6372bea26c2057a877d612c0e4d2f8b5c5361bde97415ba0da7dbee57017e3aa343729b5f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h488bc4a88020394db3caf13935cc9b4394d016c75ba224ad6d90672ce0d8e66c1c204a98ccbd2ca7149d618f9e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b4d7944b97f075ee7060d02d1424989668cf7afa279a9cc18f408f4af425870f80af9d604a89717bb5d9c146;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56a8a03801625d69b061051e0e11d9dfac75a12d33acb69e71fc69567031d330a7a936a42b048d77f797824fe2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c5ccb45c29a7650024961e9be7cc70d13be6e514b5da2da7decfa3c45649757abb4f71a49ded593366b62f4e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4311888916199895e247f7c5b269bd01212341e9a7a335c256094656080c54f3cfa0e932c69a34d4cbb3a81fa8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170e01a7c2e1d567cef9ab8c4c0b1f15cd5149fdf9c1d16e57f23b48e455a819e5b64a14c75dc747b810dba3b73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9f8bd62e4b4a0febc22c62c6135e71950b7e8441c84d73152103572ca3095625c68aea74d34255a70b698ec9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha113e9fb030c4395fc5ec5babe236133f16ba1d7cc8dfe1392551cae4761b41dfb57134b9d19a7fd67fd7c39d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e52a34a29ae9b1a96b68f7b22bba780f29ea4f82f00807932052174cc4c51e9a47359308051613b82ef80680;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c88f2d086bfc8a1b1ab7686c658f9ea603678477e7b7ac7b71b98b9a689bcbbb1ace51f710128810b79a89ef09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1152719a8193c3231cd8da0e8dffb07bcc7c3202d00f3e9fcde588d9e7cad09fb0c8ae31e55c62ba04f21d6472d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fafc286ec761d5958a90c019bd88daecc25bdb167f182d1e983db0991b205b7b617aa44c39c664b15d85c2572e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf94dda2fc7a1f288cdc8fe301398f89444629b7c3fe1b25e7cfaea7253a131e9d3fd8a486c37483a49e09d831;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85c2bebe061176ea9433cda89950aa21f9dc264454203131cac24295df6c34160fc5361820dedaa864c33d1ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae1084c593a07418759cf51211c93f5c29bf6be6fb4aab505ccac35d3a937fd360e667204fbd9cfc073b0851f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd65b57e3ca5753d365f34805e466334880b1d452fbc568a4a916709ec065b827fff9a93e8f326005cd78ad284;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h941a1bc4e3faf119290b9883261a4c7b61ab8397469064925c99b9eedf076cb0ce687b58f2cb214e7cd34dcb52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df4ede8f5e8c0fb6c96b95ec7404dccd6704f28ebf92c4f1685a58073c89b7748f193b6c5cfb0657e46d32bb35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c84b5520002105271605b524a36843e9c1f48e8797d2c2325a479941f95bcf4ac060d69d987e492cdc806a070;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he072780832906677686c96fc7ec478080f409d4bc947babc2c0fa7a0d907fad83df6726eb4720b3957c15104fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf111b2ce9fa83c16ef3fdcba530cee1973cf43d6fb25854c2c1cdab92d353b14c3698560b4b9365b0129317bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25f4581fa13ec14b694a8be58c8a150af9b15f963d88f090ed5ab8e661644a28ccec284ed4a7dfcf24948b4301;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c4a15cd1a5ff4647d7d01683fe6845076e9aa4e1002c6d3afdcfb629e776708062e049609624c7692b91d776bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94c9cd58455aba2e06680bdace59161912283aa6da10b169b526338b6e876cd92ce9b8bac37699470482607804;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20191ffc16095f99b85c0705c0b01e2d3f9869a10333723db644b27f76be12c8d014d4a5411c266f478a3b264e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1760b56b14ce9dd0743c3389abf46f41a79f95c3d74928586d92dc63a66ba764db0b4dc9d2997ca177372aa933b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1094bb25a5ab4ef3ec8f719a624572eb8d5c2ff2f85283bd09daf7c60519aa8985795c694325a8e336dc73d2eed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1300ad58d468b8cb753993e87dc4bd7ed4605b5ca99bf6580f2c7d65116340dc567ac3bc948e40c5548c43a22cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191edfc7aaf43de8561623b5c9288da2610211120716357dfb3412008eabaf92463a7ab695338578a09eeb9fb95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he30e4720f903c618e8d95014de5274b9052eef93d0cc19ce3dc954b743ecc4c575034e822eb0d404851c2fa0cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a962724f13ae22e130c545ab59c5846d4f03d8ebf950d1492ac1bb9d337391093395122a3924d432cb4bc1b28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164bffcce8ab9dfaa88479e57d5b6cf5927aaf8c97be6796bca5e870180e24381a5dec55ba809fc9dd77cca4702;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4250ac9d3a69456e8daa5b16c6c0034941249c384203f5f693e54e46bd771f08afcf7d9f813c7d90c97f051670;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2dff9cf68d262d4047fa7c614331d79c9eaa9c2b504707cb33b0cccf1372093501db3d3fb8c262f5f286646ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa4523eb7b0291b76bd5909a7b21efae6fdf214b6c825144df5586a47a57199a74d3ea83e3fb4158fd7b62ffc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13342b7289a288afe5009e684a3637d112c7c88cb489898755f132a739871c0be43c44cc12bfc2fdd2a354808fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff95796d6812814cd7ddcab0bcb60685a785997366c73f7bc30504f2df850967d75b8f1c6498a509308db7d155;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b52713186a54b1b1e91cf8c21d01111b6f3e1409bc59ff37d034e244652a14960b910a90588f64c64328fa383f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a2ed6380b788ace67068d1e5804227b7e4b4976b7e9678994a50d65b4f9e7ee3eb58bc7c2a11682969ba498a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h915c0f1c61dfea3de50342a742b023554012ceeea9b9aa51be26d529a9a7020ec3b74b4fcb0a1eb944cab03df8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184159346c344e5c94ced1fdff011e788604897bbb52d5c904e893731c662ad831f7732f59dd8f75459c9430264;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d39d0271fab2491cc6c7a07fd39aaf1165afd5ae3e9fa30751e1334c4f41e9d538130952087f60b6b043935af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ecd5758306d8be7ca4f232d7fda0ad7741c99885fe53368367620f6ddf936761d6ed165548e78cc2be383a55c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af12ba2dcd93552174afb4c281a8ebdc34aada6bcb15ab177652b7745bbb6c9232db64bff9f1fcce896602392;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aaf46b0f828381d05730e0e3db881041d2e176ce2ff4465939e312936a0f7cdf8347f7c0ee8994563a5256fa21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90348e11e5b417014454bcee3098e26e18ecbf3d7d9b09f7b86c4280e34988e7145ec46a00a1d6f1c44451c9a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb06aac2cce4fed0afb479a693219e87102c1678569697c8ff95cc5f02ddb154bc8bf30a099b0d7670f7866408;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ef76cbb1a725198344f6b9fc79f2b73021d087daa2c08e299ae86dcc96065a5a34e144017812368a5a1284690;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189850e6786d2ba178db8344cbf5d7cbe9f2f3cd6215ba133d597760824769aaeb1dcecdbdfb2b1b797deb76030;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf54f8c102cea386019d863cc9ac314b802d5249eae52a048152be96799a1180042113b0e26903eac460306e19b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d770486b0e08281e9f397ba95859bb36e482c6acaa160eb4e902f44b7085b75561129fa5e3f896124965db6fb6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf25b921526c63b5404b8ca915b7e53ff678e7a2bc02cfa685a228e508b6b5936744a43846f9e5fa9f7221eff86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15428d157fee8b869704b7fc8aa6d51d33e33d39ad2ca611b22dbdec090837d35b79bba1d8471a892d93823c84f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1164b419e4a391422b1a419a63914c0a9fdf2626273690369092eb0d3590b825a299398bc93a9f7eaf501b6eb28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83ab7f8eb82cc96e839c7819c433ed810361418993d62bebd6c696d5ed801bc688d968211fd23654988adf5edb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6d7c1a674d8ab3e4e76ecb66c30267d010c93987b6b2a7d4809533ca2cb89e2511404c2146c662611785c70fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea1e52d925a6318aa689f9da94249011066d39868795a8c89cc26ec4f35cc2921cb92f9e5377fa54b5633579e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1160c4d64bf646025241be2d50399d3eb4096ade30eb0b078641f8de85e7f40fb9a6fce6385a224b8076c81a755;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf948aad1cf94950a89f7cf367f79fbea63b6ee1d06bf635e8623c0f9dedd6b2c419655c2876690e7a39f7d94a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14952ba6109208a0bb9db675ffaf05712aba362a3d2d9a756090d8c2acec9169c30cb173c4f239aec6f6f479368;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h604564e52beef9f2484567009b4e73efbe2d006556c7fd1c396a462a98f2c47f8e62700bdc455c34ed87fe998a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12eea9c68ff1f278864f9d68961499fe9f5a7ffcca3d6344faf894792105966cd441f269274b9345ada17e66e2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5e1af15a71a3bb84425aad558e6a1153c7b0473b6c82a447bc8df95a8b45867e8ff239f191d79d4aefe242fef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5933e28717d47e4bd8012c1caeb9ad3c1ca15cce9b12774b9b3b5a837c9cb6fdeea27bcbe5af8ca2c619bf9c2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf233a0cc0babbaaffaab629b593a87e5cd5152c8da697648ee04bd0b365e07cbd8612b72c9fbf0b297ec4d4f87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c48ee3c41f6cd64b13d112d56c2c8e15856884f68d29f7748750a9abcb22380c51ba098da5ce57205be433d2d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25ebcf7143d3ac9d7640747f5a2c6b1a59372f1f79bcbb4b06159db258d6daa7e7b012ae19439340a4cb45a059;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46a22bf2799ba995a6fc24b803f04f1deca3ad9503435b3f32143655713288a16a1a8e04a4a6dd2d0de2906a8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb0627a82af286fe467014646f915505a7da1e9748239a460d15a47f1eec441695a510833231162150a32d3b2f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f46a06fd8094a8b0cf1d797d942bfd15ae189d56564406f750c335a76c7a54c60ccafccc2c46df7fc66f254d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e3b91737dfd3efb3360337d2ed1482a9c2f8ffd640256f92a5270f449b2cd6a37a982f9cc1f92a83b3eb2e73c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bf27e126061958592d6428d4f790dc9d615b86f9946431699531d08a0400f5e3ba0cb113c8d397fa813d87358;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1648e55392f8a8498969d382b0d2f1571a4580aabc265ab4e57ae1c660265c2df05535c3c2c79bca96ac49203bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbcb38e2063a56bffad3fa160d5682330be546f6b3bbd4d46cc8ebd1de6eefac41d89736e92f7d10a6b3ab01dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7eacf831e56811db2150bb2f91b304ed1fc59144a59b6cdb553e361728a58e4e9c4b5c126d18ba269ab56375c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aead4487eb745ce30b5499935417fba3045dd9d1e288fe756fe4bab3e91c9eb82c7eaafe1462d4e9ab367424c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a66146f2cb4485b05a29620568c87902dbf911fffe639b20d62d339cfdbdc30e881157412adbba6573b1f7e06a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc7c5a9335214fa4f5fdb61a5aabb46608a5b6093bd0823e4e1d100b7266d33c49c8c9c991ee14d3d2ece45bdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h823422ed4d71e491433f90bb13a61d3c74d57af1879b5fde6278fd44ed2f95b21e5c3e12499516138fc30124f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c693ebce5882e965a4447bb135b39274614305b38e0742ac522a243bc8474f56621f063e85cafd9ff7a06e1ef5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6c05544ca5bd893cec83171b88e81dc3574b7af343db2d21f6fa41cd52f5c6316d84dc32d0a2dba27cc66b580;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1983c8b13ccb7e09e42891909aa12ff41cdef57ea3053983c430e9d9c43f108e045fb4a799883a58206774c2a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1895c356f5da73638a2c9c072194a3aa51ebdb31ff5d6efa688785c43c72e2209b06fc03916470d324b9c32ef83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb7a5b0365fbcf7d726af5942d2c486a7dfcccf9f608ed00835f037fa106e344a913779bb840e218577302da4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e27bab642472dcb8377256e7ddbabe5d7cc14e637c7d9f1f6309c8815948644af40bda640edba6fb33c1211e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9c773ffa3be6371dd082f6c3cf856b4fde08ab06154e0445388759011b4372108fa5fa102a00281a69a2b810e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b55cd83771f0722a3986d09cc4f487b52659ab6040fc828caa1e28b3db5db26b0b626ad981893bb58782ed88e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d669d62450a8b7407fd7d3bd34b3eb04ac4a462fbc943f64487382da67c9ffaede59eabbcfacfd9a6f53f34c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he056fa07d67e1e92d82138f7b2d6773c094fca37c42a09330c42f42823ecc58dd90ac1fe18fe973ed6f76bffd4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c62c86fc34bb2878f9c28ad71915fa16ccd96cfe5936ccb2b5c00b9faff16b6de5b7dee9456511b70e86d39e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187ba84c13e5d62a24bb737b1f7d8c30c2bc0304dbbff2017085568369e97411611198819b92813616ce04dfb3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66bba7d9c367f39ab502bf3a4c34b8bb88924a0e5fc3f5a377315184fd5eedcd7027bb8d8ce7596155d92389a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee35cf346a5863e5ef895844e3b506513240492271fee25bcea7f71b4b8c5a9f82c2d6ac126b7aaf1b181ad10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc82c32456772a6579666e385d935a76cb51c475601a5959dab63610cd82f5a01d7bf72fd73c2588caaccf7e3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d3a5d65514300862c86b7d5c6400fa4678cf576c2a8915706acd557ea22e9b7bc17985ff2aaa7097e30ff61c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3575b43f4f7f7031ebaee42be40fcdf94e787a764c1a95189c63da83c620c060bfdda30aaf9f8fcc7ce1a0ad4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b1ad696bb388e00b6959a5afb5b10d05f029534adc80ce0b4b7934d0ed504b7c1745963d044b4c48733453c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a21f36a8844a401b1970029a2f27bf85a10909fb57cc5cecaf9fb0ec0ba273cba6926fa76f719199f7f6f342a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e1dbc1a8ad063afcda31682efa2474e403fc425d08089fb2d27172b2fab1aa97f0caabd4770c799d93be6947c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9f312bf96964783d707d457c915a43b91af2000b70e2fe798333baa4785678592e716295c2da24c56d62f0be4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b010d4f3cb74448868bd35418b899da7ce8c0376d8c84867a09a171c3c86bf4cf552d50354a34c555e361693bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a0cab78a90a6c364147c3079f82fa01b61c4da2fa61b1943ba76017a8e5825363eee56c0f4542dff0ee5192c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2ef90946b395f7de6dcbc113b48368a3613968aa73841adae3e0ac85e0a003ff3271dd527e1690a6cceda7464;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156b66d63ea0ea6c0114923dec2e8e44ea5554d8b6ed3688a4fe34aa52663ef3adb314e59da29062ede4878e343;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a977c7d8fbeb67920c89cb1f14cefe2b45c1dc897e0c2fdf2b6ed96fc05978ea9e73f898a36eb2e8b33dd3d2d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd791e35585e99802d2810a43ca0a97db44c7db2eb6af150ae04b369450b3dffeb216c45543dbafc7827717a79b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13948b3a539d1fb8812b9a9fd4f6abf31b6bb48188c93ccd5bf9c7b207adeac3263e6005e6af7bcf2ee022ec4f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1576b14aaed7985543718d176ed803ab820d0f253e2bf4645aaf1ac17a19ea782864019024c5fa2d13d2e323484;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16bb2e599623ab4645372a3dd0ba033ad5ef620f5b1a23f2eed24ca98cfcf033f61a810405bcb1eb38ab1ab8896;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79d5799435761b87d8193e902afc601d6295d6f2e043bce2401fd2d2df5f3aa3fb43930f07b2abda98944b0956;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h983abb923ebaab3c6beee431b8ca4a170bd890f1b7a8f99bed7e5e62598090dfef9edd7181bdcb65982a575dc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b83c5d39a478b30e6c78bf27c18d61fd12d6edb92e6728c95637417e48b01e0359d8480d23a654a9f4f70d381;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143856ac9d62e09f68a5a56c953dfa4c7f631fd25c80a00fb6a48b3d38738857ebe4616a65ff4acc7a9ec9f54a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b2b117ecf473868152567dc9373176cd6ae9c051901506628cc85a0582f1b144183fdc0a68082b5157914c771;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h207d30c3cc0251fe9a31cc248fc1e2c2bdb374952666d8b0f295a27685059b7b0336d91e19ed25ac6d2038aca2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6bdc5aff817a704060ab728105da106e60ee46ef39cd22a4c43a67ac28d5368c6afe7e2b9b0c04ed5591724c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c7c27d123ad902f64dfba3a66148386fd902da88830c63e4950664c10c2d1fbc46c80e34d793da314116a67da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bbdf540d2e9ef8d890abf851c8230a4db25f7d8978e59b817808a4b0e04d7eb0f4eb8d728e10fbeff1d65f51c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda47994bf62cd6074726a28363c5fe98a9cf45d8aef63019e684e26518ff413b36f4ea47f5b321dd52bd06ca1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee5e4aa39245cb6e2a97d80c0432e2a6ce21b63232547c1e74bbd29625bfd8dc53cf01c308d626f94b482d7340;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a68c27764d49864d717e50a8dd23a8694380575bbbff99e2a8500375e37ad04440b981f7aa95d831030e1e738;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9120757d52f25fd66d1ff3c96acaecc44b0627e8739485d541e8262c5c273f076e431ae7b4ba21935122ea29fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33a036b520a173deac0286e1d0c5916c724f1f11b5d1f3f2dbf177d6667761f21d491a005d071b87e9d6711a5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155e9e6e4f483e2a60ed7b902fd1446a94fed6fa041dfd6511a089a4907ab9c0499854d5da55132dbf5585d0b74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd71cfe43cff1ea7c47bec3a146ca80aeeb45d3b7376845699c8980c217c5104787004e7e02c9a524b873c4fd1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc922c7fe1d8712eff5ed3616cfd997fe6562e7468c2b408ca206ba0c2c9242b9743fe61ecaa79997695246af3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fd1f9b27d7e7f9fae6ddf9099287ecad5717a581439c68f7b296b9f75e57d54bf4ab3ba4bca14af132305be10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d525b760f870745b522821e2271072cabdb162129546f577e5660cc6a9e0b081209d8be1fe45fb19b1b3b94b24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a54b6c781f3dda57aad57776cfdd64c2435e12901e1a9602eb4ea184d5dc75c2ab4c985a62d94c60aad3de3d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6c5b34fb92fe4c097746aca84c85502489970a037f280b5e1e99eb1e0ad02129975aaaba617ad7655db90e4fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca5516a48ec32bbece2117fae630b7d738738e749e23089e1c0a917b7d26b006ffe90c537708c9c220a8b62af8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e874b35fb5b03a9f9140442c74a54212fdf5b7d10f0343558acc7da61fb11c27168532a09fa293b9cdea2aac49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba86f642412e783478986e57a3c1ca916ed7469bc955e795f08fbd6f2b0133dde3ab1e637b153f6f7eddb22cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182903cdf9541b9f883a7e265e3cb6772e8a232245aec360bd081eeaa983772657fd744466f8a43560abde1825b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10059bda09100ee107828ae0d2a2a6ef72e4e918df5eb3417fcfe35550e763cc9a25a57f7862554a0923d3a4fdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a7bec96a6d1e812634f01e9eb0052725ecea2b48979531a46fdd7a25a90ed9ba43849ac541c5905e61990fc38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d94897df68039f8920b2c57bdd12fc94686433a97004d3e086562c6e91275cf38713934f094d855ebdb7b0d1e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7adceb615e077bbc09810e3d2b11262e720f6cc7ed2c1059af7e841dc8b11f1e918a3706697566d4809b0831f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h460d4b1c9cc668ba8d11eb887eb870ba7b41735fe7574d6e66177843751fb7a739aaee9c504f6f3f9993214eb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20de00f2d5468bc99404ce6389b5c8620129d2bfc8f4738dddfcbf6fc1305e864cfc9a5cbfe50f5a869d1637e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0aa3233daf7d5e07a9aaa4659b2e86017a1009ab157c86e4330ee1d93d19e1ad6bd0265c247290425176856d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb48e38919c3813303af2751d2465d656fcb50a210d9979c825c61a2d59eab1662c8aa3f2434c69fb86f15d1abf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155cfffd006c8e297972e9b32f125300670963193fe1f55ac505b990453cd825b6d8b70a5c72cc9a9dd0621236c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h319f4b1d486b2195ed95fb66cdb0718bd7026b145d103d8c8efbdc483010d02d03c036f02e9cc8ca5c08c98c3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b0920267a2bce776ad49039d38e0f33001a14bc48284c1c3fb44ee012bd24aee90b9e8c93cb2ef4e1f2d5ca97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b46227baa88bc6814b99ef924e57bc4d8ea8448d8c8cdf46e1896c35b80dd4b1ed0bbf366cfdc0cb051208c1d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ebd536e1f9d0c16f1ca121782f46111f966073103b9625a5a7ba9cdef5e4bd460c693c26b1a36ebc46656f74d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8960eff2e6df14530d26aa915febbb9ab8bcf0171f1721c3d987bd8337121db591e99290cd37a20f9b2c6db226;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc04165351ecd5de476894643daa05a9579778bc09e748efa414a4fbf564007bae4f2d6f14a7b0354aed4fa4f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccaffd3e0e2e18192d2877d9f246fe68470930580abe7f03972c942f05ada323b487345c2f3392a05f50d8958;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4f946ce750bdd82f5bbaeeb2ccc6a64faa0615582ea79d546c5a976f849b769e87025166c35a4862be6532a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1199296a5d060b19bbc92e09814633e1573f9ec06781fd9ab0e21c2fe57200c890e4433949c5987a55886c4cf26;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68cc7317ab8118931b88762f97dcffbbf5c7aa73e8c0dfccebbf9f39770cea1c49e8b1dc9bf3d2c8976ada6b7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131511e393cc923d6cb481eeb74b26fbe265043192bb2e03cc2ad57573a72b37f2c1cb7e82be8d8c998a9a20ebd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6a829a3501fdb12b7f03d4a03706ec517514c44bb394c07df18bff492a00d3c37dc6dc1d78560593f56f02bed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13539deb18a2510402a01ad22921741d147d895920e884f03ef8d24fced2048e6f22645b90af29d63bbe0b1e4a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac713bf75e5148c558e132be802b46727df2721ec4d5bca7925b61e39210e2a32d0d2fc10a72dd15f363265424;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4b3a0c0a9e45c542f106d99fffec87a020b6b7490d3af9a964ef640ec96df89ecc106029968a4d36df1e59ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c86cc9a021e19e0bc932fff11ca7ba4d3bad802e9083eb4f9ac16093cdce0f7dae9e72a56c51cb19ed45bda22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1570ed922559176ca3474ce419a34b4b7cdc13979bef9c8e48900a297c4a67445093040670dad2afb411af782e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18aa25d8be5fbe6f388760d9885669a180246f8ea734f34a374c8f9358f171ad36c095e47682fc1e283a0afca0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf0a32d35f648889faebe76dcf2ac3b01e5426ecf4e35067ff2283a262df2ff849ead0e2fcaf5f46282d0a4389;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122281d3f61684ec8faf928e42667001f6e229f0442cf18a5d226e0868f6b6353ca6d68b34c7fa171ddd56ecc5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h96a047b522522d941b70f0982d7794c5bae5914942f8dc82ac1025ab158e1847082bdb8f8adc63c445f7c274eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1206f4d3bb48b20460dc6aea25e2a8d80d53f0e4cf9643a2ae1566786c1b9dcd022f5ce2c53ced55367cfbcbb6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a639dd2397629a62588bcf3a3b3d89e29d27494b0f41f0351f3c374e688b03ae939bc79555703f14c012dff78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ece67fe12df1642a729403a464eaa0dd7bb5d15ee7992c7e399cf3e63d2a8d47be2da1b41c657ec44eb142ee0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffb1e979efc64a72dfb21489809e8fcba8f8bde1f0b0e0a4bb7d77fb0ea79a9a35fb1f7a42809983be9626491a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f4962acd66938d90a2b3623a927bd3b5e42731906f3a4d70f6f9f3993d5ff935ca6a2fc0c9f2b10a8a8a6b70e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb74400af02c5c7bd550e26f2bc07b2b3f8cda1425a5285579b6bb9e202ed94cbe7c5e14d715d8be03d370a670;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1785d01d972dbd4662bddec8f71fcf5904be0a86580c72031d163001c8a8dda828ad644ed54a097c04e1bfa400e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e76ebf026fa27b2f1314b97eda0a8ed92cbe31797e39771de06fcd0084a48589f5b33ecb2126f961e1dce233f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141aeaa72118290b92a384d9986ba3e226e58583b04b1ae7a49d301f45ed37a236f4352f0476ffc2a14424a7e2e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c45aa0512704ec98f290bfced661248f8059e21572789361b7b42c4237693fa4b02c3c08980dad81f1abafcae6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a395121976e3d1079b15dce12c59eb7f3080ca3b46e85d057e577c7a2311b26f9c8a06ca5fc7ae895a6a716a53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14989ab23aedb2dafb2591b3acb1653b6f53ffa2b0d06d9862fed47e18de4aafb8c824988c75f421176adba399e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0a356146be236b722b82a6df4f981067f6fcb3ba2aabd6c532ff156cbf283dde30f1cbfb4564d430de6f7f76a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h453d6999e19e3d74702cecfbd9ee7beb913efda3a25634600a2634ed8e8615e7dba9a7d726d694c2723131830e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf98a250497c0be9f61fa0c737df7708146710ca39f68784a7b559b0f2f89e3c5f8f46f68a63c2112c91a8e735;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1670aefbb7526da870039bdcec3c5ecc76baecb16194d46205dda8ee425d9c4c7754e06591731e48eaccc9faa6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc716b502916e6fa6482b150a8b3e1359ab89e005aa68f6899bd3e71f2af7360ba3ee4aeff8ae0a2a78604460a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29959d5bef6674cf118d8b313307d489abab3f4d5027e81ea047650bd82636f1ae497a7c803f8006c53455e6c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148b6b4eed32a21f5db908724626f16c2c9c25b406956e1cb23124d47956ebbfaf36671aa1bd2444cd06d38c0ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17dc9dc3f517b2417d879fb61c25433552e7783d92fbf423d181bd6b9fcf4cf08b5c700c6e4520531e6bab14b4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf70aa64bd054d2150546d6b879032c6de3420c1bd2445b802a0f79bfeb429ab9db8001ef6a473ed8c6372f255;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5d11698ceeaa89747c9307f31f7d1c331d18a87cf86bf86ad6ff44e2745776e53ea3372095b73cb73d93609bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b91718480aaa734aa9180bddfe4b0d68dd93d42070d0ef36e6bb703f060422f121364888636febeac985ed0653;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14454294debc520c69c738223857a0418bb10c3ffc7c9f09c0319335e4375386deab2e28bd36be2b93f4ba03563;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb41435881c192faac2ffc23efff3378d45084d024cc7964a42cffdad56a4cf692075255f4e7180c5532adc56ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2de73cc42af21759806c6e7f2e4e84980320cc7b4defd0cf62b002ffa71910a3f4526ee0f7a1e984065827c50d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f77e02b3524547916f9b63d7f6328d32767fc6d170bf18994020119a3c0a73bee90bdefce7ad232a7a915a0088;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14080297268454fb98ab8dc4d28483530c9f86c53b0709263c2ededff06465bf30638b03c50843949de5076f280;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9761ecba45992b80db7f257552137b7a1c948ea5ae8e06bccea075e81d97a35fdfe0921de271017cb7210b736;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c7079d2862e4bd099c5e3423cb8fd247493e7a1487a2fa7942705c4d85771a47c7fdb790d7cbe7d428b9c55bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcb14e7ee2e8e330efdb1cd4c8ad1112a81d470bfa25e9e36e5a9d586bba7834aea733f19126c16ed2369eb63d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199c8ba35ef8db90b51f967690245f4c06ff70bf1681aabf6010b2d2be369909ceaa65ea7f701e98c684231a731;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ea674f94405e1b0053233890c50cd10e8f3a3901c06320b25b742be1ceb4925c04aa9ac261bdf7c915e3cc8c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6fdbca69bb2eb1b26278f1af7c40f4b2749c4c75633a1d2d7cceafd6b67bd889da4c7b592f254d7df1ac9c676;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8383f95edbe72b7b20f841e244fe2577595d5f21aa938ffa9098ecfd9d0624c1ec9499f42afc9e6d14483398fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19654bd0230b4f91fb6174dfcadce63ddba539410adf5753dbdc6592f4eb2df1a976473d234a6fc30bab738f589;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12121f18a9a3a8176c97921d388b5ba123a402d618956226ee4b653a27cfa2f60781230e85cf304617e27ed9c50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cd66d94eb9e5a4ae56cb780103a6dcdbea55b051886a78acb4cf7d9d64887912715c6e1c9fb93984673a9683b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d42c415e49664114177865da7f8ad4758527e95bda3d30a7cfdb898f32f0b7cff64a9399423d59e4fdac89287;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2995d0b08f10566830dad41875be02cc53132a3803e0449930dffcb97cae27d239e1f7766ebb3547ed4c4489f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8efb45fb9d455eba76e9359abd6aa749752ca45174748cfad3069e2ca4817de3528d0f493f7d60626108bf093;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22e1a7ba20b5e9a52688a785bcfa90c905d7997e38a69183f888458ee441a40276269cac5ec9b62e0393aef8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf6359edaa68d526712fd0c0f9bf6b57ef6cc48ea0b701a690b1aeb017e1a2293bf86efba5c067fc73452938ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf47ddb85c61032f157d0ac86d05390a19beda3f21b7205d581988ab1a1722eb93c258ebea28af99f71a0fbb56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd257ba861f5127dbd6d4db48177cf74730a25816d65c8cb716f385a49369d6f12d7f986c3ebcc3a2af9edb327;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h243a221080be48cc0dc68b92682173a36e88f412f43f93de5d9832e2d6e809382df405a7e9b8b1e98998abaeff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df67d7231fabcca420338f99a5dbb5e1c4554e5da376668de0202f1a9fff3731c30e51d374dc4bc54ee5e6cb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2236de005c751ee7c1bcdebc79110548446a3652c234cb445e9f8a47cfaa990b2945a5606e8c1d918334962764;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b72c7c8e7627d4bb805c6327c088db463d7d7aba4fa313fc407753668e08ef350f853ccc772b169545ce7efb84;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he20966de5caee21a4a08b4a3a0fa5c3a31ef4990713822c2b1383c86cc6bb85c22d1ca49fecdf183141f595ee5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d29dbcf1243586977c89ce5a1b63c4a06e96cec6e3bec5cebb43a3548db3e01370280a0772eb41758160cb867;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd04824c85f482294f2e3e8c7bc1131de5ab55a1b5ac5b3619b7a8525044b9c37e34cef49e9fa4e8dac63bb15f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81418f11c07189eae2b9a4015c3652f6d7f3de046d3413b9b68507133e69c7cccbbdfd20946a72cd964c9e4da5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121cb9722af86faca1f8a0d334edc73d991cb1e070ece2a33d76975c9fdd016e7e1ebca1cd8fdf75c174ea044ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h486c3564b5ff4db876b66390d6422edaf26d332420c428b5e292ce64b96780534a559da9e420c6ac10422b6252;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1404c9cdd7d9bd1e090b6e85eebb0a3f42784168342bf7a25f930e841da73746589f78ca20e3d24d8060163670f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb00b25788cf1a57b93d18f3b76c3cf2bb673d86623358921b32d4e31196c53e139c8a01f4647e842c164e34385;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2acc9d8041bf073c45c4a35cc951390122e608a65303327883cd02bba9536c871c4dd071b4a0a26d4a0b989d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110557406c77436b5cb804c736deab2621068c7a2969b98f5069b374a22313f06d66b2d077800b2f181a54e5aea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e355c4bebaffa1a836945e51aeb1398b9ac823d1fec6106e1036cb3a273da0cac84068c722ba0b9404ce9e56f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c75914792e5136fcf44bb87d3b1b9781c8dbb647833cf737fcab3f9b6d6259a18bdf6082cca5d44d37999df35b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bfb72ba6d2c204dce283ec3410262b4f04564ac2f3bfac91f6ec87929dcd392f0b6880fc3e3739ae27f8d36bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1148cd8c217b1ef6b2a9faa0d8a5ff7523b8ab733a371c1c3b4b5addb696439a2775a6054635e75f0c2811fe650;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea2cc5aaf76d91168b7a7103c9894ab574e266ab7332fa501dab9b9bc134a8d721b152ce171a6843f16916970b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12467f6827bbc773ed19edaab472560db3a7320205030c3c4d0a3059495303d56686751b25af3d6671488120948;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a8269216b2fafcefb6910f29d2c2264e95c634759c26a97817c651314593a3bfd42b19e9dc462b704b0358b92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd02e6ce3cc760cd3bdbe8bc764d33c950d011fcc4787c495f83a9b3f13f1c1136575130786e716dc360c17058;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafc4072c4befd6d729b0c6fbb22ca7fc08e876481808e6d505d1ece5714f2739c98d2ee7ab45a5c2ad2b11245f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f322e9892bc0a271540bff40c53035c7a818eace2229c84a89a5207bcaa92b241014e029f778ccd6a2ebf4503;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb2e6ec15694081698e69adc7808898ed48955f8fb3b77000388d40a3db410d0d29b55c417abbf2b8ec0b4bd33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75f7b7deeb49f7c8f91e641d9cb42f292b5eeb2490adb483fc49042816461bbf02f2f6487e958c0b08c2f3bf89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5fa58b95b62dec362b1300f67342f8b07145ad215c8be15e9d856f7daeeda24996354a07f5d5fba79fd64f7c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53af8b302f188fa72b087cf1a32358ad3922a8481b92738ce6405c4a0891db8f2eef5395d65dba58a92012342;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175ffa43d9fe2a24f597bed9ea71599bc255d4553f101d426b76365c60547517629d5279964834c42329bd97bb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be7f2454d24fa65920be7c4f93af310220b1e78a0a1efa2313f90186079d49834c2914419ec403a7d164e5a8ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e047e15a7f343a59f42805d2d7fc01510f1aa66bb4cc3b4cc8c80974155e9e0f19b90fee00ad5d1df29bd2929;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b925736b3d4ef0b299ad0d7d9d3ee2a13db9bc76d4c6b6f035e3f3ab28c55312a2f013462735a43111d18ee00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1e6415aa0466421cfe53fc24ebe15a48e02012f47eef5c545b116ac082bf3d5d3829ffba3f669038144a50013;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33550f3b8a593bd8d8cfee80fcd91c6ee3561ebbda84f340c64d7d6b5e24cc2df5fa851974c535fe650a7eab0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c5365749478cff0010110d484391eb49f0ccfb1bf5edefc7c5c698d44238caf59601f8abd34f371bdad80fc22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he74d467b564f433cfef4d6ad0dd05b9c25c193f4e8cd14e2d179e88512091dcc4bac8cf288b55fafbc6273b401;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19217402e215aeecf2e17875e2297decb1b303abb575885169ee614d39c2fc40f92d8d13db55293041c44df881d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb20562c309c4e4a6ce19abc3ec946627b7dbd959217c3fbe05193ce72844f2d6e85f09fd554b715096de722d11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14379374baaa8ade39c4b117bffe40cf2ce90a23ec31621afeeed8099976e2bc3600d6d55e302885ff9bb95e163;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0f85428a5c8a42f4379ece3d44403e5dd7b4a6e15c7d7fb9888a50585e48c1aa49a60eaaaf0b4464b8d63c09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ff0fec5164bde036acf59c1bfee8c957ba9d653360fe1001bcae4df8f47d7ae5753ae3ef9a00702d08e0b0c2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1374d3673c1fc747b70feb65c40f37cf31e4a9d2966ef20c21ae4cf4d24c2ff27026009cb07e8fc0e807b306d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1428c0bc4ee7d81332559fe8b7cdf4b7b302ff0ff689b03683032247e5125c6ec24da7f8537ef9d2a209b4cef20;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1694028362392176d50db43ab7f5d831cf6f04727aeb55415ee3aa988a9fc7462e31a60a2f6ecc61fdfdacc585;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173cd46bf4178ffccc42e642bea976c2420338146f4159c887261f111fa8d26d733ed91abf47db575e257ca70fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184e0ec426883887e8c1cbd473832a4c1cc11d4b9483ef29efb48313ab57ca2be2326ab74f2c3072a61aea7471b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1677ff4f8847e71482952a6d00d278500cc52eec5bb13505ad69314325f3b42c384813d17b3e2a141f47d6bb10f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bdb616c376d0708d4ecc37af037104b352f943cb2205cc994a194220c9dc52084702a667a00d0b456da247bc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117970299de05771207465d6a303612c93f65b266673bf711198a5aefa7ca364c405d715c68ede6b00fcc226e59;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7daa17fb9d5ca775e500424570871ffedc3eb16ff0504eb4b99d4425142da705d358232b91db01d181fd94523;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6cb81848d113123b4316ea70af7b8116f28e59317839d125e299c88fcdd67151d9cd889b16abaebf09a40f16d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41043afd8e5e3e08ec9a4a8a011e63f7af450ac83b1d38cccbb08004073bdca91f616c76dcfa20464454d2e12d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3505dab62abcb84ea3f2d97c81c0eba5fc2d6ec5e445c97388c66cfd3a0dcf477d24e6dbf877c9ba28f980db39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140cd709330e7a510d82f74db140e4777171712e1d63b8b5b26d20815bcb6d73b172b9461983f4bc2f05b7c130e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a914a8fde4522775ee4a3a855995fab1ec0f3a276a18f465ed50870ac4a36d42e78815245a90c960946e88e880;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb177580993d7ab82fa35bb96ce664be033715a61cbbb270656d1bd764c41260ea6a68c4d928961dd014f646f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8271567b02b6730e6bf89094f858960995cd12663a5e1298ef96963104757d407c82ece06b2eae1bf2eaa9188;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107a616bb839aa04de9e283a9315c4b6a47d1a561bc003781360c2450af8ce26853eeaed51490062821b67ae9d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75cff8388aaab49f95c1de069e41e49482fa9855ae803c03d3e51f7f5d5cac6e40736e81c2282ea10c7a4a174b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140b3bbdf054a244bda479dd3acaf0a02bc41a6f74d6d07ede4ba19ebcf07dfe5d4de475fd2c65667a89f9377cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146265dff4d38e25a48d1a5c6e86af271aa552c2017ce7649dcdc426c6cab5ce1d99f1a15a8a1595615a8702f64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he657ec3c6385328a736ec9ab6f76d33085b9b96b103efc3f2db44d169d4c58d9c1504c2005a814bb1e68136a3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a092875f9c2fffc570964264fd303062d17e7c25e600f4eae73a029ec398c93c3dc3287439cec21dd058a2008;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba6e16044b1822ddd479584bd46be67a58e6080d85cbf12952c3ea91763d5538cd41253ed1ba218d5490f1f973;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b808c6f1f7a0e2f4950b489705d13cae189592815972c4bd625c692ffdec0b2dff211febc8b896f3bfc452b37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c575a2b4651e499065f7a723f77f9cd48bc7a7b0900ed07b6b0daa4f6d3cc3e0d27ae9a2c47e3425f56adc115;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1020191654a48bea7d3c672431769e6a2360badb24ac0dd5910491eb94c572fc7bda0c5df5fc2112da207139979;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100fe56300bbbfd6783b080b9ec43b00afc1aa10b274ed80dfdeecd3ba58a0354900cc31ce6ef2d9fd32118c28f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195c7c55d3553e83b3b1ebff6b5cd74a90fcf71518ff749ab0900f95dc9657144a510354efde328825fa0856ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he62d6fdafa1a2891f541ccaff7d0cca6c150a3865dd88b5fb28db4239a4bcd1b6890d2a2ccf435b70782f81d7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fa01d94869029c06d8e5292b0f25e048b69bfc441963506cad4e88d71b40483414004b1e0e82ab374eefcc367;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab972b8f9593efb5f358c2c588640db892b53b2372ae1b40c44026281c9ff659e0e562f5afce82f5a2b43d96e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce82a6904ba7759e0a96d3f5e4ade57f30141e59503076ab58c011e8f4b171f31e97ab13f10aa55ff7f2b79f06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78425a1b6f3fd20da047c8f1ff7201cbf61b05e133e863f19013bb657d02bf719daccd124e22d84e48cc323e01;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b26c6f9b21e2c0cd64cff7388bbc5ed5d4a5a0e1e86769878350c9c11d9f4465c8455c1a4aa37f2a1800fae96b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5e7f02d7f2b0f97f3861888933a046a135ffd5e0b207d6eba59efa11e67644298c9245b12d097fdf07abdb759;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f91676d344f150afb52431b8a883bd184e1b72870f8bd459f3c52b21aae88467281090d1e56c064c29557a1f57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33e3367e5b66cb642a701d04ef2e795e0dfadd472c6a2998bd5198e55233b8db4dbba3521eb536bbca2a14972b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e61f029bd1070003b7b37afc9c592462809b97886eeec457bda8069804de7997e2728bc2bd3c2fef771d4f566;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c79ea34a0875f49f00ec3a9c325634088b8f8b47cd9fe8c797aeae6002c02f4dec526de1d6f402c6ed91990873;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d00058c253a76f08f6712cb3fd348b1b8aede1164b224828b6e3f6e6ba02c68f95b682a1f236cdf48bcf93be5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a806577982791b87456c4376321564505766c876d3a0e1f8c304e4fc879efee8c161c1e1d2c1f7aa8cb7d6eb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd0195568df9298c7c11eb3a873b12d9e1add5a30b1431cfff31e2a35babf82fb9ffbca7e552de797d3640e9c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1898856db4dfc07095d81fde87d23d516d65779d14a3baf99ce0f364e9ba3647440f521e075d245cb8acde431ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15566cc6a030fe95bf47ab009edd9324fc47c96fc95e95b45de038415f035fa443e08d08dd9b71ab0d22341ae25;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had2ae9b755379a5e6a305331e6f20e2a5e9038597830a18ff3db8c1ca73021f76b064e11c00dd52cad3c6b8529;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae0562a8112a2979d6db3e9d71aecf8270bbdd39c778fb60d21fd6403ac8e10bd613f7295f9d6c3858a2e78695;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9117ec6d60b88e8561afe727e486596612ed6dc614e4601fe9e0c266646929cb9964a04e38cd8ca08793fa8576;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a60fb281e8ff585339c340f807ff9b07c9dc9e60a74d23f3b2564e7b0b9348fd942c7c2630aab460622c3e688;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f8e4681db09a3ea3e94f9298253a10dd414db3abdd705cf9fa8972964ffe9852fadf6e0fdba20d80eff7a6994;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcda10c3453868aea272f6b6024c961894f5b3a6147690401c2ee7f2cc47c7c112baf0a5ee9e57ddbdfc5b06379;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6a38617a2e0d1f4697ec7c81052ab17e9a0efba5c70b6585d388eb1f62a67567f8b14ec4f2f0624d0bc2357a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23eb949467f6a94ba3bbc07621d75f91abd7530a19d772d6e1f53903b85368b2dfc094e0ed258ce80c7042802a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6c69d0f1d1d558ff225b4a3d4fce6c4b404a5c00fe2400b309be95168ccf11368c7908c1fc654c90689cead3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdaf921fe357d6e3707934230cba620d6ea6b7ad18b245606ce58b8df570823b9854ed4746bfac340609fec9098;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdbbfbe5daab6b5bcb54845013f73b956e47294cf626d3482794fa722c5a188dd833171044d3df72d7e586a128;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14613b978891e123b7d6558da7b0985cee7707030da8d68c484a4bbd8ff37659e112cb63ba25d88bc6c89d36855;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c3efcca746e1b41517b7a025fc10d6c5939d91c186eb1a017e595f462c6cb010acba5a532a905f1bff06f58ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had9f8b3ad2110b5a5753ff86deb5ee5270206969b9ef178578fba08f333262cddac0bd78cc61489488f3fde69f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he74dbfe66345f28bf38ff03b431c746e0571272659be9edb58d522c8af25e516d8212db656afcc154e86844908;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6bf330ad6d1d856325527f3428b988d907f53871a3f90a788301bffa1375f20d48d41ef9a28ff52186bedb1c3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1056cf19016bf482a1607e7c596b05f9fd2439cc6510ce030f1fa190b20e572ad50b1da270ec62cf127c1b49707;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155630b8a155fcd6e771c281f4cc0cc21986969db2f2dae5789c70df36b70f08c0b8de1df688c08b4718775351;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h231999a9526815ee09f9288fe0752e94e0c19b1aa2a0d1e7698b9cc88f65ea78efa29bd172a055989f079df8a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37a9cda528390697705f81fa3d16eb401f251345fad48cf509826a3fe05f7af00676292c72495fe55d95ca6fa8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b8839e37f08840512bfc22ca28f2fbdf930fa862ffc75fede1e15e28223e0252eb50ca47d590ca3b3ae7c16d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1657b25235a731a0460d83f489b73b8eda868ec89dbc531947daf2d53ca000b628a219cb028292995301a850a02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109cfe141040696e8043934302e24b5da3959a30cfe7bf8d56e361048c9e2bf2f612bf20f89778806b6851d798e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1700b7fb83fd4d53194194c8cdaea7879ab6b17b21072c7bc81e3bf9a3793c3002d72c73ea55f3389c7a7b86067;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd8a43388721a2444274f5946aec94ed49733b8b2c0b986a715ce29685afaff6f0ae4d09a0ed4ce6cf1657e4346;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3bf20578c17654962a7046045df88d2296c222688dd6234b538406df6571f1f574a484206d568f15de541a7b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a964f9822c04742f87c69422c2b73ef837ffd21891faab5d2540d62193a47600d31e6832f197ac644442a22094;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7294d6a7ef89bdc5213145523d7dfb30e45afa63f4875c6b9e2fb65168b5cfa5f25bf2070a8fde074f2114500b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a9228d86ea15956a01f0f725c8dc1f6f2674ed857b36e72b4c0cda3260fefbbef21e6df9f2fbf110f492c5f49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8c40b20117b5ff7d4c403674916b7bc3732d721910da4c64e2f946689431d4c7c0659218fdfe031b80828eefe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d4fbee43843f4c3c2e1f8a8bee14e816f4f752982fb86c456c6f9611b03d2337859b4b9d1e54aa8a010eab4fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb61f41521c92cc64bbf651966dea21d03387d2cff7780084c9df967a69b55eee94ba0d7c42ea8dc0d921b83db4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90081d9ea9496727cbf7954ba9bd85040e380efc10113f656439e4baeb896d5d22820cb91cf8364dbeb908f80a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19129b87cc60b2db02e17f875c3927ab40a7414d99bd5839a587ce727d1a8516038d9b7aab3bdb842a19ddaa246;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0a0cde1d220044c3417dcff6f6fd2d0ba5e60fbfcad937650a3c0f162707f225dd7f4d613db2f8027a24b988e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he81e37c08c92be1041dfa2f38840ec51e9f6df874f68cea2df280bc413803fcf9007b8f9e09809f8c38c8b2202;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d123d41c466c98356ef6840627ae531be15ff4c43777e65e645c5e6c1efd80dfa5083b47e92e4c412cdd366dac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad0260c4842a38a337779dc467400005efccbbb9d0403ee171572d3c17ba409d08d36de710818f79ca1723336;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13631813eaf0fd3ebe0c512ff46bb4db8d4fef7f6302a3b6697f2a2fc55194f18be9987fa40c5b675a923bb7c86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4dfb535bbe1f62e7de9cfe7e4a9fb7567d68ec290bd9a6216e6d15e6a50e6d5f13c88ce4c78f07e585a7271f9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147904abd085a07f69a035960764f31c9136cfd622dd0802539bd86305782a980d8db02621d07895b529d5146bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5ebf1ff7cd24eea1c61c17b7e4a45feac78af46362395a34938985043c1e3f2cc82b28c61f6dcad1a09bc27d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39f81679060d135b54cfa36ff10641a3982702204dab04573f161a149fc5108f731418eb9b8c7f61c76686357a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72b3e869fb0d30a2696c830f16acea99bdc5b74e6464b9280916f8d5c7d5f8a8525e0efff0330fc5782ac9ba3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he26165a67c9b0c9d4a96d1b468da32f52b00d7c8e708593ecf92bea62e8b156006208be41f7718d40791c85d19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd415cf2106dcb72cde82e62b22143ca4c3e3fe21a90492e31e07d529f9d3c2d3b9ccb297e4dd861f61682916c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ec5109c28daa1772922f7fb0645bb58bb44103bc7c9c9ea88eb4d2e2518dfc90de6b57ff2ed131c44779c1690;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17da850d5d4240e8475687a564b1401729d54aa1c11fdfdf4b30a4bc5d77255101733d032b4ade265ecf27505c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77cb008f8c4ce484fb021c33c21a2ceb026700a0ab6422a6478ca304e0ec0cc53f43983e07e843be9ff818f444;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8390a1285339bdcfb61e20da75edbcd5c3fe2201acc1eebf31fa7ec076f865e6bd74d575188411f7577cbb6ebc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d642ab5df78b786c0b44480fbc1f8f002540470e6fbba3e337f6fc1e03b5540620726303e5a21332b878e6cd7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0819dd42e948165e95ab5a408dd275bf03c847839752acaa817207e58194e39be56c33b6395da0c83c1194a90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2268ebc2fc081fcf8bb539050acaaac2054a95bd8c9ecc284531aea8fd427f6ee8bcc18a58ef4ee3af33eae7b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f6626aa65f1f76db01b3fc130eb56b4768753c7e3c8413fe2474d091421884fd106fed256194a47d6b203a502;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h855b04dca638a93cc47fbce5d89a12ccabeaddbebb153093add9378b9e7de5f72b597d6c68d714ae2301247ccd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a4c98788da0a0a08af18cd0195f94d832b55bf6cf84e85aac1b592b6c62d5a658f100b76bfb87c2ecafed6acd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8a623ff4e45ea67ccc6c33dcd56ae390dec4d08552a31d83abdddd310939269445663e91436174a40574a6e49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f5817f0427f81794a79057cce9d3a9db719fdc722579c2e04b8bf190d82cb40bcf7ec27afd7aea22ab6ec9dc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1815529dc5ff5c2f7166b221b235cd9df9526148a6378fab29c7d1eded8ff20b01c6e566f27c1d9a3b4062165b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8e120c2fcdbe136e82d6774fa851fd48c852a8cbe2e5b513eba8822397d2e32693c2548f4ec96a490905b0a7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac108268fc0bafc935c0391cd0a20498df4e308aeecff72c6015360e99333e41541f75014f80eff389a9f23b46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac22522f3cd5e6d0ad40b2e2966c7aa80af8b44a9904a06b0cefbb0c2f6afd3049112c03892e3f025c3acc20f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3ed729444025be0ba8672b6727106c8700d7f34bbfeadedced367c3bf6a13adc4c05cb3ebdea52ac7d50b1987;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13443757a442fcfa7d0bcd4e4607deb11584f7a617b82b7da80bc67b9fbddb9d275818e51335feadcc88e32a862;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1767b29952306dece575aafe7b43e3167e052c7b90e580a03f5d12ff95a6f0e33d55707c716de4b743b0bf36eb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5c6afb1de84b9fccd061b08e7fa6eb33f4bfffa0fb52b2d59b4165372af07744198ac66fddc8f442a7d9c611;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6bb734ab7fa2196f4d2ba89e8c7f3c7779b74c6c62b068e95d7d06f69c7ee2894587842d99b6b34050aa501d9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18226b6acb56ebea9bea348939e8b95faa5f1578625ba243c6458505e97e23b60432f3808dfde8cf51863932466;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1977e34c50387a3e5525df510a755624fe1e4e198ca0f2051b64bffb20a0c146cd57efa6d60020dd5de4dc973fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3fa5fa072f2dd638ed1854140fffe32658c7e1eabaee4cd6bed4df0c466fef1516d1af3554dd5e00a3c27f9b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0057c729d8bcc9ba4b07f78590199656e7232eac638082f84dfcb98f9001ac1562aaa1d96e564c0adc0a02727;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b6ea2a8550276b2382150c4719a04341a83281be15d0452a3ca9bddffc3a8223f65c1818aef9e28c04516b378;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1373d271853a0d05040e31556520a49587fd78dce3feef21f06408af65cb9c734984d52f22cd768e0482f6e0031;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b228054e50a6c666c6f8dbc40857a5c0c4a9b50b9f2b8564c6c9615918f18de2b3497a09dda4e7db9012ca6f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc762f7399571449af64c320101c0183153376e226b36ce4cbc2ca7eefe52c891afc850ed0137f68d383a75cc94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1474002853c11fed54a72f7029fd64106bf17154ae59516a3f300bbcf5ac45ade2ab427bcdabbb197cc3b6d763c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb375d95003d0420bbfd82f9de47e62bb5edcbe7dacdef4febc5e5927473642bd3c4eb7830c41437bcf55e5592d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8824000b449084e0f2b71ad97be90db968ec96fe73ab99ff73255cc66c1dd6e51117339bcd4047adfa8b29450;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0443625d4b67626bc2881afe1476c12f07e08adbe19277437890ebc82d74569aa03c45e66721d0869bc8ad1f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1781c7dd088f52040b208168c06f069f3b373aaaa69629cca4fdfe43fd6007abbf904bc2c6268435d96130d7b33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33a952452174f0b4a76a1caf985dfd1dfa54d43f4d3b66d7b36dd3d7ac690a1d58fc44ffa6dba7e25881796163;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h855e99081844dbbde6050e03c2550b097543b66d2365765dfab3ceaf296825ac982cac5f488946390286d47b28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec62425ee82d09b877583cc57c3bc2a3e15ea3ebbef88f19aa7340af1a33c8d8abc8973b4def877d8e41e4650a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7f24eb7efa88b3da44b48ac93df8867fca244501ad0db2ce6a65d0b0396c4316f9e7d66b4839e8d61917060cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3b526fa051b9daf1df6b175b408cf1baf36133f4705df9db38171658e035b93c139a89c9eb3e765bca44a23fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53f720eacbc178d577d34867accd082759456852fe7485fe2e9d70635f87143e00822356121045b9e52323bc11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heaa61a4d9cb9dbce45aa04f438185e75e76741878d45e57ec8795c19bb46c0e3fed263c868e761056d38d0c2cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffe29a1c7a05787f0dbf7a5711c019b4cb34be770ca0f954d5a7774add23f6fa702411b754748e5ecc1a02ed74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc9ff8a4c79af9a53e84b7bd4d0d81454847534c380b7a42af37f5b896eb27262615e5a8e1407d5932be8c6626;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ceae12c8174917085414d7b383f7c91e92fcc1d1f508f8d1a3a3c5bb62112869bb869966c3a1b6408488e3bcfe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f23c195a9034b23a13c414aaddc7a225867e08ea69edb00647a14fc83fa997376e36e006e22354e30a442265e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de9f79e8b52520d36420d6de4fd7249df5e84a5dcda43a3ab551681f23294b5b31e9a68887f809e0d5a7ac5559;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1345723d81787ce77aec43a3047466fc7ad8f5f00efe56e62e2edac421bc5b61c4dc0f5b930a873118820fff6d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12061e0d6c167b475f6d8e00fcc1e77116d4c92540e2039e30e7d3a0caa5dffab4d6bfcaaa1b4824a5e6a1c4b6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10958436b3fe0085c68dda59c5310048614a304fd358e569c4842a2bd5434bb4554e1bbf34d61ddea3c5c20093b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha27691034f2a5d5f631b0299aa76d4fcb1ae7a159ebbad300f666f3b298595e5d5a46976e306ac343d930160d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f28dd65c148ca2842dd010b5e059a7a84b4bff2a0a1dfb5a70823ce8eb1b6fd08ffe368226d2636ca8f95a77a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34a75da25949fea45aab04a6e83bdb6853f175f4bcf42fff628e169da22ab66d4bcad99e0bdaa85876957eece5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ca57c2a8147797c4dbf0c39cf48fd12f2fcf932fe176dffae02d8f0da3efbbf5a4d7f8fed7270a5736fb36de6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5c063654aff45439b4250493d187cbecc97af6ad5cc7b7bc1a46b9c394f7e809668440482bed8f60183fc1943;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hacbd312a481be5746f7baf56d9cf83e1ff793144d5c9446d3440de6fb04406326c41f98a5f9b7c6aae0a7b53b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e773d4f0e7b57fde8994794fda9cc59ed1b0b149cb919a9a5c10c7b7df4cc68a98b3af4004bc768788307af410;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h673349dd519dbe12ceabe8267e7f8aaecdd757a1b1acde636148ce8647613c2bd7490be70d29fa1dd26131f4da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc5e459604541fc13fce4decc213382f9927aeee298909deb98631a254119c846d022079f093be5ac4181f9409;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5bc15b009ecef3ba25e2766ce8ca1005cf461b8e7d70c3adc2624b505e5693ace4eb7f02961382c4309900a96;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1384f58676172a890f8678f5d2863e7271a6a76af2aedabede5d4445da557ad1804e4454ff98ff48d7b77e13f6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15fb825482e645ed1af6797485694ff0b9b015dd4a0402e72afae29d207680355c0c017f0de153bb5b2f4f6d241;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d2449af2dd9e52621ea9f3944b841e8040d3481aabc40e1d88a62edf571f067af132db12d92babb471cf2c2a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h874d7f9c2906e5c122329c96bbd2d584f78542981cb143ca2b4f7420fd4e561dc8f6f7fd5e595ee4c2b8b7d73a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3b77e419f9a8622600a6675d12e9c8232de470db72eeaf7a6ca25bfd37eea1a21111d745c553d4381d0229ed3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf19a9324e5fabf5a2250ce97977c71759952d7faa409e4499970b86ac62e9d5654010542c8e5d8e948b4a09ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb94d654b05daabcec5d64673ff2d4cfc671cf974bd9d803cbc8d7b3003c56c8095c0f6436b84c81a57d7cf581;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef73c5708ada1a31f065421d9488ca476f931d30f266ecc33077cfcdc043796e6efe6f8b7be5c061616c4a9289;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7791045e7c5b0f587bc6a09d2fe581d13a02667f97d94d4820e76989f4f0e3b28f729c0a0d6182f2c804c8022a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haec530b2db78f0500cc98017ccce04d503d75f00faec3ba656d8974a469a36b5dc707568881ceb4aa7c3bdc15b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f2bd97d97fe374af4acc94a38b5c29c079061e0ed7850b52991e3f8e3f8d4abdcb7a970127fe1f581b2a5571a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2bd60a234fcaafe50b3bc5b338b4c6eac93404bd647d15e0b1e09f150a8d7f767657686066e108485167c2ca9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98e4d923bbd7264dfe54711f9010f9a6aba70e1453dba1fcdd84f4aafb049acc8a36cefd8b2547f6334618f8dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f6af2a22684eaf6b5acf4fa90dc3f1d5c15082359ae22e3395f5add0fb0bb4f0f884e88c585f47a399aeff7e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121e04fc4d0592abde5ebae54aecf98426a4e140df8a8545efe8734765674182ca3eadea1d5073d703da5419ec4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d954bb236e4843affad63c157b4c81321a0a1c31fe317e796897d1fbd53bcb45f1713a99c077fa42534e7fb36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ed046f84e25dee1fc546c49e6f850af0b0a83535ac6c66f89798ae3f36224c151ec2f7ac3a971c62fb3770f7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e6b9f56a90ad4c59fd93ae2113be2be58f78ad296268824ab6adefacf4d9fd4c99060e002ecaae1e655bd567b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1854444c537b26419045234b60eb33d8fb9190653fd5ed6cc40fbb523a2ad284a08818dae9b19aba82e795d5e2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d05f5b4823d25f982d3c3b623fb0d3d1aa0ca9b8b91e656ebb60c8fea13535712011b21c2916a7e8c4ffd50200;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128f63f2844c3403e1b19ada15c7d8ca7a4333eeaecfae79da3ba397a18e9b96b9f3794cf39c0e1db67ee0a03da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3794116d4f787e7fa25270329958b215741cfaf4696b3cd7f6f29bf9a412d81a8c45a76e801e5e13497c89b008;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1050248f4ed5e1279668de4a947cbf632770031e6f68cd73d0c2ea7d4af3c3630b49d7e0b81ea30fd243c3cf55a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10baa5e679c77e10b164a8cded9c0064621b77e7a9afd6c6092a9c0d1bdcdc12345590116e6b175d81bf4ce29e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf067fd5b2aea8d8a2edc7c210391e7d4bcb6794f3d0b32eb3d04045db0d7737bd576db6c4642983665ee9925fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f6e3eb8aa927fbce59de37d24f5ef4b313dc0b697aae2916959d5acff1cfe66ebe5d1af7735e8a0e0f916a9675;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121b3a57cab86755a42f3176927b6fa0022f550f81e6a95b5795204246597ddd018a209205afd51377611223871;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1300fda296be92cb251f599a278df0fa2d7f8cee68fa53f5dee5d866b8f1ea42715fe9d549b1472803ec7f432e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10af9504e7e59fe79b8ef06c8688ab65763c9f8d823a8d3ec952cacf1f1522dbebf4d7005a42271bc62cb657dde;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b58c15666b12292f57a30903049918fce4525510c4de4387e72de1df4ed200468db7e1d89bc1ada81881a2d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88f5ff97f633f9f63506a4a655c8b5be90bc0f3a909273882c267b7829239dcc7aa70eb6462dfc2aaec4af7c54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e5ba40b6893eeb760fe4acfd694f9ecb0e343a149be64624b85462dbfca5e7d433a7870df9b1f0ec5fb54f94e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h634a21d72c300be30a383771292329f47411938f61f7a6243d79bbdd577424ebbc213d11d224390e814e74e6a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbfe2f6f464ace846ab8d889ad4ba789267cfef889704e78e6092ff892f2224414d946441a49d5d927dc4edf5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10661e5c9083c3ee662da24ad267632a7deb71b9da95674e752dbbfafd941a986093059eb57c96f8b9b513b8d59;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db5f5c6d2b95f09d463072dcff6f531fcd0a1890adf528281a51740c834909dbcd9318e02a4d9e298b3870b15a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4b6fb569a3acb21e571875c24149f9d95fef48ab97602ac98bdbe934478703ef3b419c63d5089d3e39dcb5ffc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f1aa3ca6c1ebd6abcb8491530689117d3647d63eebe8ec55ebc22ea5d76d5a547cc76ea3b0de2aa46b78c7210;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80d49894f8ea0c7404a4c72e35a3f766255e130aa293482c3f1d2d8a4f21c309ccfa377b746a4023dd1b3ccbb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174a82ba353a57a874c5acda52a90ec6d60cf312254c8d19ba14817ac3a431b11b29f96b1e078745f5c44cd5d98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df171b711ca7495971acd400ee369f8e99acf7d94ad88ce9b5805146bb25cc94e3ae926efd11d064d66736a545;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd479bab2b25138b4a43efd83388dd919c6799314887252e8821ca4a87ccca1344cc76838839a46957ad3328c06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f996e39c8e2b8b6ff264108145ef8747b8a82112138c1cea4d5009d936eb498a6c583bcb208f0bc29c8208838;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h702e8c2274d469b17899eb5c951e11e4371625647cd9ded0c5440fc5147dbabe846985f5fd052cd9a356eb841;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b8b37b1cf75a1c21c718019c8409483bb4cb30a33a16531dee710771c6c939cccc21af29a81940fa7efe504ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h454175a0fb6ba99a621decf3c697e7be72dbf36cd965892852bbb9c6cfcf1a1a3c259d371d74e1733fd70f86f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee037b25ac407e060f105397b53e2418181b41878140878e82d4e4e914c770891e21314173b2b8fc2c5fdfb891;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a74377d6319ae2ad83b65e4f756fd4684849923f565fbe77aa11e498912715b7daa9f7145abda100e8e16d4ff8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he498c0e3bb4c9f3ec72557e9f1f470a6c085517e290dc7df132f5df4c336947fce027a4b2999d9a1ce8c1afdc8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f84f6acea04b7e5180eafb4a000e2f39e956ad5b5a77c78537e147a8e9ee61af1e0f8576fbeab209c8f9b1345;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147d073e52aad0add0f57bbf013b7d75a615c6bc5d5368613d42f0fc461562e929e6818936bee6aabc69712e83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e68a456ed5126632e38d84a1b9eee503859e4e840c61d4ab5ac8a5405664be53798a5aa677f1bdb10f0280518;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94ac7638f88b2246787cc1ce782a89ee1335c73ffd073d762231925ebe5b61d574f4b4b67355290b5c5b0dc75d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b1c65edcbc1a205a56529f3fbd42b3dd0ddf5f8a23fcfca1a1333367636eb720a4929c867d4f282fe1a899a2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37a7d320ae636a212abb4eae9eb2d2ad055921b97e451eb76893488f377ee0a7a62c148af5b66d16d8f8913b03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c45773447b6dd64b7cf3cf50661eea56850f4b0a323d7973e8a34e8c249bcf4d751071e766ee4259c082b561e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3465509a772023a0fb711e2799ac96caf34edd08c01e3001f62a0c1a751288cb72eef5dfdd9eeced0c23be0d7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dec2cd3e506839cb19fd99f10e4e82973104693bd39423d7e587eadc82e09597cbd966f8ab8a62a40de93c945f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179e2c339fb59eab83a35c093313824485d78ae75d8b70103dd1aae0a7478266c92650eebd281540e53325ab2f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hddfac98ee8d8cc01d89a6205fc37574e59a949511922e45c0c08f6ee0ce2c6902b62681823cf8f76121c052979;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146f82af806a966a5c4250cf372dbb0683e6145a70ab6cb0c3f4013facd007162dd1151bd11030d0d56f9fa35ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1cce23d6429b51ae28131e009288711323bba8b65a8b2bb5877f7ee8e7e0ac0c4a74fbcb69fe9b7865494037c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebacd9ea251f35e06beb447277b67eaa4b7141b7ad38a19432610d4ca3ffbfba485f556c6118b098d8af38174b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a77059f5d696a1f7a5e4c4c4c97a062a18671c03780c419b6dd18a997f5cb0d933e8ec7db0d6390ae1876f6d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106d22bae1504897eaa32f0e915af648a5da6a6810f78b403c3d00c380e771ea9a864658372bbaf82ba9f9b60e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc814e5b46f5bd0bc37da56d840737e0fd34a0ebf5cb07d00c8563098124c047dbeeed7e1571ed7850e5bb5b9d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147e186d1b4dc60665861ea0aa4e86d2ee629f2067e78835deaefebb1633d66729eed6e24e09940ca5fe5b97fb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2e049b01667cdc59e33f46590813005f916ef224621c213dad58ecde4881a654506a0c9f852061b4e87193ef3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he61983e6dd0eb1fac99e0069075bff054bd808be96d9be934d21269964c47a15d79962f914d9ddc44754366246;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64d7a7fae5bc179a96c6d1cb77afdb0cec5d6e4ba3fa99ba95a46888ecdc904b3cab9aace700f066afb4c8c9b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1cf93e46239ae5a4d8c905becdc4ff875e762447503893ca70891efc4256294a38bb345f83376904e14be5499;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70c965aa1fb63ae248942507ecdcc3d0802d538c2bbe9d9d3852bfad30e2276d0203203ba31c83de2bb4943193;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22c838ed1badf8c237eb1f033be1fd026b222fa491d32200f2fddd96fab2d9ca0df50f22249af481a273be1159;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6069186ebfe04de9044284a67bb4145f6b6af7f407eea1cd56f3f50c2b08275cc9a1e828dd307845a5f89e6a8b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h350aa399ac8e8a36568451b3879d7d6707f0c6ee12e1db59ebab05aeda0ea5c5d2427460a82ba7aadbfaa478b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193704ead0695af54aa84d087233e81c3c54c118336518451cc5374a77e94f15fc92e7e5318937eed0c5e94d07d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0ee130572f8a7ec119c8b305d076b288c823357912c7c1ab67f3e99da7a5db1e30455b518cfea4cbd89ab74ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167a037a0776a506f85f0dfb90827bebdc811275331a53b1e0003e003ac3b49ffe6cf1c870e29856d8124f2f3af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdcfb78085e4ab72bee198d8fad3f7d91ac070958e3d20ec6f8d86efa44641b30283118938a954d0376ba7be95f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8a8a45003718a3e0ce69291f159f46536e5307654a8b64ad92a1c64e3430808f2eada122c679c801d4bd72446;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26617764a42cf71a700dc0dff470ef76c0c700057bec65a0c54f536dd618ec7ef4babf48ea28ab2bd5c0400d05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4c44d1d9b272fcd6658cf4806dda821aee4ffe60a4091d977241e7c84f14456bd999bf539a05ed9a2b17baf9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15527ea5498a3f0d6e9fc2e19b9cc5ffe04a7da0757116fbdd7b278aede367c3ba60759785c20853fc4f436b9d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcca2ffea6f07164b6263d8a218ffa1e62a8de9dd017d8ba5d4b8d55efb987ce52b94400bf91f1d9abc7afc85c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb625f65ff9a848a5b659fa482c474caf112f9efb52e56b5956f833306c47fff57012e1c452f4cb895163069392;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c8e5d10e40599331748831d4ed87e38ccbb028f28e521d9ab2c5aa30d0a64c4a532f05d543b1422627f11d57b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4621187734cfb2e8c45d327ccb50d4918b7fdeba9a41c29d5925daa1b674fcb216a103fe56c0907d4de1cabdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112fb8c2886198113e157033d631795b7bd3423005a4e7ebf878fd268cd49cd365e974255d79e9bec9da4a8ac8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143bf94e10892748dac72597dd741ecb3c88eb0fbd7011fd442dd86252c7b2df028230a8f9bfffa2e822866bf7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a1b4aa6ff344ecc052e7f607002c6be580c7e74b0590c9ffb875556e62102c8010e0a05d3461344bb8267af7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191fab04bc095fc50f20ca95276626dcf4f5f913834abf56992270e19bc45a73164e0491573fc34457f19b04989;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34f4b8817ac299bc7108a05cf03bc0033170a5f77a1fca55fd48f897e1287fcad8acd8ff914420a23571a91714;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a54ec7cea777b36fabb425eb5c6ccfdf8808660f23be20f265da206b25925ae54d963f8745763f0cae2dae24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f11dbb3466d629a59e6828fd2254a9b401ff6866ee6b66a1a895431c289cd2e23e7aafdb526acab8a75098e738;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17188b7e4e6234d6a3a7a80a6e07537d83f794f9ed24ee6b4a5e52b23895ce06d2bfc453a8ec81a29c1f34c0054;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e89d186c705431d16d18e248f4949a560df7fd8ac0c97297f83dbe76f640914a4121d6deb067911bb33dc5c22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146a927ffd8059ca55e81dea9494ffcc86ba201858d5ee340080f110448cabe5a38ee03984ecdca4af13b1532dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8eec5382ef0461a9d7a5224aa6d192ed0a7488552eb0c5bd9eaafeb55f4b094efb924cee9b458359740097f612;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8fb5a848058adac95b423d1f2dd323c2f42976f5a2d4ccf1f67fcc2f18d2dc055a22e4010cb9a1e2aef59489d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18830e238777efbd8fe9cab920c5f30f607c0d836002992c9ab108afc7776beb11aeca49ed9797c288fc938259a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha420bad0d2c1b07c0a09987dc8b2bb009eea1e23680a034d0aed37868de16fb245ea9be39d518dc3c7b9d79b0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1103e75e8afd085f28fda79c3d9214e4a74a592e171d753b89d1b902fa26b2cfed472efefcb78886eb4a8ee98ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afe9edfd10510820d7b818078fe8d839f06b79b29cee54d501773a898dfad04518c3ccc2471af69c539ce7d3ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7e954d429f7d48e289aa464312796985549d60176d8a7c91cac50f763b43197731322b500211ceb7bdd377011;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcec73d4f3daed42d3a6da1fec87ef2955ba2c8363de393c10a2d254cb42ba072f0b9040e40e25c06d061c9c568;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e93c70c148beac9937529a5b8997a9fbc7c386045eca4ec80d45cdd6aa30ee71b69ba0974023b4e2055eef8eeb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9019da7ebbdfdb0b9b51146573523d379efed0a9aadc8c4934c09737cc45a5b2a17022dae9cde64ea81ca05fb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f668c02cf400c3dc1ee66c9797d0ce63b30ebbddbd30c4bd17b870f53fe2a8a1df896f46f1869ceca1ddacf99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dffb952b2043a82399c4f4cd81fc9b31623a870a2d03b8cf6d501bbd757fbbad4625adc23d09ab01ff41f2927;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b1efe1cf68b65e721277517d964dd0cfa6d38e7fe19af1fd50e95cd68650121f12628991f5fe6057fee721890;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131a89e529260a4a5487a11fb0d2aed5c87bbc46e133afaff79c416befdd2e200cc74eb79189582b8282adce7e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he73d2cd0821d501a5277793f7ee486499c08dd197fd94304f6596c8daba1470be957fec56fa6175ee1907ec6d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9bc1d27cbc3ab5cfe5a9bcfa26734f0a45dfddce9f64fc52c85e5d1e6edff42133d8b4e36816230496619039f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8a1bb6323e4ef7a94335d2be4968d8b6e722fd3bedfea05441342ca95474c6205150e33814f0a094ee02bd63e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194c2bdca084b8ba3c14d471e6484d736c0ec7d29b1230d710236fa305b1be43ac07e8ba07921201e09994e2d4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1981345a7dbd2c5bc24037a034049336d079478a87639734fd2e2f73e1186f4b485acdcf63b25fc2590b37803bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de8cb0fe3dadb4420feffe22ade16059f231a67d3a9d7140b20b4c4c8fcd628e6d4a5bce818cafc79096db1b47;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e89e0277f0efba9dac788601d51ad20d3f52c4b48ebade6616ee90bf40b1783f6852a4da37d55be19715f142f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca0f5e1b29690f840bd121a1d127d315c76ed0a6140c932ed94b66e125366df5854177195553ec1cb5c9b8302b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h715ab479ba2cb7bcdd53f4eef86fce156b3504cf11a90639a546886273123513d101cbab05010828458e85aa51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'head6c1be659380647d3d8dd36fbfb4ece1f0d2d0a905e9907fa4f84f6419a4bae9003b9c8b978c2bde1a27bd57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2303f1a3491e211f2529a5f166dcd66a5216115f89dbc210b4aee28a81dbe1f9aa9525fdccf39b79d043ac78e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5934d52a8f9e073e38bad133db1c37daab425bd1040ccefe12f07a5aa8d53dbaf80dbed2abaea4f5e64d3ac51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1592510a986131b1e67d33adea44690ad9fc072b6efa9857cd55e2a6889cd5d0babdac4a21d5dcd957a6914b96;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11827f1cf9e05316e1bda6783630ed5d92944cb2d59f4420a59c6218eafbcfdaf1b1c7304a9677605c531e365b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa80a2e9eb4e2e613f6ec5fbed344a7e033e3d9c3c7ff2f6981098c7e57e518b09ce6456b23c85aafa925fe646;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1b6f86268c30142914d7e4f89cee1b279feda025ab9d79a88c42400b4a7d0754923e9e20d7f4e151196a7fa66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h552813ec4286bbef86612be4f95a8a2554ee91382af09123ae51a2ec6fc2934fdc72611aa5c0a28fca836f51e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1983c3be664b6bbf4b30ade2aca97ff74003e3acc09d18665adbdb1d0889c96bcabd16c11ca8670cbc23e68f034;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c9f621491f5393562fe14a8d65fca84674f0e8c7c21d5ea6fd4e3214a9a57be716ef54a78af3e5243cc66c68e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1162d59ce61750b00f39bb4d2e4c013a566f34970f362adc144934081998ad76b5ee70b0ddcc4e05e0794361c10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f756bed901e2381291c8f3075bc8a1386a4b93c02439d56d0c7b0b9d8612488d64be4a027b8b5066d79deda94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6bf7777ddfffab0cec1998ec3c88dbc0e4ab475c081e9b0201464bbc4be099a2b098ad94a4a91b83896f8a6724;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d9250ad0a9821bd8e40c4d0b09f0b64cc5832c70f507f965e8bc4d7371cbb137fd649edc06fcbb8dce42161fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7b9ef1999c67440ba5f628cbe1d5a9964ff5232e333abecc0cd80a38ff4ab6bee0e3d2b6aba5ac138e3058687;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14abed949b4e9a1f2d80719bdc362750e7380ae7227ce7550cddead5f8ec56f890d30ed70a0e678426be2673cee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6f0be6456d03f430a9a54efb35e5ce48b4d914f94fd18be4d0885217ce32986ee55965e5459a86829b8ab5811;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8aa172ce22f18d4726eacb860e2058d7ccbf57b38959f2413629e0a999413544118af5c8ef12032f238b762a86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e46e4c5bb7ac05e0ac63db1e820a10d7d37f6c0bcd3703f0af2991034c24a748cf1a83b3d09f69ca1ae95cb3bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe3b12242d94c38b32eb152411eb26a6170db78e8951a86ec21315c7898d69ef0f08b3c99c78f74e69387c98da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103da5406842a954f45408225515ded186aa97fc87ae1cf5163bc7bae48d0bfa068f6df5421c09b16da5d80a730;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f1fc5ef86e297558d5f9b860dd9507859a1ab1cf4f8df0cad58068ab718faf70608faefe003781c085d7ea1d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2567453ea12bbb472dacf38a715b5989140627e8af14c369e89b641675872634fd1b701c6a6b825b767e3bcba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e8fe1842514269a58d25b8aa88e7a56de446792100acde31303af1e1f36687f5ca871e6cadc1a3d9b4ed82db7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d8fdbe422151f8af62f061ac33f2da4603ef49241fbe7230efc4243b4627390fa8d588156b45745c55a0036e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14effe8c9755988b2e96599b4d2ea5b118b470c9eb7686eedea381300ab53c944035eca219e1330b5444df628fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f05f261274ed0644d180d3a3fadfa971a5b1d1bc5fb0206e198304f05ea49a28a252ba026dcde6645b6bfb3ac2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20585b7e16088f78d121ff97f79304d076ebe5b04d6fa60e934a9e56c6534c8d290ae3917ca2f080d8a3f4dff6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e18e47fd19681ec5f877d7d920f85e02d560d198abd62836879dc4b3f0cef3e4ef66fe4e7e311578fa0f5adbb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4dae58bb19d6cc2ca9e96231972c2f2e1341e825222dc5ba7fd6fd425f090a7fdf0ca2d3954488cff73517225;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17837127d562b5441003d7366bcbbc09caa88c1ec364dc6fb49b5f69946b085ad0977781e9e5b8a577567f5a942;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c8f8e53d7b965a2a29b1e7b1a6ea9c5463903788d080586fccc16bdd0455a19fe21a641b6333d7e579a5f479c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174b210e8ca1ea4d51b47e56e44835e32763ecab19155d9c25d6bf59ca88b49fe47bdf78dcf5afad176951024c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a23aca403a5e7c5608cc9305e25d1aa1933e7dc6dfb0dc93a88797b0398ba3d48d874625669a5fefaef9cbaba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f90b3be280bb593e60b6de63d77f4702190cd4a48186f12864022ae3d27dd13b32562d42733ff62e006377df4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae0d8651a31cc44a38dd6305d9f7c9950e4c0a9fc7a018c81829381683f9b2eb8791b183eb3e4b35942854d495;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48957b364627fa53496a31239da110742ba0364a45c413b7eab53843217280371c9ec41a0777e3c3f10a205ac2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed43e1e1fe994c95b42222390cb240efdc9908012cf94599fb3c4fc3f05606aff50434d98d4e01ed16249c0a9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d16238032cdb39e78f8f4de581098c6a4fbc32d35e083d08236449f04c775bfcc0d12dc83f52bd845648df3e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b16b786f69c182b26419d019b6558f1ff9f2c01ee2d857d0dc2c65792ba77f979eff4ee43667818653bc031d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b8aae69ef1c4a0befbedde826148417246825d3ad47cd67f558d81cd32a39aacc7bb5e2620a8663caa87939da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117d7d18cf9274d9216d41168c9bff8cb55bb4e223a9aaaa4cc8f50feb906e2ba9b033c554f868001881b54bbd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17853bf70896596df04ef911436ebeb64686f63d5c19c6ceb6173090586da9df773c00b7c453fdfa28f089b4a85;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb632cf5405cab58b3ab9497af5a9311fb3a92ee5083064e47ff2030a473f8145490d1707975d61145f2dc133a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ee2c52c3b7b10e2083a6357cb81da3bd28eb7fc86c403777d62de3ccb737f3fb81785d60ea66a4e6831f402d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec0d05d77eedcbbabe98c1e7823f77e5c0c1368d9414633be34bdbb3a5b604dd42cdad6d3493023fe5a733c610;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11304c909cac95cd445e18b82a1b7c16329a9295c92a361526f59c7157ffa9429a3515ca089d6d08da77ae6222;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ff4eaa606c7f55552aa84e123963e23bab0630ef83240fca34a6c460468ba5f7f811b56fd1502dded8f73b9d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he83dcbff6ee1a12d46f5b0d8fc7f3835abd049338869dd901be7ac78199f38686d0c19430ebf0ed9ce44797d55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha69a74f2a322cbad0d570ba5da8014edfd29cc3dd78af944d16c3924a5718ca2d55dbc4d99491991e0b6d4e33f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4b5810daa4ddd24f6033bfd479e5bdadbf6d1dccffde050a524025daa2a61a1a695c8ec4575eb579fbbea56c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc98e58e32c1a739796879dd8eaff9df8321eb855fbf7e5ce09cdff1b3624ce06990bce37cf3ed85a6bb9eb8abd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80cf189d054e0834fcf2a3e77aaca85fdb9b07a1a7eef6d04a88eaed9b375ed84629f07b612749f26f10833fb6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3d84c22782062e14c52f454f9c7897aec14b83e25f1769f5f1b66242773818056d94196119b4cea90f0b81278;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181b60649756b93747cec94cdca14d11ab37f68a39e22f13dcc21383ae3bee4c67461e19b3ec1a418247b29fd71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h762d826031a423ef68d8bb1f5c245674c48506699413bfdcb8394a35fe00c8e680fe281d153ef45e5f549f7571;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf05d87113ae205694e5e5a47653e3c25d0593b4e299a4744674ddea56ad9484024f971e2d04905483dd39916d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1305a8904bffc09a7910c11e498047af0c4fe0f9ffa0afb84a2f8b7ac8e717b6cba522cb506e22f4bbad05fdf7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189cf4e7f97706c2b9549719edb4ad57a9afbdaf3347921680848d01be1c7129cc70454c515925d214f94484324;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cef5b436e2b11c7b17ffec74c83fc5b14b25e77c858737f0cfafc0297c79f7c167e693d0e5f7d8b1fe3b6fccd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1689f7319b8b98fff38ec8892b6bfd5f07bd6dfe775e8c2d8832e6eaee0c0c28861e42fa8fe3541a510d80774f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h848eb31b1f340e960200718906fab5ecf1ff9a9550d9c610258f8debcd213fb6d910b47dd1aca932b1be26a719;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b37639444a8cc6c80d3cf594e2109a52a77b7beba0327c1398fece00d535e8b70153dc138b63bafcea9e3a2933;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1adb14a5fb45291cb8b59988a17c4856f3f377d6e226187332a8c800fbc91982e7fd3f0dad10c3d97343b2ec0b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h869f5c4fd2ae4db4f5d121c7e8424ef619df78c571fb55b96078e640e6ec0a4b3a5a5984d696388b6c5c9458cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11374f255e8b42f70779e17fc50df891de5c3bf777f6d8b73b1575327b6c5a4df4b845cd813e3595fa58a2ab9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c66d275caf45910ae4138d168f8565418a1d1aa41c491e0d972db72f480c9831d9e9388a804d417962fcb43dc7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94ac3e719035fae9011aa148e26eba1f87a387f3dc7bbb0ec1ce1913bd587546f08564e51139a8ec9f351c74e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f611c3454d7f81621e5246719911b2be5e8e9f6324bf1e20cea7eed96d3b63b0b1520eba769b6851d6f88f73f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8daa9f952ae2b172eb382c7d49ffa27c1c906bb96d1ceba200478263bd1c80c491035d4272ecc27f4939ed6a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f751ba253710330b2e0f35881d0a411e4d556efdc795d1370e41d58093b7f0fcd1898d6d6d9be3d759d5bebc4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9531c86cf9f3d25546b61df6ef84e9ffb02cf95b65d9af2f1644762e09328653b5840beb98421ac9b61f54156;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcce12bd27a3f25714555a2e56435a0c73027b1611cd4730fc564a39da01b4786032349d1eda378fb808831608b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fe73d48e8e515d5eb7c1c71af198bb28fa7d250960846e101e4461704db45c498e9452cef531249e2ba32f75c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c50d45cefe3b98f507c50db5ad9df546f011b40cabff05d541a8968589782757511fae30c75557251bc885392b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126d7c664769deecf32f5c593583a889ce483b63e389c508efbbb8eb43bbcf00d5b3cec2d0d23d5dc4617e29a17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ce5b5e64ec990972e656a718d6f55a94d29a5df22c848461d300ce70f8a55ea5cc2951797c8770f34028ba0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb92d848e0d75384f600dade2faf577c2369fc33acde3300442a5b677e4cbb326d00fed47defc94b4a72004745a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25b20cbfbca347958555914bbb11e6e10e2356ac420307a8299980934fa2f12494a5321842c7b4b0e450b1a0d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9287cfe6dff566787b10b50697fbf1350c4b22c0247aa517a3402bae8dab8c914b3767ea1dca480b4304c8d3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81ae963337147d606156c4f7022f520c69bb3b9bd299b9de76bb662b6f99535317141013bf8b2af68f5c89df66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6a9928b1f2f209dbbec33b5a01c32820ebcc543cd07f500c08dfcff55494e278fc9a01fbbd972d6a2dff44462;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd2f0c1bcfece3555e1fc065b703117ed433e544cdb265c5a8fc8edf978eaffd15eb05b13fc9b85c9b918bf605;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he66aa4999943973a2b8338b5f5972dbdd00e13fd767a9df6ca78b1ec71a8277bbbbaf6f9e9f58b1fdf03ee9afd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h750b320ef78ecdd8bcb07482f85833f7e9ac08a1dead3be50067398a59f51a0e3385ca8db1f7bffe360d6d4ce2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b617a7c72ae03376d1cc93b6eea6a4ef59191bc8318581f78154fd06dd902cd71716e4bd258c4e99eae8d8c83d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c40ca5e54d74601a81613cbe50b043a73c4506e6e4ec8ab4221921327958ea8247121d7eeb8ed702e86eaf9d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef8261a991b0722f65e906b83926de6683a4e776f02bf1e8a6caff712833bbf7385327a3440598817b3ca25022;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf78188769314e3d6fdcc388f23ea8c4aa2bdf06395f24abfeac48fa70176be02050c5196e378092c7c1efea81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf23e09aa9cde23ce2e159e437f3443189acfffaf63fc5c9acacb23c5b3209e850e3b0b2f6ade3d542a6ece6f9a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d9c5da6288391b160e632e392a98de13675ec9f9ba6e2d30e173599c89636eff26c38653bd5bd53d0fc9eca77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f153b46a8dbcf4f0a89bba08bea75c17532aa99aaf18c4e6527782137011f64680f3c2de7bf779598998bec22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3a16c20f1d9aeb4d151304bbffcb7a06cb656a8a53917a294cfee4f20592dbfabf6b498a0aa2b628511ee513;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h649cc0e15429e1e238d0ef26ddc95ffd5a229f7b4277c01480a39a8578814d2b21bcc6e686ee14ad84a2a9f32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99ab60ea5f34e562308153e0b84763d2eba7f3c94587bbfaecc8444f67a91a4bf283c8bf98e0be87f81f4b0576;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e5f11d536c01d012f15df81af9d642e092c2103ea78a54d66c1372f857333bfc77fa5f5d086a2173e76d91ec8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1405cce5509b4287a87461849d0d88072973bd59d2a20993ea1b6f80ff4be78e3945d87fe7c0c4155a97feb5a40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0f3fc5de2714c9a466173304496c3942663dd8ef5e361620758fc7e603168c0e045547c88c216332f0afc161f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb34865aa2328843bb051e1f0db5973b956aa7de6d7030262bb91a2131e13629fb0ee60d438ba98e8cbd9cb7c28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28a807c764b109d2abc8e3336b6caf0dc9c2cc9309f35375372ec449465df933b4b5fc3d78177aa45b12764c76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f14daf783f1743157432ccea46e1a422b5148f8ad5bcace5d01db023df6cfaff08bc814793a61bfda05a78b145;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f74f6bb7a206b365b6bee608996fb3de071737622f9ca243665e12b2d8ac157d418f629a3d8526996be43a2e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6795407688f96e1927de62760d3969f27963926cedb742dcd11e04036d2257644ea8be465668cd23b07d951369;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcb260422561378211bc9b299b3c4c7cec1a633d3235b6cefcc66eccac647b8ce76f54d93995e4c0db5683cc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7311d2277db8e9cd0c21bc87d0ccc74aa7e3e74a036c67e46abd564a777602a58167098f0a2acb7ca6f0fe8dac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf6ccaea5505c888262e9576159d505c4d5f3319332b9606d07e11b678600b48fbea41bdcb2a38700fa7f42720;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd03ca4a40e7f5b0b20b932ad1bed016daac8777a1c0b297494cc88c5df1a281100afb28104799ae89447d7560;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46e2397cd6da1e1c5e85dbd779485cb21bef280b9a5dfb033be29b8daeb8a5432d9a6411b7b3330a851f6a58df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1603704501e4a3a3fd7e3b6eb5d4c43a3174aec48bd9cd3dd063b38244d121de1301f84fde79300e3d1e1a13c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e435f2008131331d463d14fcc3a1fefb53fd02dc9bfc479e0774da3113f171c0268deaa33eb6c9784c7deff7a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1ab363357c8455ae74323ff8832a43a1207e92bd6a3bd6d3b041f07377688f0725f0500c55147a562e18ca45a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf8b7187a473f6bd81081ce63ce97c102beaf0349045cba82f491d90ed60ffc00e830d3f13b4fe4a6e1a53cc6ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178eff7027aee34fad4aabc143b520397cf3b3558d1a2e3ce4e7565a3b51e300fef404755daff010105b6cc9635;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12687b92b3e9aa340c0831a3cc130c6568da089b97ec1c400898f2afd1812fbff7615f67b5070e3b6fe2c178916;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eec72f0287d8838f8f5d103b37bdbea329152424d2f41984bc6de1b405f2b9ff245e50bf8080b115b43e0fd62b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb4348a6063a8732dd0411bf332429c3c00d41aef0ee647cde3de936f4a145469991955b4d161f55f4356c53fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b39ca0074bf0ccb7eb547f48cf96e6cb71f3c2cfb6e776f0d9844f3c9b0fa5eeb8353a838f379219e725117778;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h242bd61e0c9a63cbaf6dab8c913a1334299dfbbe0dbd9521b7abd68613c2ab0d1a3a10ea37cd560c3ed315631a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha88dd8a102bb111853c1637964aaef31f5c72faa3d0cadf2852252df5ed4dba7128d8e7d1601c6d33a86edb3ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5dc648f61547eb9a01a1c18062ba96a839c8d9ddf367ed59e6c779b5238ea95181529b2b5b4dddedfe8c2e78d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfbf5fa19f51c7000a9323a5d679db87bbea90171bd4d182e973f9ace6d20af56b2e26e18ea686fd8f631b75088;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1b31232b264ce288bed716a0229a5a2f02534447f6aab521c880b34badfc3ae870bff78261a47e619dd6b0d9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1319df3821c96dc4335b110f3a1b32f90b41a0a378fcb3d0d9cddde36627e47644a86d47dab0bcdc9496dd592f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h157e4a1a774f341b0a0c7b38303358a078d8fb0b64a3e02d49b98e5a3527c3de6ae2b644153317fe89c0044a064;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a292ef67886284889e09b29bbb656b35d8f2dc796733bb17643b00de7d691077522f918308aaa2fd645f6b3e23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf8a65193b8522524a289665f469278d399d1d98389ca46346ecf7e13b08dc45db389c700e32047ad540eea60c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7eb4ffaf87e08b01394cd9c96cada9b0f05de89077cf8d125a12d1d7e70cfe849a629663efe9598a72831dac4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce6d0502a0f1db2e5afb940d733f400701d4a57f725cb7ec6ef0077314952197e57ab67519fd9545b35e2b1cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16806e6692279eacdad76fb287c92b9f8baee56196e0beb098c1473c9e6b9d25c85c42c4e7deb224f7fba568f23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cac3438a9d3c5112f75a5a91ea984d8f67b7d6ab483c185e69e9fa63e1364352f774c9755d63f65a7d319cd1ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5839a8767cab9686a4802420b189f5e64ac2af94aadc64edd5a1debe184f7d06012cebe944524e0aa1052dace;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47560008b564b101a1d9dd6e4d02e65464a9baf3336f817b1d88e279f02669333c93deab5c895a2ed148ab1299;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1837f4ae99cd5486732fbc6ebd82e255274fe8810d2d64641e4119b48caccde247fefc0ef59c88df419332636a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b16a3fd358438d08c6add1cf3d24517d7e80bfea39be4d0223826d21499a781ff7451f52b84a3f027ee8ce601;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf3f354c37d62aa39a8199c17537e6277af7e019218b0ae676f3babc20d5a4b39555cd4c4e03775315b6593867;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1201f08dcd09bf693654a4300e2fd9230ecacde920d67d195014a5fd71a954dda963998406626605182b91e009b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a6e674c720dce8399aa2de4d50b2390f28f604773508d84bfe5e8e33ea5a58268454ae3752ee3a1256960300a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb11178be144870f3e95f3c542fa343400672789b6199c1bc94e9817a0402e77d1f7bf5794130c0b247fbaecaa3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d169365d32fc3457b9f835ee409ad15afb5f3f06d76da8f09a577e490c294ef590859cfcdc6d543ca97529333;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b117272c7668095764c75678efa035a770101b56ccba6fdd59041dd81867690462371c339f5c5b1c68932eb06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17dbc76a1f64ec46cd0f42867b881af668dbdb5928760692eb139439b53a684698878fe4e7d251681bc1e3b289a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11996fc2191d5e49151f6c2fc277cc1cb77fad8bb3de387d91c954c50733488bf69d4f6c6ebc8009293cf3b7f31;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h255d3de22077f80d358dbfb5837eeff729ec8b9a3f9b1040c3e861e718c1e9e420025ea6980db404cf18e576b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4882c4d10b43be44775f4a38cd41571a701b695c15d5df09275d5a6034c1c5b2194361e43f3d887c987c98b6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f053e5df5736803c14b96e0dd58342d08ccbd22b8d8ee1d639baa430b3a2e4995d2c4be907d1f37012f7602c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf655436b2e3598d59f389c57a64ad3e2ba1937899eac93d0b9d5f7a9faa01f4570bbde0f0e0428e85437d8b4b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8638024208f1f98dc09f7238c481b5512bb4c80a9c752eb840c028981c7202276b838e4cbd25fa12d02c346a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1080d0118403544a8477a01e582114b08d3fbac5af11acca86b9ee148d7a43dcd0e46042b82483387622793671c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6b01608c5c6bea1b6971dd1f18b57c4edfe60a8e7973bfe35a63730ca0ec6abe08f2cecf8130b5fc97b48640b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba48d7bc55601a654f7e92ab5ab7918cbb3e5b7ca773e450f324f3da1c684dc1a6b14a89c66d7ed19bec71a1af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14495a4b75a3c28a224a663d7851c0ab264ce7547d1b1b1a7951ff57807bfe2872b77dc6449458a21cf429aad76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa6f229152afa1851bf68d3bc33c4ae3419e90f6fad24c2b06cae5caac49c36bf0dac32c6fffb278fae9019c93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2122fe2d77a3b3e4176d7979b716a751ac7722d1132299d515a7025eb916505227b684ac1e64cd203fde22041a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ae2eefdfec80eac3f087bdde170d65b019c7a2eabeea8b209ed744db2d03346e8118b867bd952f3e84ba05442;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22af816368bb3964b7f233f931e138d0807d7edf5d59e5b0f3339ececc66b6c0c2db72ebe5e9482c719467a960;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c06a124dc4afa7a61511e7f9956f35994241c551d6a1099aee3832906e41d545b4df18a5003395968fac9048;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58b269db9a26364a8c584d02a708ab30f5df25ae6218c914ed6a430b389a27d9dcc81e9fe4e9e1a45a4fa23d4d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac927bef63da13eced11b12ded2c85efdcfd5cad3ee4caf5abc0e6e5692163337a8fd0d6f530092ce1868a0cfd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha76d584bfd1dbbf68766ccecd2cbd36c74fb5b61d7a40744a3834c06141fb1f0bb1932cf05dbf14057c2c4079f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39a4212500132de1bd169fa0e75be0d1a338d5b9ed4fd1b5e8d59b5ff0c7dd8b2854919ee1c17cdd71c5d952b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebce57135584346c23886e6de1350f23163d291889ac717798b4a747cd309345ca5d2fcfdbd5eaaddab2bd2d40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h778f2c124059ebd94ff86bca544f4b821015a55cff1565997d5e53554b3d70f85917ff52929b33548f81dd6c3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fbedcb8e1e2e87806528811d3340489bcf629c0c5bb353daaa47215856f057d44eaee48e3ee0cf22d9253eb53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b71e1c73178c6ae7d4b8c87d00bc8975460e562aa8fa9dd0dffae1bef869017660dfba09bcdded95e58d8ff0f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h894ce83068ff9fd5b98c49fe5ce32c6e799cfd867defafa089c7fd7e43f5bbf3709f0012f88a8d2767f4508c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1811cae0a89757b902ac74683d57fd4c14bd266a60f25d3da1f6c8191a746cb2d90653a290ec20d4dac8dea34cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b2989f33fa175f0115bde9e32a9ad25d9c7d9e220195e822331de4afbc430072ce7add3ee198c2a1eb01cc3a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50f24ad1c205b53a48eff0e87446473414b0ad572f173aeac0cd17c4ef4874b7e0b0319df48fa9e13df2f596f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a229e5bdbf2852db06f0f45ff3c5e09f59fe9eb28a07228dfc653822eb0ca663896e3fc31795fe319f6b5a3f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h384727841ac003948e78d64ad802502530215ce6c3b45bf3cc4d3559d5ab0768a12bbf80fcd3eac0a83a1bd44b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35f8869b6cd61cdd7174a2f3e93ab661da171447cdb985347d5160fc63ee73cb4889c64752ea99ff2ba66f835a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce893f412462299af56871f2470e8df59021000adbf1eb6dd96c302a4f5897b342925ba603d8fb775bd9165a83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118a7d02870cec801dbb8229f3d0bb5d90cc61c68a2bf3871e67088635a14e7cf62f8b8ff22734df200c54b7260;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b63e30d34685a65d06e0f4b4a8e6b09760c96dcfc47f96adca7774939567108c1b35a4f90bdace55e511ee467;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bf79b4133008b97ebce1d586cf69ac3043ca030b45aac49e0314a6bc2471a9ad532a0e9c2d6cce34562cba70c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h553a9ddb82e2d7925f925b19ee976ede523ec0221dbd1376fd61f53b96fff089773561915bd779cc138a446f62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12599524f00f1a547193b83845815a2d688cb978d1d29199c2ed9d548e372c39af68f6b5542bf30515cc9e44c9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a7fb2a3afe3e1a9b6f0db0d618b431326a520ec351e100174632f8c9abece6f5255ca71cf5790029d820c7e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad675a1f436594aba2c3f18d4aab6f132553045c5c897fe26043a80f5ad4fa066448a2197e326cd2c656ca828f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dfeb5f2e1f0ce2a3de177acf47e1c5a10d69f4f41576f61301de91bdd7e5a4327f171389354e3726a3d7a01b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11eca03c3c2a9e4747749f818d13e9d5ab3e56d47a57b1a95e8f739b5131eb395077b57e43bf6f73be682dd33d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d4856db6863ca73316f9edc998c0b6ffa15a6579b81e243ac13ddd3ea7c94ef26dbdfa259a3ce70cd777d6ef2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d61dde0924547b0fa5953803fdca9245b770d43dae7a6785a04c3190ecbc320fa214735ee2e2068e5d1a0d572;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a9af843494e75ea1f77f5f4847ddb0f94b203f14b27f11ff4a0845bc9bb4731baf6ff3625683c786291ac2ca4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a5f528330215f1bb8f1fe1da9d85681808a3727c4cbfbb3606702f153c2f9d40fc34522058e5e989c2f6b24d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bfa7d646c6bbf85baf49d24b8c30023b3d77b102e216690a33dde039baccd6f9049f20311f8ebd6e00a66849b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88b434d1663bc5960b62dce78fba5d46691697a939115f115a9ecd09d2156cbd64b4834887c6de3a0800041f22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he14e985a0139cec38443c5af687e3e0988e5684fbad87bf1e4032be5cf593f13f36e499aca85d6d2466421ca02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a08cafccac3749c80152e55dd522b25e337d5d14c396acf83c8077d76719c34a88f6a2724e7a53c39fc1cadb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2110def52c4008164f69325fa527d02d0d41dc349bd6b4e3dcc7807b7e062e18456b572d3de7fde3d0f248af0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150fa33cd551bd189ec7d03a75c1b12f0c852fb9696673d9d3bdd376271934d9dfabd09a89045fb9ef9619e7312;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1588a121cda4b24e820cd7f7877d9f4e156970d0bf273f0ad8329b4f1ad1f8543b2717edad14e804658daa70ed7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf67315e912613f0f6f2ec726a75d0f23e69d38a0678291ac2205fb582bea9ae0d85093e62afa94a143fa1a66e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea6a3fdb69a883ac419d87a97ec50336d394ea6f6f7e63f202d10f4a8c88a6ede46e9aef12f0260468eb2a697a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d45c1f17c710a0224ed3092a795402334843624548827f3f5f4fdbf85d61568422ef9a0f221ce9c96b78070d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18625fa1402ca9af01adbccc97b103ad23581accc267b6f2e90b090446f5906b8bd1108bb83afe597b3f88eb540;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb4c0d66a655eff72779cc4175b0225419c88669e31fd6e714eb871e7bce751aed61b6116e26ea0df265d9595d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6637bb00730c8655cfd6e0f4f05913b97a1b1203c103ba0f85ab47ccb12a91d7385a253e2ef02fb59241f416b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebffe3891de4176d51aed53a5d5ae63f72becf90ce5dc85647b75f5dd91d954748a50fdc89d0f4456fd1c53290;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcacc176cfc83e5bd50cfb18a62eee72412a90a22454792f8aaa646cec1ac00b3942e66b7027fe65bd8ef26d3df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c423a994ec043cc9f69d50316c10074c33b8d2ae1edd4e6c25a8f866df21c725ee9a0712d1ae0dcf04ed170a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha46aea14d87ec788cc64ada7f6642c55a8b32616de21a91da93cc3d77f390a6cf1468950a359cfd94fef89ae25;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1853eb3bab66af79b1bc1511ac3e06f78ac8d86e1bc1663a33d138b062a7ae7d3810d0a596fb2e018b877789273;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116c523e4102cd2550fd5521c49652cac0466fa7374898dfa05df8a9562e297945ae667b110bdb3078f6a3c641f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a4437ed8b70a1fd5bef2736cdc2722236efe3d149d1659d603dcb28dde9167d9e93aa8aa96ee9b89db3a9f029;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6db5a9bc127759556ffc676e91d6c497abfefbebf201c5c3f339e9c39e30262a5d5e2f2a2b8d399d181693bfc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12832cf968805a706570644d702c7adbb4459a90b407bc675da02bde59b78fe367f232b977da40b1c1f405bbf7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be8e439cf0600e35f4e45989d90264114b4df064423127ff44bc4b0ae1cd9e3e6f2afc8a9706353a29b14ff5e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d192e0da4997025a181354ea2f9f73afff76c9a3c367b77c679e5e0119f9b38a9d84deb23f221d02add828c76a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ac438944e337818ee2e7b84923e1c06674c5d3fee3a66aec2341e3c933cd159fb15cff9a6991a9e7425968881;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1280d12d186f9f5f02c2d1c44c6cb4c7f80d87278d9bf2042fcb2db673d118fd053a10efe334b9cd87cb23f0228;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1569b2e59ca24fda77057f4fc89f7c1d1ed511fbc2accad0662b3e620d8ae7050441e28a4a6897081048c1ec2c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25e94f07b9fc4c8dc793f736bf67ec7a9189fca0ea87df4e5eea82a3e07f5660deb3fe9875c334ec375b05545f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ff1bebbb612b38ac03f154ed7ca28bc19da2b7b54097bb8c18b12f2b71bc3020132de5080b975cd0d71b5b78b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dec6dc7b285ece57017de0a2ed83eb8a09ebc02fec38463fb5c541ba0bb75ac0f27a9d6084e8c7003a95130d2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57f38aca71295845c08c48c5468389a9099c60c20f09666197180281577ce73311e2bd26c5be7a959a6839befe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc1750c4d028c8a91fb58ce7bbbb78e4a5ee3ff12869274601fbce4fcf9dec0247777a6db1bfe74c25cc3f1935;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f6692edd73ee499d4e86ecdb8b9073165a55e0ddd6bef3bb8f790494c4229e373bf17bc62ff311c87cf974f8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90c2e2ebad1c54f198b02421a2d359a22b217a8a760e6aeefa6f2936498ef185ea6e61e5c2845973c02e654779;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1727588c24cc72f5dfb3034cc2d1ae06d4718f276a8229b9ad6c6372cfe3fc252013e8d787f782900cc2baea331;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fa2fb1119c08d77d6aa84c9faa0b0a17d2119d2253f6207672d248b640a8c2b2a122e0d9f017890e5cd60b404;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7fe1dcb6643334d28b550d2ccc2b27dcdcf72dd0a7b877c4af4af4155a8a0cdbd950e9478b24d0d9c1b7e85b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c914665e1a30e543101dc08ee4d9cc601198f57518ebd225adca8d8cac6d49c86955f1e7422ab0df45fb0c56b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd200f8ad126998fc8dee050306991a557e9051aecb30e1f810325d64cbfd02ae957b3f3a87381b0b03a0a998;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ad8d253e2705f590f8efe7c615feb8ada0e04edae2924fc4fb545cf6ac3cb795c563419473a6ff49739b693f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152e41aafa681ead028caa75c1b72774b26a4a86feed8e16f3852cfb246c0259066283714aed52144b13a5953fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0b7b97245fba8f6154c644015fabe8d002545c0d545972a26cd47f17e914abedf53c8fb3996f33295166ca2c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3abfa0037e07e5d4f2f1bc00e105cac45d66faa2ca317773b0e7b1718dd13f0335d59ca59cde52e2b0c1871a78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69be564dac86991904ce89502452e617c143dbfba15597fd9a128657e621cd80f81c0d62e29e0b6f2c931fbfbb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he07e402e4067190d1deb6e3a4f9b7c25e218d7882384edf626fd8e17533b20f7948e980173a5da9990e4aa6468;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fff36fc0c8423d9b4c108cbe85cfd05fea4e559fb4ac523eb25262f4d98af9ea080a6e2569a496e67bc27d2459;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198bcf68a036cc2819b09f95f4c108f8adb5b486d893b4c9a50031d6e2ed2ce197e429a170eaf0a89a0cf650274;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1030f80ff4c86ed2c354e847429f0e2cdc8ceb163c8fa7b685be7944f8ef645bc821d0b7bd0a11b736d4a67768a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h771fe2cd135e3812dc11f53bddcc832518d6620498d50df28343feaa105eea7cafe8dfbe91bc1694e227ec3bea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d312b8f3a10c3e78a907b6ef1c8a19c404b650c01fa5cb9e8090fdd3d873e2f1391dd796c478eca9fe3df8994d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h581594bb75f3d80aa4da3404f4313fa0c2c754d6d86d2a85e2b21fd46fbb98a29da8dbd6e51d4409751f3dc14b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bf3ea086346e30bdb8d8aa8d64111c12e75f0d3c4967af34ff966760afd89d83cfc8d946fd69f72b4f3eaa3dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be5aab58756aaec2f6eab0d771a27c457d288743ba2ba18846a4e93dbacc54dba35f53aa796de08a74330c1d09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c4f1997f53e3902ef0495782a68232486c46ee76fd3b4cfa7bf43bd62df05019efeddc6e65a459162bbdb2112;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd743c5f8c9a2b4eeb2d24105fa02dc5c11d7b724688ff5941332f69e2b94471fa286b1f854dc22fca21e24b40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7656226a7afb46c745eb26216cd95c797cba6d9cdacb7dacda8ad5a5f5fd45a2472b2de496d7ecd77e2fea521;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbcde478f14ade44d76f5cee2d06d334962980eca70b9464f426a54812cad8ae26369152d101661c56ce652f18;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haaf93925f6776429095a047c3f171a0f77ed2e8c196476b8b48ba210e48ac1c9449f315925b119181cd0c7ad78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haca3a9fa56625ca158ac2015de5ef81f0ab9a31d11188e18bdc932115559aa8d42eed348f525ade69439f766c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68993d0c83e1f16dbfe8e6c2b0f2b2a01ea4da31694f1e70f2eef4f100dd974ce7b84501651b63417d56bf8f00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198b6d5f90cc996dd2e56c37a1401ed91581fe5ac5e4a2f2c113ab2ae4b390bf58c2408e2b14c7126212d8fb750;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha9f908ef46426c17406d468c8990232310c7f904fbe224379ffaa32764870f40a12b9f7e74b790242952fe0996;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ee068fd16d824740fbeadf5a820ddc7febecc88609bd72c01e1120b9e708b7dcc5d58b84b03731ca3e3bf0ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7a079d2822b1e1ea1c076d184c144fe00bb349ce394b0b6debe6b205e2a7c739bc9302b6e4844ad45523a98dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afcda89d027526d645ea776ea511a31d85556cad433eb76ef91292ec0d77d6e4f80b9432cb78fcc9c37c1876da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fee5536d18dea8abbe0fdc3585116c459b447a2e21504d3ce6131156d22a2a75017a2f77824af7e74f408f8d82;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c532fa49f5cb1f3f124c7caccdc3c8f191e498d09cc8feb5ebdf5a68323933ca984baee1287d559ef8e5eadcab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadf95d885aca03bea68a99984e4f377cfb38f85d89b07790330c146bda4bdffa7eda6fa585244e77c8764dbc05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e013a628387c585a0fac704a4092d1992d2bca2d12344f6dd185dfa29e062fdc4cb4e0f8db24a2654ea8c65af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd11cffcf81dba2c818f5cfbd26289b02c806ea7df1fa6c47ce9dd7ae9e2ade507f49bc8cb2133e14453f194030;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f76a0d40824a6342479a81a520d319643b078564433fdf83523e45f36cfbb618472e8771b5cf165c96a4211f1f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f6616c0f303379c189967ca7a4553720483ea8e1c4630cef8007c8faa3a81df6e856b6666462b6c2616cfa6aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92caa4c90f79affca467f694630ce3ab2777271186012b35f54f24fa6956799022cf54958a591d3669029fffb1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h638b4e2a7f9a99766b1b4c49c4850f6be2d657f50d1719303dc367b54560cbf94f0a476b22ae35af97bd18ee4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b27c543d1fca08899d79201ced0343b619c0d4ae6cface1a31b5ffb9efab37ae9d737663b9bdfa67f9d51c227;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7164eebb3bd5ab14c6c0bc283aa7efef442b5aa11710fbf58f23c8bb2e932122724ee31161045d385599aaa25;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195cb413335369eecfc94919b0c7f6c23be85c24abe03b1e2696b6cc99ed1098a21c7817d20df043e16c6098a0c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107c857c46d7071e5b82782099a355d3d9b0b532e62321a2625769e6ab09c00094864767a553e2c1f4f47442d1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19004d82c225276c0dd9b5cace8cf104071ee9a6914c80e45675fd8fc0764c821bbac04775629349af0d3bf55ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163341b3c060cb3aa4cf2936aa64f4fce9fc75362a02fbb7beea0799fa0dee18e2ad72958d838cb75cb25103e6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11dc9567fbe6ad80885c303ccadac3deff618abd54f978b1511690e6f56089e483271306bada6913f77263f6623;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167dd69ec508773011a5df8e90a4bcf23f053eb8f6686e99c6ef59b6da438cf295a02e0cc073edc3e73917386d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbbc2054dc5eab7c0be43f02ce9bd88f9e676090d147bb57ceee0c09f440d7e2e113632788da787f2e095f654b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a205664561d76b6353b85b3bebbe521c3e28603bd8b561fa07e3490ed000f7b01f2cdd943b1d20fc25e65e309;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a1e42cc77f641746f4a8464a1efe2d4f1cefb0219f536282be2b9124d152c755df4739560d4d44c3e6a67b9c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf22d0deadd430a1268ea686f529c917e05cdcd793fe1e212ee80520034cd422ebea35701f254bc79bc60645fec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17fa1708bf9c43e41b65d488198a098edfcf8209a459ae7b94d573f2d5ab149cb802ce67d1b077e9ddeda0d0129;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b6f200bd210718b366fbf5c2d3fea03ce9b0fa1ac0186b7d9809ee485ef6647da1e146c69260a1b8101272a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9151d0734b57f247e24066c6d5886b5e64dfda65e3f976fe4d1087a71114f31a355c29e4034853bbe6bfb300f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd368a0f0680e0d445a190adb0a969bf15a788d04a46a5e40d0c52de184fbf30252e301d2c788edcc2c7307e2f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he11711ce72ea083ccceaa9d7b6d1c9c232ce1eb0bef9e85845f6f3699bf86b1397d59d2a66f5d32dd80a9ae778;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a909e36f5e0ffdfcfa03abb2a0dab0037dcff7d23c94f1df8f94b4dcd345a2c61aaf3b0c539f6ae7601b0c65f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d7369535411170c978a8723af0740161ba3295dd61fbe4d584dd9cf61bb57af0b20f1c59bdb3e7c7675044298;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h158ec1612f29802c0719ea2d165c562e0777aebb3a1d06f047cd126fe0e71683407312b56dc36d8ac9eb10b6f37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0517961cd67ff6b6bb22755907799caf27d7f2f31e4af2e215db0b17960b29f7772fe52e488872881676e8402;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ded95f8830f14841379a7032a89eb9e91d20850f641375134474f1b5302acdd7dc093ce6f39793f324e3c10cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab18327eda1adbce57ebdfa232f65128f4aac6f9a80a7b8712ccb59534d00fa686caa67e6767b7c5a8a8e82147;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5f2e012b922bb8be3f0796063fca8e27ef2c1702f216be1f59bce011036bea4059c65743e0396c83b45ed6f5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186bc6897f54484fb0b5525cec16f2d0ef1afe758f4925919d9f74a8e6bb8b6e500d6e8440b025d5550c1dc1ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188f115a23f7f930913beee3b610f2b70180f78b217d5c87b3dffd51d4e81c2e1ac8396acf1dfef47b49c417c66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ec32ddf1d476bc7fd9a1f057429e990126141d06a97a30f67c48481827734c952642ba9a7ec0f6088971120cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcab3b8a18237b55b33ebf30db3ec4e0c7c95a267112755a3e6a4528604dda40d891235457aabd21c7754a2f9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e2b8cd20c112f1729630e9938bd5e71f1755e33bcb9ab6e683b40aa95dbfda2cc00a77c352bd96eb4b419c5fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104e621e48b859324a900a6b9d1a7d4cb73536d31b4b956835cec01b05f695bc3ca2afce0ac81555c2dc067deac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173cffbb96858d0ac5aef135ad016ffc2b6576836dad35ab2d46b1ebb5d5dccbdbba50f70f76df46f4f5cd8b64d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161d8926298876be91bebc896e705d221ae278772dfd7083d45576e751ec81796b9f9a31d294ec3da3355553af0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f3d5148240aea2a614275d04e0ecc177689288faff2d2f539ec8644e4fdda7bb7660e155bae7c5dfe420ec5c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab10930d75dc6f1ec7ebe9da7f12c155c8cae053f786ac70de95ac559c6c71c10f72ad255f01bb121c3e447ac9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33ba7d7e99d58903b6345032a1ae88b2485049bc10264db19c5dc2b01438682a12e55c1ed03d15d8b33f222694;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2c0af7c7057bd57846c494bf93d086112e8881ad9ddc951ecd300aacf7c5cfa56e4b366849dc87bf023bdd72c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca88c1365c7456629df58783a0d694d5d436a44e25f60e6cdc5e0285bc3b91c3a4915d42e49155914b300306fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fda1f3f5e3bea3d234d86cea094bb722420ce69881c89eac61b0a408f25abf819090df133f6a5472ca57f77b4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2017776b2ca9b97a5ac3839674815bbb5d24a22a407ea2168c3a4a6384aa5387f4267ea07f44cd21a44cb2445b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb56afc5de610826c9d708ce83de9124260acd2fa16f0b157553d1e983d7c6f76293748f9bd849da968a7ab220;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h458d4941701af6054c26e61427ffc3beba1fb235c2b22a38594190a26ee559b7bdf152a478948fb16985ebccd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ec79c0d2459c86c7a9aef98bc464a25ae50ec392b04becc88201c265f26f8f8d5f2aba2a1c4b1b0df28e849ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29efd4d52f45019bd8a883cd17578550d7ad4a592da37f903c1d7bfc5744d74775b2ca0b70f13790da70c4e5a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d2e76ebd2815ccbaacfd21ed3a3cdf562e5b7a17a805148a5be7462b6349402bfa0cc97ecdded4e9b193e252e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb13f0c0d956de4ef68a3287b801a1a8810d7ae3e858ed9b4799cb2c81a435d8e00fd3a86212b8e1ec64f20650;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115c182a4e6b5c49c3114e8002fbc0b9d4a50cdc1045546217eed051b44779aac6f93e4f5941d04aef068173fb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he327cb4c268b34770940e6ff02ef98813319f408bbf7c25eddfb27be50cf1c94cf8c2163b11e0bdf4a1104cd48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h789722b6de46db3995d059b48545208182e14ab68305a9e36ff6ff41df85fa55bc9a9d1fa440aad1b108ce0ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2c31f70de53a76641a7333965a44ba40350d55054965630ee98993f362903a5aa56e3b7dfedb09465a9e44b33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h162c51bebf23857d6bd3ae1968029ac9417f56b73b28f04f13f55ff097edc57b9e96c0d1d416355bdd1a0693ed9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1072b4a5eef370a4604138e5a00bca2b98e3a9dcd7c0a635c267e4014ead8569452ebe02c7bbae2cd47f3e6a93f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67d680bd2f9811225c01210bfbef82758235f67eb5485713dbd672914c77c1382f782d3667905d5f4b559e07be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ebaa30dfa8cf1b14ed0e013c3816b1ba263edb2930ce60be38b76d55ce01450d44cfeb7582a174dabf6321dda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9259d9b5bf3388c2dcc701d5245848a07c98ffb13d213ecdfcfc9f9150d91b8cc8acd20b941caa0de8b925a7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd2edee8da181473730a9d55dcc5a1c9a0548585cfab8807f7aa8aee1ef7beed079a18c1d963ea10c51cc8d707;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb4067d231b240cb38c77df322e3166982f0254b424306ce354ee9ea5cb86b553f40b85c865ea15eee82db92a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134b2ff81381b9582798c5c4beaa8a992a22db2d7fec37c3224fd5a0196dd6e596ddcc236979a06317fb7d6af52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d88bb44919926cb6954f88956af1778af76156b1a9025e61a01026c1b8da08dbf96b0a9f3f70358ac3bb0325c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfcd9e7fd483f03592c426dcb55adc40b5c9f2ed595dc0461ec53d52fd67daf05b6232a7ab8643a44e8ab606d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9433f309ea716b613baa2bb49c0a2a71fd9ecc1447da3c5e8b310a857d0603e8ad2b5556d2b470942ff492ee8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c09298afb78b00494feb56bbd17ddede6f15cfbf869df47c2dfae2c657487a9ae6683a2005c63704f4e2068a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde04de6c4a1d9bdac8d11fd363bc63f57c9dde2fd201723db4475c037e9bc9e606b123c2af449863f40b1387de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcbd1ee900098521d658d8b774c0e21888e5420f3e802f1a772e129291a680fe7bd5429e3fb517fc90c3c9036c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dee3fee2558702cc5884ee6bfa28b5193df179c0b65e783ca41b1ea00c61b98bbe7f9b68e2c96766c00d633d57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h456a16bd500ec84c3852b90e2d1cf39ec139fd70ebe1fd82808f1735b6a0d686311efab0da24fce84e6cb886a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16221995842e8ae73ff93cea91463631d1c85bb785f59f78d85ce001181a4563597b98595bc736af1155bde3a62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed16e70d9fb4ed58f228829e1a5ca60b405b36011e43e584e8fcfdd69bf602b1b120d2b6b561859c5f7b211035;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e664ffb45b0d711e44982ac96f44c126c56c94d6c21bb9656baba30c916a2793786f023811df30a8ecd256f4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h73bbf193c6c14d431b32e215e5a40742daed16ac24630dd28c44503de9f100ab87f0739c159b0fc81ccda98b38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93b63307a045ae2750ebe5fda8c0dc03edc8701329f8577ee1dbad5889dea2482d32caa0b90350aa8294708f9a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1caa4ba999872e56b11987c23916ad3893b014debc4bc46cdc44b170935751dfd2c8ff0c4db6950e16fe6c4d234;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbab4bde43166c67ae62bc3ce4ce9e451ec77d5a8680cfaf09e358e46e5acf56d9a0779e690a9cb4a15e78f38a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1508e65bf1c8a6a7b4870527433155edf6e7515a8defc90a520fdaf74067e98999fa89f25a6b34a3af604cb9f8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15546f1e64b2c8be58916a12daa375efaf8a1d686b4a458e8518373a0d2a056bc4766a5b8ee11e2de19bd87427d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195ff7979a54d36a040b58b3b12b0e6163ae9432f0de81acded942d520a87034dbb52717a3ebc29b055fd699bc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h113a9406524d87d07051b06b99e04fc6bfa4971efdb34e19fa5d893b632787275c315629377dd2a3f1322f5b99a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6b07783e10867013250c57baf1d56e3ee315c76957851a51947152277132f6b80173f89f58eeebff2af4dac3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a4fa84c02f6ecf6e314c9d89e8a2a73bb46c7f4e56eb37815db1bae033d45f078e78b6a7a90912472ebb28481;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bbe080f45aa8a1df6b04e679baacf7c6f6d931d1f34710ba7523fea925df2e2c7725d44e49a307c1db45575158;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121734d1b3887afd50b40ee387815225374f1473cd29346b86369b3e53a146fd194109469e7134daa2b61d44ca6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f39827e33d82a6df602e2074a4105ee258c19b728d7811ab2229ae817e328aec3e604cded97656f041b34e562a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30c0edd9925e3b5888917541a49648f7531a3a53c47076f62f7e923837766676177842ac7b101f9934620df090;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124829bea90e43803f7989e5b69462bf151498329d836407eb8a9d4b12e9cb074b3f865ccf9ce49df5ca18b0416;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f203c97421aafa8e5d8d24fd84d5b7531da427d1d6ee1ebc511488b6709cc8157fe599f656969e84935db9ca0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ecd84df7b5be8f3bece82bd889ce0b96e86a3597133247e17d8ac940bc6efd3addcc4732acb081bd5e103476e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e333ddaf0aaffcc15902edcf4c78ef98310a09f0ac53be457020082adf5d57fb1c00dc4fe22c761f8a99163a4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19aa15d61f6f237ed4e3073ba518a38274353768a2a433de05aee751abd838a74a92b93bc4170b7b1f8439dc01e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1705e2d09c82cd53455e16829bdcc0869bc2c002233617d71a0a923c85898525603e7703e36546363a04076f711;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d16b0f3408f6c941c423f6d86a58c4760b890e2bf660e51efd91d1af9bd8de88313d9d25fd542684fb41ee607;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cb7ad0f019610f7ffa63ddd3a476c8aeae9eb5d3fd6b08fd15a7d9b6ee3f1e8a283f2b58db8602280e03ef7c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10639a9ac91703a4a2eb3952e3e974b39d8aa6c32c21ce19ccb06afb2030c4dc914c714357f2aef56c166c18677;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9458c876afad37f8c62d90e72954e3077cedb4f694889f2c7b296609e58ee9306beb9dbc6aebaf769ecfebc92d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1adb8a66276b9190fe729850d69abaf1b66098969f61830ba262f6b58573f80fecf65dc83b214fe5eda918fe8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd80e49890e71105adf6f62a48d2a93d5a922faf8f054b3e47a2987598bafb983c2e1f1617166e79f5f3c33ede8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha95649ba961c87cbba455bf690bedd347ea6e8444b42dc30452e1e8b081b5c9da7b6f78ed3d287a3d239f20d2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd897b4840e90be2f9cfb363fccd5ec410c0747af0cfa05ed01211bc271771d814c08e70cc965f19d335263de6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1292412c51c2eafddce9c4741923eb6974488b5b6b8a7cdf1cf407c3957a2ea2cbf31024521dc6256360b08f0d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17522e3f64158d8fc947b6816e85c3b4f117afdf5d8922cab7f3230c069a71371e1e3227f4a3dd4e32c7eb14b90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3f883692c124548e4937a6f0724df0d9082f5607a25c2612b8e1f6fa25657ce39d4d62e934797bc3bf1041cc4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a2f609c4da8e3f4d7141717e0fcdc0c57cda0fa46f67ef0ea8b87d6623dbb26b6137f6dac7fbecd62418e0921;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ca87c925d0b9368e1b8735517a10cf6fa06cd2b87057862aad9884e4d9107821227ce063ebd2a5fce444fee58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f4f1960e74861d184c7f0f29f7f17d3d313fc1c590b98285768d0ae58f4c9d8f53fdf49928540a1ca0082ee48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89fe0bdb53006c3359c4d52cce4c9291f52fcb94ac229415f5e027c6df1498fea5927bbf85fe7ec05328ebafae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1378e4b454f19110e140b6186e7e43307d56aa53c3b3bfbd03d606da8829e184c0e7f237775d93926cda7466de7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9e6dec1ead2dc7af3264a54fb3296f6312867f7571cc6fbb57521c0f3c8def308bab34b43fcfa6b1e57b841aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca9f617198ae03f0d9385b0ce1d74a1ebc01a1503d18a417f7dbeffc3c0bbf0d537dd3e3d0d3af58ccc7fa85dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19016b63dfc778810f162382b6ddb04da99c460d2dcc71b1edd6f5f58e16e61ea96b78e09e2d404a6966553a858;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b9907a5171e0a44a11112c75d9d0d79c019730dc8be0f01edea2c3193da7123c08eaebf5ee75a30d5b548b1ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0f37ecf42876c3ac3724dc2b28a6d43c7cdd70b4f6e213a3cdffa85163a5206e42078059a3d5b26a66b60e37a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181bff3e66814743250eade9fa4475c1f4950b42e7a73ea660591d25015c8b00bdc163e192d715b67c3318e4f9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99ae0338ed73db078ffebe6cf0f0078ddccd7fff0129375d89bf4db8516dfef9cfad093fed31a75408f8ccfc4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60ad46c582b163b72096812d44039d8fe3586f6744031001e56236b47b2e3c4fd0c1fb4994c3dfee9a5fa7cea4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bbd1f81bf52faf0a419567885b2c032e37dab16a66a4ea30d9bab9947848da5dd090c5e2101fac4aaab25bd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1419b4d4bcc0bcd2ea8ad053f0b0e49e4d43ffc8cbacf8707f5402627f7041df6e593429663c0141d13be65133;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he20b3d816dcd60f2412c43f5ab14151b67b32448bb97dd7e00d89b3143051be8cfca0578cb93054ab1d1ea55b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8d76c1d6fc420a6e6bff70cffffb5fc3d875195c467d3c9db6a391c602613d415ac416da2b73952a7b7d75a94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8fe2b027bbbfd942ff8c05d48f3dbd4676977629562d51a5b762ff15fa942ed4e2d2dcb5b74933392e3e4023d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f6a7fa6567fdfb94f2dcf0b167e353d299412b1520c9d7e679c875e4e09a96001b374fd60bbb88803c5cc1485;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h936c3340268eca969a3a87b95830d55e3c2e4bf19dc2c0c8051e8d1d22d6e2db610aa213bee973100651ca98e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c079f26e0272e35d7da1727edcec121beed63c7edb0238de2248496d770dd15681a88316c8537fb8a1689a662;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2a55ef90957082385a162844f07ee2f0bcd84896f65f44afd1bbaf0085bd1c9ff4b688566d5f18310eb04be83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef60269a38aabadce3c91631739d8f5cb8d2b97db90a5156dcda5ee6587cfd3752aac9dac5329590d21f9143a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150e80acce0f5dd9186d20071d33e5d5d29ec659b772e77afcfd129064169596b00a37f21e10de7fac490c88dbe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196a52ce643afbc23a6312ad2ed366d0b9e4a4dc934922c1c77ef4f1ea44f7bebfff71c4551c2d48ce97ced054b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1591a78e81be619f71f82d51c0e273d63d9d72c6a986f7d9f6ab425c254d2229919970a20d0750debc4219311b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b0d06decf1cb4c51fff92e639caf4601396acb8a125c5d98b096b07d139b587d1062c8d855c4ee0bba325f4cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee876bc7b17d561eb81377f9920e1c6ebf2dddc78593b608626056560c8c5713cc52955164dbe7036171efcce7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae57d3c6b0220a4eaff458fc2c2f18fcb9b66fa5cabf8a038b4fa08233b29cd4cc93771e3ffd376f50c9b928bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf17ac839b4cf975a19bcab1a760aa575b1d96413f010320ec6de35f075477ced23844b191c147430d53f1af737;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1270f5e8b25d87da589d6537afcce5b1389343b42311095fb019cda205fa4780504385ea8c7c90278604c19a339;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7d9e4a23b6e71058a49c7d21eca26b2024c4b30832179ee6e602ec648bc07889a7a7f3badd0692f5af4ef5615;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c5ee6968aeee9dcdaf52e574bb256b303b24e9df39874fd58197fcdeec5aa2d4fa9adbe04d9d4a9ea5d9ba731;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc06b77532fc8079d4bfc48b018d21b6f2d84b8aaa3fede43a421c65e8bc73d4a5e93c7c6bb1185f3d4756f43c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe517f87330b33865a80ca1bd3a09c546554077196f891675907fdc7665067dbe791a8fc28bb41c681bcacceb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee76bd946d918a968a45757a56dbecfdfd565a8f2885d8c56f7ab4129d2c374764df3167ed8f7840ce9cfdea2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c6b42b2d6bd17b754981ab12f5f1d19adb39be33c122e6cf3f8604fc267a44d453855b77bf0e3128e59ea16c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf42f81baeb652c609de3d41e0237abcc8e5ec1d2483ef23b97cddcfdc57cf05db46a9251b3a3713119a3ff377b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148637a9c0d840c27e0376dc83527e28f786a909d46fc9b151dc532fe301d6883fc0012375f1b705938c06b08c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74764915c1a1f5fb2bfbea18ac5866c2c3acaaa98309513cfe6170a861bd0ffd8cbe1898dc19390d2f66e29b1f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h700888e3cd7edca4310541c8eb1acd1ff15c9582077c81ee0051f5f03ac66ddeb599f2391753b6b939aa5eeffc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f76a10b8db22c6fb6d3c0fbe1b8fec071bdbc969d2543c014ae6d5b821a72def7dfb896573030738aa52231ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a30f741d02efe8929c052ab87041a1e3c2d3bf695fc46267e6443cf205d75a4d0d62fa6477282b77ad17c38de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a12c2b1110f1fa9b85b93b781fb4328da348450ebce40f24f65708b905aae126c3a6373e98d1049d04c241560;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f00f127231e1f986c88c4ef67c5fa620d93bc9c0398867a48f2ec608d673577e52edd2ee8c0a86104761a378d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134b5324f9d4cbcdc98d4eefde16057e1b9c498d3fffe530e2229e22a80179b48aca99a4d1460b81ea314a6ae55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c42f7a817fd1c7fb8449f9e671c8696b9fba77b2d5c254100039460fdb8c24185e8ac9fd07ffb63ee5a98c9f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9a05ed5134ee9aa2493d851c3aab2c61b8186622377038ef0bba7bbea1f4f53aa91d00b313ead12816d07f9fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4529196f34bdacece2a9b2735dc40a4b5e30efa6f262438f474930aa7b33ef13349a661f5cc01a32eb6535af5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f385ea2dd0df337f22622338f5b3d18ff82bf9f2f0f0eed34be129f37480e7d8134301c5a2b7516ba1d68107d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef454ba666b825242656973480668d9e630765fa331ae0149e4e0ba049975129d25e23282b72b4592b315b9f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1696067f781ea9bc8e9e3cf1b8fe8cc5c529fdf5e7de674ccf830a0c689ee59724022f3fcc3871c900ea7365eaf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba895bbdf8677bbf95a4dbb2ed66d237bf6cfa18a9b8d25b78264ea76bc3cade5b9e6f2df1ba42d9ca85ff22d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6fd808c4651b46e2da2203ae62ed49bad78e3e438d1073866641c79a168a229e062ed35bd10e27ff8865e18092;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd1f5c2b0e304f088f5ddc02bfe2662d56a470edec74cc0655e5fec5524abb2205db112ee78eed692fac9c9218;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2292eb5d1074678267a157d1e1e68dc727bb160cf82813f91d561290ee3c0e89bc23479eaa6bbcdda19dd4a639;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172153b361ee5e4675bb2af762472dad5aa4af1b34a2380a67984995513c9c3434c44b6bb69acb3e1c5a4776dea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94a36750fcdf1ad92cc5d7f3b86e82cca9bd21ca78885340279b32d8a3c1982ea29b2927a2ba0a0cc9d5fd01f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e56021598bc1ecb192982b68bcd6bb732aa3115b52e1745f5b8c05d9e357dbed2baa702584b24ef0eae43b21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f51662ad8fd674ef444308418da1e72a06656e44faaf01303954702f402a71a704f178e5ea494e27ae284f4cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4213c990667772271679d831f83d4a2168246cee48d3b2b1c768bafe406e010811e4b8d9037baacb1000a2450;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1768bdee7417e28b71b0c80a8320ee9abef7c7e5ba83c68c5006b805741f717d0b3cce91ab575fd7ff33b1c1b50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1859d4fb95403ba2a2da4e9cdd3a0d2bd92f898539598a4bfc8fb48502b971ddd0f170f238e38515286faafaeaa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb68fe267bffff30ea3ab1437ac9be2fa17e4dbbd4f0b75c0751441c3b0df476ba28d396691bea273cccd8707d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108e162e274adfac22fb3560e448893f11d4e9a556fdabde31d99c2de137bd42cf9a6a8f0a22fb547632748fea5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37d5e05d3bb3dd86f893f0425c8e832faaa93cafd57a69024f2ea7e42842fcdc49ec33bd41fae914b30afa9b9e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b2d8171395a8005c7c6915f3ff09432553713c94f8922e598d6e17902ac2952f0473b8718558d6febe15082f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1292c59b9550700cffd8449bb03707a8b0e31728f95a4c9b0c7b647f9db874b60700b51bae468c2e5fce7fc8b82;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173b2aae8ed3ae7903d3bc1bd77cf5d7a7a21ada1750125313bd9f08bd2c1f175e6a8517b34b5468a2d9785a6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dbc6282690c92640211c5e8d846fccd2326db0d2f89c5c3f754d6fa5ed6de07651d7efb1abb16826ea0706608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf38e6ac185c2a96c8d1114ff5be8d12349069a537cbd0f7600cf80e1a94fcc82fbcc530252d92efccab83ab3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187c0adb1a257efd83051a53f2a1038fdb6ad00f1c7ee73ac37a3d38da191d97e4d319f14ac6648daf03e83682f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c89566b13bd79498d7fd1a99e2785a5f3ae81a840fbfa0c65839e730b8dcd1b2b80a7870ae9ff150ce7aa9c91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121f276f7a200c6868af58a3efe71d262df3a2b5d11e8a2bba0ceb155e286aadd2cce0ab364648a53ed1d8e1144;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23bf12cc164051733fb42c413a1de0fca18a9ed383a6cbeb8858526bfaf31dc631707b045b55fb808c27bb21aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5fc07a368e4eb10c84f7f5625278c5e44385ecffd378467b9476f6e20597ca3084172c001d83c85d555e17a29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd7b9dbfedc99de3a923e97db54b027443f56fcd4d218794ce3b614ae627aea2b6c59626287df1b260b220019;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7e8f86727282ab1fb29595fc22ef31fdc07b64b562e0ff09eb6124f129a4bd263a16b39e6a4200178b53d5046;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17836003e92fa1c237269821bcec2b96e849c6daaeeffba27427c572ac12463891d4d6232f7a280e619e61a6542;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1917d1b78ffdce9d95f5bb512f280fa52f18919024197370a656ccc6fbff954fac38e5dd0f388e84576b9edff86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d48ac879d8da1ef379109a6e5c3b7a3291bcaab028a5ac2c5fd7f49421552d4ae272da652523e813146d718491;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7c580cbbe24478148f20ca4f718eb6f37f1c3a073058b60d7581102d98193e373dd5e26e93f6f9ca7dc6399b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a91290c8eed8b80bacd19749276b3082becdeba13e8488278d5db8ce93261de1712a8bc07edf0e9eddf969de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51a501c6007c31a107a05b89dbb4445188f2216be23413e622b3563ee6e76fe38656f2d9fbb2f387dca0cbf80c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1d1b66e0be8dcab17e89ad63216a0473aa9d383b84f45be3bb8694c557bec8966ead410e528998ab0fc1da331;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1958aacc967eeb9657317de2ab6c8f2e3b8c37e441e64edb50df586cb503604642db737bd9a573446dfc997b4e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0713d3a78171c7d5489ce1f0f2d40340fe0d518cfc3eedca0176d3ba1cf74010acc4f98d43c57d2d813f42c88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8db2b9ae9f0b1bfc5fd4a5a2196b457ea87a6cfb1c4561a2015dae79f8dfb83703b0bf7a82a7221517057cb4d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5462e4b67baacb2c9075436b71a04ad4aad1517dd065294d4d8a5ab9ec51f940a06704a90ce5d670386599e30e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa6196b1a2a80ae2a1e969d36e141f6e2b04c1419b5f796de44545e2b876955689c581ba567e8b9f6c7999e856;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce4d2072c47980152555a574c410be9255c0595e8987dcb0aff0effa4f53f1f8a7cb92e739c3cc315ff20c66cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160dc9ebaa6738cc3992084c348ad6f2691d643bc83aae3b3190345eca4b6a34643435870b80ddabba65c9fe98d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60f8c28c8ed663ba57a64475e72aee4ec937113e7fe7235f8adafe1aefdfe924351c1ef41b696464c16c16b769;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee6f62ef5c26d19f762cbee94032a11f1ca2a03569fd8f0d1a14fd864e3722ee07a0c6574faab5c25505b432fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd9b14659f0dd096889f31d5e6c125fb9dcdebd79fdf0e035e71cea9161da1ae4dba2b1cd4327a9e00483eaf54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce82e5591e8eb5d93a459fdd2f283c931d1915e19058696c90b26936c59027f967eed13cfed1be7b51de95d220;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d0540c150142c5ea2ba6774fa5f9fbd028be94f8e1a366110131fc0c08fbd078fe4fe1780d4b4bee78d138b64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6758016e7eb886cab6f23ce713c06fdb1a602efdacd02bba193aafc31059e35b90c7e726277f205a98b7e3eeac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8004d7e6211f60c4306434ee692b203ab3d6a843254b28a130f1c9e6e0abb85682269aad6ce1ff9989fe30f876;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7f20a4f0dfbf845a8b5f422b2240260b2c0f199195bd04ce97e834842239e424d159f41d3b8fc17a0835bcf67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193e8fb9a3e0e6f081adb4b9e3d5e63424f640360dd1f5759bab07f74d01ad510082755e7b38ad11324c2ae4b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac8e92ff460dadc91426a94161d1f9eb28d68c3f532cc1e8f861dfab49e8e0486f656baa8b1ca341b554e40d31;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8bb2ea8de0ae9c9a308d6c60f07841d14c2fbd8c63fc1227233f87c80060b8e0dab9b403eb9291141397aa35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1630450274f7af67534af6efd6b7520e2dbb3c0e80fc77379ac6dc3624fe64e8e521ece6af2546b2e6e84fcb96a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13678a84028a33971c340ec908dc09d187f7412b528f168c8feae2663cf0a463b355ff69a9dcc1cd1091c6496d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66d6bfacbdcc1d4a61fa9ee3db0d092199c60698f8ebfe641514a7199b3aa75ae8610bfcbec2071db24677b937;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e676af0adf268597047ff332c487378bfe2dfa5f84694b5452a83789932c5c067a2dadba62d97822ce90a070a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d266a0a6753147a5fbe6da2da6db9b3b48bd4eca066a47db32f050011670ccd566908f3f1cb0a605665de4fed5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35fa1173a521a716230f7a4612661048ac408661ce8b38007bd4ffd0a3f57da2a094b38bdbc428fe5da982cff2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4815c7633653e4023e706f68d38a4180a1e0d05cf0489ea8014eac1f6c3ccf51eb8b11e314b04d9e5f1a95e362;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bf2114d4f42b2ac58909d7e4300ad04180ce8e75695c88c93a79dd29dbbeb7ac27414b2a9694a8e14a38f89df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8cac66bf0aad49c4e40d6b50dc216cc884fd59ee87961664134f6630ba2eaf4b89f2d22003c09a15a3e6016a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd257c638d6453b4619f02d44e3075a07ae3150cc2c43ecff3daefac6d8340917da2f38023973f562b0dd00e65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f393f78143a29bc9875514fd0e6cff0baa699069b458ecce4cee1828f3a34c59e85a768bd5518a68b8698d09fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb909d88ae3eb0fafeb6403df2b6786543130cda3bd3e04ce53490a3e207b10e50a8be497a36ac5a2ddfc9df254;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1953ef8d859e16b2cc03f56db8c0d2d8e56767b37af31d0bfc05f31826177933536be4d9d0b4bd95cd0a0ed89a4;
        #1
        $finish();
    end
endmodule
