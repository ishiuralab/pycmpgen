module testbench();
    reg [18:0] src0;
    reg [18:0] src1;
    reg [18:0] src2;
    reg [18:0] src3;
    reg [18:0] src4;
    reg [18:0] src5;
    reg [18:0] src6;
    reg [18:0] src7;
    reg [18:0] src8;
    reg [18:0] src9;
    reg [18:0] src10;
    reg [18:0] src11;
    reg [18:0] src12;
    reg [18:0] src13;
    reg [18:0] src14;
    reg [18:0] src15;
    reg [18:0] src16;
    reg [18:0] src17;
    reg [18:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1862303a009adaf4603aaeedbbe45638de869f45076ee38e47e9780d565fbdf754552e22fa2ec45484c80722923;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec13c89fce0f2ae73dfd0c2d033e16873f90b70d6f47ec953219aeb3f258480d6c9f82f2b5d3633287dd7d7ee0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19715960d2ca6569a849c2051846e3c102ea88dfccde7373176fe23712c54e340f9b9924beafcc4b5b991af7c11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdaa1fde476f35a2fdca60afa50c5d4812405261f76ff21399b35fa5575f90a23bfba3f12904237fd1670db1315;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c0cbaa4478570873d699aa6666b3bd737f5b8de56000fdace6328bc13e2af1c2135eb2f5acaf5392ebf231277;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcead26cd0fa0676a10b221e524c59acd8858e78737855ad1b2e72d473074ed09ff5930dcdd00b4f7790ebc11a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa1edfa1d2ba3adaa3e6ea109b3b4b0ab54e1b15db9f3ce5d82c9313ed3570ca712cfead3e1345d46af393301d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5dcaaa61a8016dc79ed7092297e89b9217b58170661d2f2d495dbedb7827587f9befe5bc4d217d65c0b9ff73f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba852b4354fa0cd4b59a67eed51a9e63dabf8295e3ab61c11d40317e0b9293e8b042b880dc1f8b0763c085973c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105791f629be3ea271dcff747a9958bb4c6d755fe06833b39bc038791e2aad9dd2d123958cb0fb66b14bdf92b0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4940a1685a174bfffee6c0bb2a0c5bc86ffa939beff2f4c55e2e362899c87b1cc2a4fe3f6d283b803f977a0b66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28eac445cefb7344146b741ec3309d32379ec8d6fe88b4dacb201c7b8a800d71ddaa7ccee2da949103e6a91a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b80036f18ea0b396812a0a23871559be6ecd214cbfec7751d7f67f0ad02da184fda712b689e4f0de932fec77bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d237ffec0f77f84d9bd240bf283db976317c142d4a9a67f94e192340dcae47d5d2607c86126c084059969ad459;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e057e8d31f63ee5034d932e40aa073f7437437dee05e8781d31aea9d84cd659b110b299b60d66327d40799cbc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha9e9c7abb2591ae5d23aa3245d60d2bfd1e404bcec93d032a3aa216b5ae19e2d5fe04fc62a50d9ca94c16c7f9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44f31adfe48569dd57e9bde773362c100c805193cd8ddd9f8e499adac3725e8de1004c56d1e51a1d9e171da11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b6c8bd918c359217f37485c3ae8b9f29c7bc958416cc4f78be228457e45ba5edcfb27dfd9d6329cba0c6f27bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7b4c58d02c5ff1815687166fac9d91a3cfeb9896066edfc67ce8021f3644f7c75762b1625eb941e756c6ccdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c64c2e8594455154050f7e9e5f48d88aeb7bdef92feea542961fbc4df62a979d37154363a119e9212b238970d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc71ed098fb5ce9dc4b89b65ab6c054fd48f0640a72d6e502fd4d5b973fbfbbee78f6bd35bddb886c576568ecdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbb232719fddb18eb4afcd2acb18ce4fddec240ac8de442e42f16694a28a2d2910ec1b2859019cbaa15c39a8c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10dd97c5466850895baf0c40f13ae71e4f6a95678f555f3c6376f68f419e05e7f8b965efe381de3a93651a9d7fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfa60ae191058fa55206eabf2e68912bac43a5f10097367b1c4b03d40ddd26b65751ba99a5eef57d225803e689;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3e88ebf1245429ca058324c2b626bc9416f4d5be77dc23319ab5cd1162d6f86e12005aa683fa1f2c221fb7847;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193483a496eee47c5e97a6494d6e0329ed576679045906a14b3849c86ba8032a5d012ec6f9c376dadad2ab8ba9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1248c045cab12c6ab3d1b9437fe34ee6d22ec8949b3258da4c97f2b1f1ba64aa592558588c895bb19729cfc398e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd337ee2135af46b84c91b81da7a460182d98eab2754fc839a8bd205206d72fe1339bcd314894f26b5df2c954f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6132aae543d33b1602e7458542be951417c2d9fde022d6d1fb73661ca11512cd932b5644476f58faf7b45ae1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6be7270201e340f0d7cd7ee6912c87d139e067aaa846e1e4f45e01e2c352cc16a2ef3ceed4da280a33ef924f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ca9575c203777bb06fa3fde227391fdb401fb06d10e3369d79efd0ee1c37221033da20c781fed7e0050fdbfca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31821e984e664e4a4308e18f0f82f79db1b782c3368d7509c85d59a89db5cd1192e7c55a8f93721d6d78b90abc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17123dd13e7ac823bc492772b8613c6b671829b57418e0721ee12380cdf6911084d867716c7c6c7e841249c76a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1637ee6817c53d725077849a9827e5eb8e0b38a403e2c80e06ce71f6d377286ceb0b63f18617cf4226010ee4005;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125717a2a7c52feb9501663db7882fda90b5aa8e4ca1668c74436b0981321f7c46801686c78ce0f869bd14bc2a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfc0d408920f661ed0867d0f57608fa4eed4e012d648843cfe31a9e0b2f7544bf0d50d0221849c08cfe0d42a83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14968ac0ce7e5c60c56ddc2eace013439bd2d9e3627fc3ee7de137af1968785a11425370d0788a1b7bd58c7614d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae00e2925a02a7c336fc0be6c551726c36d41296e7eb2980557cef3267490e1d8fc3f41216a052ee271b3c67d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d66fff1bfd9c4d2c965fcde6a27b8bdf457aee4b068897811e6b2ba0d2fcd5b93dad1c35f3a88b3a701d5e4229;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c183dd231d7c7005bfa7672f540ebcff77f7eded8f8678e63ce01eccee9df18a8b1f7ad3491603ab02558dc74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4801a84cc6b5af05c5c508f61774f22a94d8d8c164c8f0e8ea0680ad3c644bd622313ea0d48172374e59cecdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h391093e3a9c12ccac6028aa70bcd962f5d9b0a0efd0737facc3bd7de85aa5650c8e82c317ca630919353af347d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf33696d9a8a3aadd4b9ed9bde57a80cee4ee885955bb81db801cc8134c18b2b8c7a58e531e64db7c5dd6c31e99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fde3b083858188d40566c844b2cf39439a13480c97947260f58ff209505029b7509c6a5949fd7f603c3166ad2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c2379a33843efe4e5907c52c1ac6c920a9c8571e38d761aa3aac0f20b87839050d4b07f5df65c07433894451;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha73fdbb3f1244009e462f7e38d1f6fdd79bebe28ade0a5778dcb7f2e334661484a025e47a958562de7ef660264;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c6e82dfb36988079ba7c46f9b9bb89bd1d25175598b4a5fe6581379bcfbdfdac20a26dafd8219a17e155ea57d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118d0aab0433e87c6c3bec8a92d45c3d9403da96f92fe75ffca397e2740caefcad469557e444903b71e4b72ca93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he828ba3b6fc6f1d5bf98b6e7b6ea2d0dfdc2a0225f8a471550753dee83c870e2f3ca32bb70cf9b1243538f5654;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1beb18acffeb87075a458d8e17d78958c3b848fea333175cf7cc6d95a69c8c85d1a13a79718a94923af3d3c763e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0ac406995c7ccda83c284a30e61e4aa807453cd2b9217b0e2d83464346487b89a0529bfc80275427c46b1b512;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1996ad7ee80096c420219873ab964af43268aafd9364da619e6251fc074859729f6b3509529327c693777a9f3cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172c4ffd4766b911f8b10a5d5a1937435759ff6c70a4eda9de0c3e42fd5af78d68a7867187cbc01e3b02e10751f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11907d3eb4e6d54ee988d415ed5876f82f4a5beb087a2b9e8077d635cf687dc3919637851ec035723a580e0f27d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf69e021a8348f57f22a522611a35216dad533794376911a0af5c43a144c00b999b837c1221f8d006768b77c70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3226ee266be47da4e9a72c553f41d122b901b2ea818ece51fbdf50801d9faadd1f4495adbbf9b1dccb58e8c5fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb18a22ce6bda46d004c6814075642aaec14441c86a9da34659e9ddb7e222aa61dc91c5e14b27bb1623c996ee3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b634edeb1d961069081ee28b55781851e8a29bfb7f09f21e4d6123444887cfd4515ae4db1d6abebab8b6a15bed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5a0405b80fa888e737a302a382f68516239fc35e53e726f5a15ad18f1c36655ce980e7d64c41b7f6a50f2e13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97105dae291f27adde4373b4fc8bb7a1fd68756e6b93c5dc02154afe3225a3836a53e7846b642996c9c786eaee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db0592233aad49976420ea648f4c47438d6a05cea17f4e917356ab589320b3a0163a263b7d875b8e6b5dfc8cec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1018fbfafbad52330dde26ebe05aff8806db5c3eea76d6c195ae8a757e12bf1b6bf9d13e2907923c5df730ab038;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f85b37f53e37b390ede8ffd1499dfcd70cad9a32ee15b87247976b55b25b8e3ed9cc9374ab9c84f4ee3dfc9e3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc94c0fadbaadc0fe0ba30de62c7f98ac498fd352313e05b379927830432a8a0272cfc7e3ccbc5a5968ea4ed783;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cd8003030f74053c8d88aa871e69899cb7a46898c2266f64160b177963060073858d5aae1fe86f2d4810cbb6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198fb16a6a65ee9a020edea883f421b7935c0d6d1de2d0677090af9d25e82e9ffdc3c8179745ac102f26cd6df05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d835d4074956b89668eb3fefc1433be45502c364a80f2421ec2bdd9f85dcab79d8d2fcb1e9ab2add70ed305a81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f1f5efc65f972a614eabed189b4ad31a28d904b4d971e058f94e3a6eb365dd03f0c1170b4575501fda91cce74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80e3c5c71924dae943e262f7ed4e9aa4b678f0eb360856db70d53e5663fc80af7db4b62e676789a21f8460cf8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac911433d098cbdb5d1406c583b10def2d78cf7db1afb60a11213396b57f73e4d933060e3baa0882ec05c280f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13db7ee4f015378c4dbd6b140f0a0c8786f13122fd3e68c98c1562a12853024f2e52585c10123d3e2fb3775371b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd292eb8440d458361a93c563c58db7646308dcbcf3ac6ff414b33e56983fccbd6ffbc26c2627d55752bec2bd26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d6902619a0fffb79942064741732b6a328f4f38c4dc04ed2454c030ca06e3cc9c1df766929f1cfeb3ca97bf81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9b664c2fcb53f93aff39fcc4020a9ed4b6ceb84d1ffe56857437ef7345e3f3d146350c63386bcb84750711486;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4aa4972578fbd907e27906619d61a104f80b5857378243012a68dcf1ed6f996eb72d102635fcfa36d8df142f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a3e1f44a720643f4785c7ff93cd5c13d4a144a9fa23b1b0321959aff5d50641a79ee2e860c327d0d5d9a5a504;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b306cf68ef27d8070f3caabedafbb5d5dc38cc82cff45490e32d730dae506a47dcbcda6e83d3d7b88477c865a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h969240fd35ed52947ba47439b6d9ec32b050fb16e255bf21bb26f0ec86f6e95aab1ad9fe75db19c95f75ee6428;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a11ea0d56408ec2327a51b9b7f14e11a872ec74d2a5923d17ec05f230b4974f1cccb5ca3e85de45083a289e85d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69ff4c13936aec8a7b82b7eec88418421f5b9d6791bb6509e9f537ec3578fd4d5a2b4a7f1ee92a0394eb0f1992;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42308d41b0425db746020c8524d8ae0be865343153e13ea854e56546f68866dde79a0a41b6c6f0fec9ede4504b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df5522e7c02c038f551a3e1c94843234cc3fad3584daf2ede55ba8a59d577569a50c9351a1d1b3377e8c2999e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99cf18185c68b9a4791c614c3c450e64f625a73caff1b922158b6f182023fb1a26a638f90c955dce41f3d2486;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9e0cf24b1c3493c4e397f57d2921caba426217b99a976f064296c4729b89b9c0192531730f2eaea29b6db53a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d8aadba775f5b9bc8f1c3223a989ae36565056e035bc3e69a062165a7b6a55a05d4dfd28b6427eb6a774dc74a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1886dc5a77c9fb528c479e7823bd406e93a7b4eb5c02e009ef9d310c3dd230de47c5a3f5b9df7a9d0d72406436a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133953011131d1267a1aa6615537a534ba60f36380303930f75a23475204b0ef863e48a57cbff76eb7eb9b83f4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5214bb76981ada3115b84c89a7462baedf0c2344d56a628d4915f6459dcb7809de8c328955c46362a3cdab415;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6dd6fe209344f9dba69955126fb6305cef6ab25f70c9fcfe14158bc8fb23112ed4c95ff7cee079c8b63b4889;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194649f7cdee196498dfc7bab90523f5df8231f3b5534ad4b48b58d6f39c70f0edafd8af637f45f8f01b3f4b18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182d691c2650aae70d43e619ffd539bd2f9eb0b788991367be7c62d5e0aebeff4d10b1a3d18c0e144999108de9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acdacbf37a67c1dd786a56f61e4e916557ab4d83d0f8d9144ca3795f1e14456890f13b1e098f42f7bab6a7d439;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45662e747dc1e731999c6648b8c4ea3bafa61bb6dcc4632a6ac0f7e5868cb3b3d2afc7eb8ba8cb2b64c8898cbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f65b339db8655f10d7f7f3fbdb41e2341f3b9a57f24268a6cf98dc3677eeae4bc0120c9ed48b3eb810c0529af3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecdecc8bf91caea0c6babec8e083ca1252cf34ca75a97638fe1a0e42257f2b2ccb0b38ac0696bfcd9a0707f20b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125463f295df3d50edd09439eed715b7fd61aba2d9fe319a812a3278ce33a84bbe4c919c3bb5abeeb5c366d6e60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4dace651f9e8e6d40b274c36a730933508f36a776c93cf72b227264fb1b769742f4a657e9ff1d9ab2a5dba218;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb79c2f40c55511c42d88dd23f939bd993b9775249cbffe8e2325fb065f74924f6d34c35fa565b061115ab3690;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6ed6d7580cd1a0d85f65cef649ac6425e19574a15830fc556ad4abf67f944a35e5041ff2142382e20b7dc1e23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he84f27a83d50022b6134fbce90310cad4acbb01be34e1169dd9a09b6f5ba3c4b6b23925d95fc6f66724b220ecc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1353bbdfcf63d5a65fac1ad42d3f483a2080a52d0e8551f87a7dfd5a794cf4a8f96d6b874a4d3c3ccf5c16aeff0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cdb6a6f9acf75a519223d20768d485c815a20802066731e8352dc674bed6c46f9281cbe81906d59983d3f2fed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8ddd48404640551e6652d5d040bf0ce626286ac4dd04defd460bd9c4e0b4c6cd4b17ca11fe4e83e2259dc9d60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72f4a432bb9503ee8cceeb709baab523c9c4c553bc738a67371a45f873eccc0b45ea180507163c30240964a122;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82b454ed160cf03b1c62a484d8c37b005a0c83421a07a91abda35d87d0d4bb7959a40fedafb0e0131e51a3c3c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b32d236df0f36086b2e4c0e6bde14e006e0255b2b093af3868375f15a59a29d690ec54d8e62b3cefe1d4ddb46d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb51c043dd44901eb609686293b90cb9ed9371dc3419f0e98befe512a9e8e6680477ef7f88be89a0c56a7628dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125d370d5ec621761b603ba79e6cff002a1586e6ee21b28ebd8095eff523b9726e23fc79b6c568d9d8e76209cc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c80c8f016c80878ae3a5cca01fd45f4545ff3bd7740eec6c215bbae67600bc22d6569283a46044ec0fa6719851;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134a382c8d8ee84fbd27991f8a6ba941418ea76853546b189b849542bfd9c6c516cd30f0331f0120a6d93a0acb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e7541ca03583fa272852a36bbba0a465dbfac7854ad370b6a8ff7d0a9a3fc0e159049e44dd829274656c49cc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1356dbb9d214a244c23a1ad90aabc5e94b47ca2ec2ace16a0afc916f43cfb4a4e41a706ba10d14324f43a0b4a39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6c141704e8c829faf370994d13f5729404446e4c60a9f383d7dc6e5d8147f4877a61390cfa4c8ea68fc82a302;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17526b7b36a720e906238759797b32efb27cbfdaab042b8a7b6db9a418d573c4e1df20633488d87464b867a4875;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h680092feec59f5ef5232a4111875094c443a0bf85821f78a8ce8a645da7ec6cfb6af6423771e9d35045c3c6fc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147f968a1002473c40498654dc5e3c9160d27f12247968fd32afade6561c0e40a826e240406db26bf5529e3880f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3d76ad775bcbf2567742c56a8d1fe28b1348468249b6707f1a700f4064d79877cfd3e3a141ce890efd7551bbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183ee124d10d2daab2117cdb409e2bb45fa550cbcfcffff61f89b4198e927d2e9f6b0f24632790843cbeae0c64f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h842abaecebe0c552454ad7899eb76f5ef0764487ddcdc6f489c2903f5f8228160af5bf985616d8b408861b3434;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1651b81e041a7ac6c5c7ed7698c2dd36a009f36e8abeee70d0ec31d995daa6b122e55ecc5115092a1d1ecef8d8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135e9e19bc61a4dce9a223a6473676991db94d3047bd3d43e4a4dc4fc03b1ebae30c82ff6128192d7458ad83685;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15bae053939c4d26e2eddd760c27f7aa8720ec760567cbbb7ca69c7843c0ffa2cb9e8870693f9bdfd76da22bfbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1707826452bd754ccf5d1c4c276f9e31108fe8aec0dc8a153ed796774586bcbf3237fc43d850046edd426c447ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3540e81f317b8241a051ba693adb2f5202a44ab59432acb7035fe3383c68f62594cff4ca40af7d474e5bee99bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfae007c3422f87bebb479b276788c793f90bfe3b439319b961987f418345703306845f355690a661a74a8524d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9adabf9bb5c58dd53f73a88a88b058c35ce2c79ffc505c6c310b37d35c529594c97caf0a2d198cf1924585d7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf656653b43b16d8abdf41cfb73c7936b36e92837d5c87cbd94cf1c45720af96a0617266e5a520c0f7162a59be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19db8bdd2a66bc984228d49b7c45950ba97971f082d6a44517a8e54d9ecc983ed1366d08dacb2db9abd9a7e5b07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he09a014fbb10273f8ae340265953e7e1186e9988a38c85af04e7f201848cb35532b21a57b6e07ac993e5ed3fc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1550a2d047cf1741b0c0fa4ac971d291be7ac7be9de8e362823467624c9a21e066f49474b854fc2dd6deea09720;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ce996b5026ef176a4453c41a12ebbe65e5a2a9562e545932d89f655a14259a46c4cc946f623c08a3c0b1c2ffe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a542a242d3548294ade452a20e50b9e4342ba0da4a2d3591bc4ac31455e17964bac1d3fde9a92cdf9e2e6d59e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb3ce39af7b94484d843c8938dccf3ed43a31ae1dea5ff392344ec3215181ac4320db753806bf8ac692db225a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de1f1b657ed5138b216d3db84337a13b4d2e6901686936fdeab34c5e494f1c2b35e14783b7c9b4c16e077f90d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fdcbc1a51bf9db48200a8b0f83518b60664252a2da8c1bb68e2ab885bba18c4793fa39a4339dfa649bfcc855f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd3acfe70f2c64f0df7678852ff872c96cfe80c55316030d1d4c30c38fdf175cf1de1a275ef541f000ff5a4239;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb778965d7090070b1397cf62b9efb0f7b11e4fc2c12bc7f37723372a5294ca6d33a9acb91d259894a4cfbc30d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46e1241390e940b7b255e5f29b3362dd306fc1ea5d9c1916cc30944dd193bf1ec1fdd031d1bbd28fcca515da8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b638a75e92dc51ed71753b0606710bc749105051666c7542ea1d94315a8d0dc323e7b1cf9e5603bd729eaba69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17023d69d1477bae954159c0f936293d19b9ffbf081b3cf07f2dbaa2c262c52dfdb5c015f4b9ecb2d36b505ce22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10dc84df9f3ca6b760afc659139b886618ba5adea2035048f3c2f5999dd200bff256469fad7892897ed65cacede;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5aa0c80066de289e31dfb98380828727d08bf42abb4537d7e9e89d860a1e45531eaa9ab79cb5eda21aaf9d6329;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad6e3f66cec7a44f7e9c1174f89876ceb089050464de8191750c641478af89751538ac8b1630e677749370dcd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81550862dea3d5eb0d62906819c575babc7e2750d7e3e641f61cba14f6c617feb268518cc7ba649978812fdda9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77f0fc08b0fb16059a449dc99467d14168c3cecd25ec23a02b19eca6778a1e17894da12f00605630f1596244e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0d94c165b53b5ca7adfa3a5883124ca58541e7c9059d2fa744879693ce167ea10321b2a7a784bab418e403212;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c56191b3845187781b2029c8f535147b5492d9dca06dc3485c513538abe513c8c767790300e7aec206837f5378;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa34fca2ec9772be5d6ed0a2c63266b1b87e1505d5b35dfd6d5c78c7767e321e7197c4bf772da0dcbe0b6a8440;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12624e832eb9c11fa6de723a16a1eadad7277efc41d9f6689c84b556bf1345cb2b1a378a2dcd3bd56854eff2bcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e105f48fc381e48726a913a3062122dee4af143a2c67de9cf8f5fe276814cec6c32f8d6fa4f385e300e441650;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4da589044b08e88fb2299ad1060d847f96ba0491a66008c93384076134062beff4f36b6e8966a0e7ce49595a0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e9b357813e52005b9b20597afc4ad9ab6c67452b519e035a5f54825718adef10875e732776e0aa1b8f4820a07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8cfa242aa9287c598d7f6ae3335a1b7996b7d9f3c884d852c7ab3558ab490f2965961561a29475c1a441b1f2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103ea77b05f6a8fb09730b0509b58b711e8c5f93bbd0f732f6a5ccbe046b1c5169e0aa318d2ef320b0711284ea0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a1cd46b8839222cb654a089f0b1d71333aa69802a50d6fb5a0c12afc263d4b5cea989a902933c0c7702f6433;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad8e7b0781d72c2a138a9ec5c2e5c39aa3dc6d263ea2114d947df77ba45c8d609ef346d989879a3b2da80b0e50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefdc1bbe377fdbfe4bc2dafe333041891d646fa38ce1b9d7fb01b899b378d84300608275c799a60dd92c865735;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf7454fa530dbbbb018ef953d22db2e65915a4dfe057b14229752a6e0716e15b07792a227e53aef170107f5f08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1f4ad15460bacc402aa95207b04931d4b72103424f259e19713af9d06a6edc61e11a596a8bd0ce4ce8be7b66a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1325a3f355c9766807ee9e453e20bbc23ed9f9455d5acfc224b48bdf5db6e8ca6bf919826364d611b4f90bd9fda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0fc0f7b1f144abb2ce16448b7f525d101b749f5ef4c1a4bc75c2fa04e3cb166f9ca5f351270cda1e076843e3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15cdf6a16972243920b6e9842468fd5e3d8d9c912be399f76f0d96440fc4e15dba82c85fbe3915303299790e585;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a738369025b008ef48f74128747d3abc28733003a04da4ff2bcd4f3da8361ab5403ae8cba7070884df531edcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14bdf40e1fcda23483a8377fd3aded51db50ae28ea5ad44fa5cc0b5ad86152d6f717aaf0f7c1ebe1db6e786fbce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef2c56e4b5a120a0819a9a8edb03725b8074ca407f3cc65fa7f3f558a8df68011f9182d494b6a6ac9433c2058e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186af41db8e5359aa9c577d9636c2eacabe6bf497c6c4e414c7c7dd437efe76fd1dad5e7e9172725216cdc7fd94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35ec76f4286eca233cf409dc7e4476b70afe16a7e06be6bc70e1919d9d6ff8010ac2b3ddb50b74529864750658;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3eb99dc2f43aa8cf22ca4a556762c209250fe8c9a2b646d32ac99974c4c36c40c32cab11061f381fc6a773117f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d2a0084c731ce2534606913a74220d9e152db22682fa936e9a9d4e86f6cd2758f8529b0215e995233a55f8863;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1904a967d813b9a841a417041a0bad65feca685b8ff064db6b5f55fa3bca70ded76589518024eabeeb8f5a21914;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12eda3436ab44d246b7ba8d5bc078818b18105c6f64c38985316af0e29ff782e5907402b5c7559d9ad81076a4ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fd0ed7b4ccb489e0d3339d2928a6a5aeec91b64664cd09db2669f6553b5b04a09ca73ff6dfe862f405369d101;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76f47972e155c80d90067717405bf8fec9478567e6e75d6be87ea76bf5ecf522d93ce33e0566e25b12d6b9d78c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f01c7c66a20be22486a884dba7de3266f89684333bb59663f99842aa6cd5da81f064337410ccb486dd00893d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128a7fe5d0b29dd92a4a554724d52dddf92e9576d9ec4724fff0b4bad67ce782ca2f5d5dbf6e37a5e7e0a06110a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h920dbb876e66869ba07d186f3f0a68cfcf3322e94236e443ff52ab7940d41ef9568a5adc4a414e57fa419cce09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2490a984340d37e9e0da18cf43e2bdb4bf2da9a9fbfc0637c28f347c3ee79cd40a247d8da7ad772b1f5da0dd11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd4ec1450c28f69d9492cc7819666950b30b2c5219dca580e77058eb72c7d8fd242c21a0cc69a430b429fc566c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d691d5c7efa486741a81cdc265cdfa0758a7f43be59738a6d1c993aff5237435d4b75e6ff39ed5c8bff4f3a91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f03ceb04de7dd3b43a168eb596329a04ae4bddd9c84ae1bd64199f02e61c2e32ca1613c25611cb4e8789788f8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1570e15657d593c157dfa53daa9210c2f5693754dcb1db6531c5728049964404e64efa36e67468b325b03b33f31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c8e23ff93024a673d275146cc3425e894a0cf6bca96535139e623c0e185049150848f538118d4614d911b23b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb54ef282adb8d787ad48b364ef2e225bfa3469d2a5f5378f139624dd5a85cc0978514327f3e89614d403faf31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3bf3e86bb38604d57909c84c1c35b6a4313ac21cd79836a192299328d939c105047cb4ebdb140d124aec750fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1055963cfba22ca819d2df7745a1ff5f6e99faf1809f8941b85df490651f59c44bf43843900f3de05ff23173b7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cbd0e50bd092776c0f9b2bb539472027c2c62feb5272f5fbff21aa7fdb5deb7dfc7602ed6f4463d2d98670741;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a98b768fc172d9c76decc4185043e3058e9762434ccfad4a80815898452d282df2e85d3cdaed8e9f6ac07eccd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1e4d7bc196f6c6c1b81103f95b8cc34d54dcaba039be8f82cd48b06d597460b0d159f5a6cea9ee6d63ae80682;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136ade2900a93507a5f86307011d153fb76f148bfecaea43bbcad4e1b2962b72436d371a606ea7997e3e4de00ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b455e0ec13b777f4cd03991b06c2e656fbcb07e72859fc89a3c2047b90b516cf98673d33bc6638a00078d8f59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d49d2e776fce15c0e1aeb9cb40e64daac62983ffe7f87ae99e6fc20a11d0740c5f39da6ed6c8df371163a332;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfbd90dfc3c916156f2c5f2116eb86ae782d8acc4e448275ce1118d8848f090f3486e3ff52e6bb786e7aae417ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb47b54b605bb5c56531387a8c18a0ece3067a86711dcaeecea50ec65fed83037ed22edd08dda450f5759530d38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15810fb18e0a4a26e04e700fa091407cbe5ee40e7d503046ebc08c9ea471934fbcfa5ef55cfb8a2ee04401e72ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1771f33179c7b7143bfa7af301bf5bfcc4798b94b575e702d59468b210ee0571313290107b4d7ec96c53c8b4bbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc53d1cc23b39da0b0bcfc02af9d81aed6cfc6a7b834bbb99c2dae4ecf59934a567ae0dd94d1ded4a423c77bac5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af86a20c357599b51bff73586f2bb73c2e0e664949782eac3eb45ed24f950a1200d3ed1b799ee798dc1b59366c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae9f3442df2ad35888ac240c8a6c05ced7861228164e944ebba136793c0014f3303f3458bad4761840426d3ce5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63f9367a62518ee651357f629a0d4ffb4be5b6ca29e054168abb47474142906bc77068c5be218f0ae16d1f6825;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1108b187d4c72af03105d3a484e0ddc32025a38eafd69079eb581ab9d8f52b5aca09bfd18c0770ccbc22cae7dea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d26818ca4b9a494d337786cab393434af3b612706bf825ec4649dd3e179d9445b9585d7cb3981c93ece8cb3ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39e74743fa4d31310e0fb4b394cadaf4415922baa6c059c71e98e2d87718d83484260ad8d5379a12d086016de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19edad4e8d5f61c1874ff7eba9645e559e6ec34b8842ea1c37c5929e602486aa0700d3c1f3637556d363d3390a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12785e4076bc7585fa044cdc8a6855df0a15414a451697068ab35a39423ca7cb00e6ce194f5570be02606d61ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f738fb59be3bcb90cea80eb7f700c02bb37111ee1455fb077d0816f3cbc6588a4f50105362e80894a22e350cef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd7bb4578a8d2373defb1768fff7b1aed24e0c07bbf0e8f685ddbfab38e813b60c0e0e473eb2b75c367fe21f60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca19f93f1fbe851cfe72cd2ddae0c4234e20327ee2e7b836dfb9b94b88db5e6b6dad8f56e8c12109e199029d92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fb08316acb4d8091c35daa754e8831eb9b45590003f3fe12c7371ee5b9c657b205dfcaca6164bcb1c941354dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha94403ab57db4bf6176b6c640cb0f856c388561791f8ee9fe8a3b8364d523a415ea175f37c3b3e3618248878c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ded32a75dba7caf1855ddb0b29cdb1b4b38acd9e4568cb4f047e5857ede408c5467efa30175de20652ff02a4b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ea793d4ab5a9609ea2dd0a8b57431a42aacb1b94e16223200023512714db8138498c3800870647ad00fbaaf8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b22defadf4c60499ec1eb91a4a17c30ea66896682593b1746efef8ea9f8007bb221cec747d49e468702b82a074;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfde86630f9707001e9388cab9c7e89bab4cbf29d704b0f086f67052b0f9058a88e315f04474e0663b9e73d3799;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2eb2a83f153fc3d0a9e9ce3005995bce910eb6e42373c5b3278279104921dd29cb5e48ea3ca9d8cbe24ac10ce4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa4f03fff7b399cd77521cd522eccc1e2df0e2494cf7ea41df370b08b57056179cbb02b1be67b35c92d7b6201a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8dedd61cb1023ce80de15b8fab41d8e7945ad3ce4c9214abfaca345c79eda737f6b764dd1f756f7fe71938c46b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha63bb1040bed4e7083324fc7aa1c4625ddee535c65f81baf37a2ba0570eb9cb9afc8839231b376d84991048524;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8b60604506a37c911473223fff5d0cde9d0a2fb6b9e1b4f972f9f79c6879e2bd628fe7e333a62bcd5e8c748e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175aa1472a02bd783b6563eb868817412c7211f859a41d5763e29c8ba4cb5a0a0839a8456ab163fcdc03ab20c1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a54fc061ed4d0b1591d189cba47fdd7a0ad6f013d022409db5cb05f943e2f8ec2cbb863274ea7eb70ce18c52c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ee06c381e74e54347f8725a6dd9f1ca4dec85b65fbb30f0b3f5ec49d2d14e20912148ec096e1eaaa5911fdd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ac5c1f26abd571650bba8fcf581260e6928560538e9747cf5a03568a6a841f18ce6d2c3b36d5584c85139301a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd1c54ff098e506844bd0635fbbc2a9b4aa96a7580f094e076f52f45a3a6c5fa9dcbb66e9875bb64236a7ad870;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18aecb8140e4aa8338f8eb4a1b6d0330a2b2dc2c546d9ee1c0f417fb174263fcc92973683ca0fbeac333fd8e505;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2a1bbc59ecc5276914b71283ed1ea8a430fffeb7be4e41744a5d17ed6ab095c6bbffdedd164f47f430aa97f80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ed2c5553af963b4665d9be20004654a9107c16d95b23e1270a9869ab9e42822d1d0dc3bd23a51aa02e6ffae24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17fce06c0376f0d48fa54cbe2fce363dfd29b81df0cfcd184eedfdeddfac7539cfc355355f1ebceac7620865ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d8d931776e36440600774c478a5e1201b356a9c2ca7e983e7c572b305d0971c97b067e4a170245f671c9ffc0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e57094125c0f777f33c1250ace9d35bf75bd96478b9aa42111d0911b53f73a91a1ee247952d6cb1691d04d7620;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50ad47a26c5f752d3dfa011bbe04d4f4f9b42f14401921a1951629c9c0b2b492ccbb6211863f5e34015a513b96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b05cd1c2f86a31fbef92978089c7e0e759dd142dff17019806a01544dc2f4676e5887ac12ac27dd2c1703940d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2ab0ef87f0cfbebe58930700bbe3a4efdec1968a72944dc6431a2a46df43aca410f813fd23b1fce553793db50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb007f60be60528d4ec247f6177b5d66b01daa878cd283225defdff475a0cb66d8db605ae474b9fffd5773a809;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6c53a7220ab3d515189d4187880b7776df0c2ad812c3a60f217c4a830092aae41a2bdaa9c73ab4403120ecbe1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80ac7764fc12ea6acb454aa465d2086edab11ef597b7f0c52d46c0a47c749e1bb7b98b4c2af5a675edf8d1c298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b121a848b454f496951c186c8f8e499fec9af7e533640774261ce92c95043741d582cb48677ad4c7dcab9cdb7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb8faf7eedc5513bf5e00745de23f2eef86c70e0fb677bfe30bceadf83ab0804a9c1ffb7f690318a178948b489;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149168e0ba9de85895f3b4c81f0ca9fb5b8497ff7090825f6233279b0b828f1cd075b2b953fd454d3c755e43abb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16afb99c7f26cf5b941d9383e92e16dc4f8907be52fc73546bec833a0838809bbe51d22e4db45223c0d436466fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffa656c73f39ed8703f7bb80b938e4349c434840bb54cd7e5ff742d8059515640e6c9b768d883d41dcc5a945f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebf56e0936726eaea436c4be830622669eb2d82282251c0f2abf76129d4de711c4c099cb5ce3d4738235b23dc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6bec1af7c44302380e758f0dc0315e43004457213440b641bbe7300ee558d79d037e40b681922077974963ed5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7426fd781e643b54de6368329b78c050781e39f3de27f6b86db5f215925fc8a061f5cea6fcb50d7738d89401b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f47aebb6d1c41ac602ee99e3501497c876ebd93cdf52dca78663ae5207fa21acde3d0024b9908a445509324c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf81517e251cf538d94e054de1cbb01cc4b556c820a500d7928306fd505ddfedb4f0ab44878904ec2bb42b1f4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11322ad3b628b83d1ffd690d2c36eef2eac96ed206f01b98056818dda975c8515cc7d68b69f167f8948cb636b6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3eef61f95b0608fd974548876936e0d967b050caf993eb4b3006a0f8eb3ce365e65cf8d56a9a02f7b2b4e0abef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e23b9d5f8fe2ffa07b1da4de636fab23c80af628f1d207790392f6d6aee24da2400339fc8491cebf44dd78277e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8868828a75785abd7ab9f8e54aa3031c1e5e2d5ab95b5d94ddfd9d20c717e135cc3382a829aa13a3a03be8d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fbae15d6fde63a071a601819202116dccb79600e685162ef986921d236f3bac3a2d85d10b0cbb3daee7bd921a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8bedbaf0aa217ea625f307bf47f706d58fa643e9637d147b9ee15d67520a33cc5c30cb10346482ac787b5b88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1040627751dc378665b3b8a5a1d8ed2b1643ec2328e22d6b3706b5ca3e72c7b202538862242fbbe43e12eb83d17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b5407cef163a6552a15912522d9873c4156468ba656fdc06198077d224718be1df8d1efcae7a173dafd10f80d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81bdeea578a6b5decccad10281689259a3c7298f210354efc687221670d28928c8ffc3c991f13d8b4ef9626bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bfcb23a1ce46621292f6abd23258f2903fd35561fbcb431b5dd60fc733b8e0dbe080082e0b1dd39826df71ec47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea8ef7ed2fefc4484fff9f6c644f5988abfca490dce5e7784dc5ce7fcaaf571d2a7019a06682272a9015d2ecdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he149ae36abab09d78adde5dd74577945be7741a25026eac5de52ace0730ae73e961595b90e88676f6ca1174aae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3d0d1740e2093071af9222b855a1e8a2361dc66b7bdfd58b9414de84f6ba43ac898c19f345744815812a6b55f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1406ed07def5ac0d6c2689c90d0e65f564e037d329b52ee83735f6299c4abe04459372d65fbab85a7818abce292;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a25812cbb189575cc579397f9c7d72f5b55e70d6515911c7e2de2c9bda51ffa4658663f16e8e5bde188f18f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d99995994dd17cd69f08c07574c64f542b915fd02fa7aae579d6917c4293f06d391a586e4cdf94aa5fee671499;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19732b0a156cb458c982f3497bb584029d6125957ed805f206c9e3d88905945c4146934dd83850f116cee40fb01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f4fc3b5b8596b1af9b981a0aa5aecab4bf51954361ab8ea415264e7a244bcaebf661c4479503b00fd764601e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51732203413c8e2b6357c286028fc134edd00ad247e047bece9a1393721c7677d8d67c684533847c3b99d96906;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20bc98aa020f229ea5fe08c3d617c6fbdf0a936d7513e0ab3fb8ea3a3af4a3c4948b492cc757bb690da3acc92e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f296046dc956cd39e4c4a5337288d7f1af74f5763b342b618bc2217ccbde19d94d63204673a6dc5b947673e096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e6abf7c611aed2bfa4b702720792576210cf50e93537e1884c55f1847034e570ff4ddb7830818936e6f204a31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be020710351bd7d353ecbf2b680833cc0497e69aa3e0acabe381f4e79cb85b11f710c857cdf3d452dfdef5c359;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d398d98df399194f05649735ad1c0d4ffafc8d1d50b938711852a530bceb654acc62b1f2d89af7e6625f59d68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had6250d85899046e58c82f9a1b2ef177cf97885d7ab883080a02e2c8e5af80d58bb293d868ebb18fe90fe0addf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7a1fa61d7c71b4f3edc6915ad5924c2a4c560cc48bc9f452993763936f53f7948b2a49e34c9ef074301e697c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35e498f9eec9a9f17f9ffc89293f8791ccc68b05d1f19d5c4cc02ed425e360d3190a9616b847387f8472dccaa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11cff7f7d8aa44fe9efaaa03330d7ded3496f74dbd6aa46dbae923ea413064340efb321f9c15ec2a611ed001324;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bafa12489a96fcf943d6e25b12237f0b63a03d077e827e82df9d14e298c902b260caa51b920424c5fca0421a8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117ab42b655123f69d15beacad805a04a9cacfa2cf5aa8c0174467a98d2c10aa952d9aa7e9f99fdd02c5bd1b93a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131488844e275daa58a15be01134792eaf34e5f81d5a0054721bdca85b282b6312721713f3e8859474160539f25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58c3032c71629f0a2162b69b949fdb04a614565deec0713994ff3bfaf4c0412ca691d6729850cafa1d1ef01f39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148beb79a5647838f2ad6d932f6b9cb7eed9771c32f24a87af5712eba6cdf10b8bfe72261e90afa14d5ddf74cf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fc18a0a816814333ddf9e41d6b7a4aa0f65d7c1a0c9adbd31efbed23c9af349f2f2974163d478d8a689e946ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb46b9e0281ac7d4bd7dcdf66bcab97c5cb3e214769bfbeb36ee1b0800fba4cccca7ff80e97b1884ad4e910ee5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb2af3b9bb706e6776ac9a65332b840083709c8637878c366319307a1ab3595b636ad14b9265e0cdbf6850f250;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4bd167415036fd6bb5e5d310b0b738b3d9955e2d014a00d8077732435769177607f09c6b085d28e4d4458a64f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185590e5fac501b4b099b0c063bbe2f78ac5cb823fd25862045b18cdbd011d41a80b7a547ff3555e4ef9a944809;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d351527a32d79539b47a4af536429e33b3bdb0b15ebd63e05e2232076450c042b4a4711472f7a634cf49167a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0a62290743abbca55cfa620fcb55060c44cbb944e19dd34e2330d23e6b43512cec81150b7b6817dfabb7ff116;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fdaf9e5a26b26200c91624f646accc865a93382906df6cf5b44a79f7d7bf2786633de341161aab86cbd6ca15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h21a67b5d3478a44f042a591b9a412099c6850339fbe07ff73621e25cbcc4d4d9fb8c740d875e664daa09262ce7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49aa7aa9d77ea7fe3f389339f4ef87c1c12b8dfbc63a4338ebb26636d0224a1bf74c57a73b2fb34449439736fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1540449822b5e8e0e1441854239a9c1c364d681810ffd6ef58ed97973d9d72435d7cdbddd8a817817e195437be9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc4581281a6bbfc11492c8cc931aa769433b75fb051382e91341086177087a83d7582f3c4c05b36f5489d1dc81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15116c38f586625bce31d31f2b06808a3f29873dbcf83998707b01c8179de6e5e906b1956bbf0b03e755511573a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd116ad7df7efeee8b40b47e3f92bbab3eb9713c2ca8033fce438c653c06d8b9a4c68fe5ec48c33d2e8aad9270f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5d7452195cc44f0f8775b9dea8bf7000b9cc1af9617a08954026d1828c85f0f29dac4835a3f51c68f05e88e47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7052765448d154b9c40a5c577374759ae8449b45d23fa33a579e73ef531992409af54283dfd270e453c0739c9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h162993c9550b15ef9bab4403ce246b5da4874a7a0917c229cc679d922e299b7326f8dd3c7e8e5a8b4e4619334bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf314de9bc8887d4135557c3a416346f6175b1514394d43d8614ecb9ab2d7674dde8ae7f0cfed6a8b88aa455bc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ffbc59cd89ca9258b08d4e45ca2014fa7c2605f79cd7a0732edddfd68e8220a728c99a28b36430fa5c0a8def3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1234d28b9946b0bf490bf48d8804d2367a3204f3cfed32589b75723c0f9e92cc5e68f3742e0caff6d1fd9a57687;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd60c6bfcccd1e290b5ebcc00d68d7b054407929b6697d13d8d93c68a0da81d921828a640a4b0b2a02e48ee9c3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c680efaae4d186e5435e98ff590c077918e898d546e08e1d83b406aceef13f8653ac38fed76cb341d460aa89bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa94a78f37077f42f1b7b44995386c1cc815e71bb0a560470348c03b82d4ce177d0c805d6f03744c076f6bc36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h869df8bee14a0a72564c054f031c3388e7a53fda34b1eb134e8732eb9fb187a273de47f80ffeb3e1adc8441cee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bbcacdb9f5c75ea2304fa424cf000203722455b381d9bc841ca7f4ef2d1065ca3daba30df2fd384109821c8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109632b084f16e08ab15aef492ae5984ff042c198a841d2059789b0c27a122c95f86f772f509b744b5de42ffb9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47c39c5adb84aef2527760baf40e501e5b93b7772d948a6918f4868959278a91691cfde38256de926b85af3fcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b7a14b3d59176d92cc180b2ac3e79591431ca5321ce1da7395a2287fcc428176ce9299ec493b79a11436213d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a698e98f776a263f2fdb234ca01509f2cc37f5bf4f29b83aa93a3853efaecc1dabfbb210079465883d97f99aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc02209cd14cb16ced83301ef4b5a4f61f0a942b94ff7ad063fa3943e49a44f0021e00bf1c150261ce62a3a48e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19db6aef3374598ece975228e9010380bc98cd5473fb19a28366db8979ddb424dfc30ec8504a5faaf2cd0e6e007;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eace807c00c957687236155172124c2e7d561380a782e436f397a1462c1d9073eb98957a1eb390365e461684e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5638cad8a1cc819994132c53108abf0e13db441b9ecc3825247b654a501e723e8b72842f53fd0af1b07c10cc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h633120585622ab2f60efb6f43928fc7899fe336b190777210e714380eeffa6232c280c8687bfdd337e4d6e3e9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a221c045214b65d4164f297d914becc60a2562c5cfdc2d6bb328dd78755f68125daf04e1fed22b245ce2127ad8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188648fe48b9e195f79849051b96fa4da24d993b8b8f382ba44e295fe7907c512413fb0006a5620d3363ed55b84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3851312e063b407abcb7fe536cb8378919812c5f3ab020cb91524f95b35dfb704f7397ae390ac75f6988ff74f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7b631a84149fdbe7872ecbc704466f50bca3242392237d8dd5210c9719997d6b23b9f43e8b8de7bb36a1e9021;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe9c68370985b005a29bfade6186f68be41845da0156df3f0fed3a02da57a5103ec383d67812c56f43019c4322;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1689ef12faeeb43248403fe9e4eb7a5f194c47d0c0f2d35f739a75e02e6c81cd4d7ec3507888a9c48e9e845f34e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140a708f5e0bb90cc98e868f46f4acbf369a99bb102e01a7eb2a0cc4e5373f3497274476c1100cf677324de90db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9edaa48fc91c071808fa154874e2b93feadb4929bd9b55d8f3745fdedd269a32f59c442de08d26c56469138fb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac806f0f60608bf7356fdee4fb130f181b1cd18cbb8399f058b507832878dbb569cef8f626bb2a7748e3f8159d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2553e261e23e4b40e63e7cf3a0a9812bb47f5b280bba62c157e4a1d9cb72dfc735406ff65b34d00d6dcb7869d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h904eaf3ba8e66826749d94cdf658d02a609413625faa4a8f32e1bd38463812f8c600874d2cdb15dd08264275af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4aca4406e4e3f2625965a45be534b189df9b5e2376ad3d0241c44280ff75e5cfc8fce9bbd4701aa245278d46a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb385640b4eac4cc1730963e78bea63cd69fd32f87997f4036f98a95582e928afbcb4fedfa5e9cd18bf72d3473b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cb75c6bc4bf817a8294cea925e56825679fe35aa6b5d3a73895575a9c72dad8745038e99ec69742064429d5f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93d5947163e2349e8fe95843cf39d8c9807b54a402098138dbbfc16964dfb2f3c99aff4c6d17be855307c7461c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26d5fac47ba6b373a75cef38942657e53c4932263d9bd73ba394a35c0451c64de225656e79b02e299d4983e8c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a198ca0cd3581d7abec12426f7f8c37e51be1d47d97993a0d8f25556d7cea9a2abe281865b1d8dfc91ce0586b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce773eb1120a0ff28b04f463e56d7a38b6d9402e09975e5b75e08285b6f722fdb5c851d4f68be7e99be005d594;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d978658d83894bc7a51c41b19778b8b9fd3c14dd62230e98db965e2b2baa4294f6d59233128526dc3b00ed6ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba73d0fe0e605341ed85dd27dc649ed89b32391375640d8443a1f89880444d4eafd12b847efd2ce5b85f3ba085;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1787e4db6a95ae877e95bc8f14bd33f52098077f37122a1879af647d787412ee55a1bc40f50754e965f3e22eb73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cefd14af8fc20901da15c3e2c5c51ebe63327e3e1d0d69fe72cb1a572794f8f7ff0c59b59e96e3fcc736984055;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd06137230ab73e240c217e0ca7bf24c52d17a2e06bae8d21e5147e41bf04316b6e776be29fcf3c4c824d214136;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3931ee9b1fd777ff777552adb984a617b1ccc1a30845ea7fe21fb8e07a6ace5da9edf1a3e9da6dcae254d1da64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecc7a6d711c5159dea7601f2f6666de7c077ae34ad09db331a9e49b8559d1530fc95ff738678f4431eb6a92e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138e547567c3b8158fdda555cb2973ae2ca976dad99fb0f9aaf43ad9f814a52613d4a7cb67ae23500078bdea1d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118f5683204b8ac6acdc949e9e11e0cac10842617d4272c65e5f46b11d987ad03fe2bcbcb6d5f60093a5e99e169;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59c4ef0af824c2d35535b67db2001c9ca454a8f20162460591c9e8f748d7f41b769b994fa96b27714e9fb2ba35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df5347749e648d265a23b1834fad9a4a622dcb7afefb1e7076d83686e0211a898e18450a9befa42e7d092b94eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e4c976408f62a758d649d8a9b86e2a880fe9d33bbf3a761e59614e124ab6ce691ff0e3dde5ebae83d124ef1b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf417900629b32290a484882846934e80dc13ffd489989f5c455760dde0a0c258855da99df3e54285e2d0ae624a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195a26441482519db8e8f772824588fc4733403346ae6222c0e0aab44249c04191a4e171892aa814c63cf766729;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c74f3036c8fb95b17331c0bd7ed95ea798f9332b0b6a1adb2c514c65d66d033bd9694236428f53ff83052ad387;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a337083e14d69c28427df23495a6e45660ce1b423216af9c5c9054b1d801bf599adc19c7b41bf4fcc946d72cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d71da40abbf5cdee5fc092053010c756ff06b4aef85795ca7038bd5ebcb5ab73f92d6af05d27309482656e111e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e79fab38738fb999a55eb0bf0f338e2178817263599a582c4bffe544b52d4c20f28cc10c382c7e2d12cb1ba2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb6d4a9ade4d87eb9bc4932904f9824920efa38b712acd8247d770fbbd29d98c6932e610c29c1223dc1bfd9713;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea5bfae492e9d8240d89bb35924af21b4f8f3c40b70a4d316e3f6061f176b43d7ab0315bf0bf320a4422b10999;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1632c3e44f6b7d427da326c761bdc748c164c9a67cc064f9dc9cee8636d9b1f93c4d77a2ba9b12148c3856527c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156d12057d78335fd2c2fc9638af4374807d681456a485a501e32c538a74ae595509caf5d8ef2a1fb191df4ebbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b8bdbbde4b1006c6f3b522d44f88b55eafa9ab4ffd9519f75332698b5ed1c0e2b5c3d5e0b09522c49ef6f0265;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ddbbb9780e86b591c6a9eb20b46f7725c47b692c579d172030603ff305acfafae94021420d08d75c91825ee4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a25a5beb53b234cfa675aab80ebd1f1260fbf9b547493f9f727ee07046197f3faac7d737dbaa8a9a6413bceff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f9c1d9e177845e7e2db8a739e50454a7733de27861ee8b0633363f413894b0607d4bab124ea99d32155528c19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0f22fbb7fcaf660a0bf4b2834e732a3c2df210f16cc3c21021a1c8fcceb2897ccadff3168f5ca98cf70cf6d5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc57247046093b630ee1e15d24f16beabd584521985cf210b6e9dd8354c7bdb34645f6d612818487e1b0ffb6a46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb414d770f2e8ed7413eea3de2fc0c653e4d4534eb67f82fd9b4bb9bcc7ddfe715fa4263db4a277f40b8dde89e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106d4453322fe05d661328f7df444fac71bd92ec3f2b9768cf32bac080ecee4ac225bb407e2a0fcfb4cd2c7d512;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcd6991e836a0a1eb02a5942656e91ea9b04668eb37be560700694c35be53d9c342d9dc6ac2486c532a2047213;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57477c56c268540a6fde588d2681b8aa851e21fb558810e3811cd1d0abb79d3e94b71d435c46bba505910d3a4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1664191be63ee1993edd26e3679b17bb752dec54da195fdb6a8fe526f05d74e210bf562eaee2808f4b7e856e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128903447f583e43e8b81284665d008628627a77e34571c3067b8b38543a54a1c7465ec9a81b824aabc8e0353db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c4f105624ee3cdfd1f0b6dc543a447089552012f46760af499ec11e7f0ceea10f88b25dbfc71a7b2d0e798a30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116d4760632e2cfb4d7c7c2d186ba6a9c4dd279c8e8f95626d9404345e25e2cdcf4dc5826ccb6e3fe7c103c4195;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd143f9283aaf562e2f540adca361d53f9f1f1b193af811708baf4e830ff128bb47738859b5d6db01f75451582;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c02852aefbb6886ea1935c11e4a8c983455738fd2b275964d249f9d31f3e812e0c176535d284d953a893493a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1aa58d7903540f096ba9a71b15e981d5f6b4fdd1fc96ddb98e9f3cedbd73b752a747928194b3ad7dbe3f0f4f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175d1613e9293912f9b660201a51622c4bed7fa1d75614e8a4bb46b7392338cae54359c5f26720757149242b64f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72e09681be2eb03d4b46dc5aa060605eb288bda9bd19649f734656837181a8b59afdda8f2fbedb337e4ec02ed3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17dc45a080537f865ac91ddcff0778587d0c3304ad4c8f6bc757d686f4daa674db2958787aa67762e0f11ce2b23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c33e4781cb568e6ea800996672d3c7b5fd536a8ed91fc6a122e9a6d1bb8a91f956f1980c0e30cde8849b5745e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0ea15ec5ae3fda53e388c9e4593d44e8c0f673f70c27032b49584220876f2bc23c6f752272c3d094b085b63cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef9f11786a8784f0c376200612c2f557f39907b6349a9040f13d0f7c9d2373b855c0fbcb6ff68b5ef05d231982;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108b134539ed6f955990dcdd8280f8d103c1842d462631881aee232f009e125600f2e96108bb780254b02178acf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he46b20a59a546f74a1df48c9ffde7cecb937e877cb2dfd25c089eb9182ba6eeafd447880a90c63c2c0d0d14720;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c55864af0725a33cd14fc20f047880606196da90163fa6687a88d8fd8c2048578c87b9a376ab269bc62925b32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c9cf6d4540b90da0c73913f44e498f4add8aeaad2bd1c2759132a97a20c04b16a3c9271ecfa46032c4d0ab890;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2255ce62c26d901d80b603a821dd0891f7414078715ec9f8a0fc9154210ad44ad0a5f2dae95cf6ba21ae4d2ec3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1165cc4d3a41ae5726b798cd608c785a5d853f4387f52d6d21c5a19422b760381327a57ded4f832de4287f67665;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fe26edcfc825ac57ff3704b9937c591d698223eca688d29cf43564b090bd2dd43eef122044b275f235b3238ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea3386bbfd5d5ba5c11084e70eb47a78b176614f7b45cc609e91a4886aa565995f5b43a3e6d428506dfb661480;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf310e721581031e1347e70d4ac8eea6bb978d5741285b9e29a6bdd2a0c639e29368aef6795af83c356520b252b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a8a3c7d59646fe96c1a845b73223d0b3726292c96d90c90aac8f22cbe31f067902547b2d531e74b268f9955cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a4e88a219b23eb9f3c4c9e6ecdc8a2bdb294ccfc3f25a6cd781908134cb2daad9935b8800e11b323100b7612f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5284c4977c68df9a52b5b7463c6cb2ba347a8382b9b95735b4159aff912e2c18d721742a06b07937672e86ace5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5789547ac0baaaa0a32192ca6b02bf0bd0e14fbe054a83bd7b6458d5a939427d1139394f31774abd8ec773a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d28d1ae4a3e45cfc5f545c582a89a23667b88c05391b503ef7bab2f778b55dbe2026e237a34c6e5848a512c10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e5d986cbbea7036e7a4e3034db412b133b099cbec07439961d25b409e8c51671f8990d2228507ccd93b4279f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f37cad071eae41eac008cee6392545e3be71ace931c5f79e982e1fd97b4e5485d88f332dadffb904111417d5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19baa9d1d5781eaabbce3b7622323a60ae61e74f284dca1e109ce652449abd753f85263c0122494aa815166cc67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142f0cf747550f64ed3b4938cba018ca79eb22c037e6a66ef8986434410582191bcdeb34045ba4412d50c8bbc7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0dfd2f0639bb596946963e47b5f726082801ca4fe80af110819f0b20297fbc9040dd085b1eb451a09448a8677;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c5de292329089d098103416db879fe1f16e22de8403c1b20971a0c4005890844ff74f9cc81c18950c258e970;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e424c0696bfb25e11e762838833b3d8b5d0da6e6cfb81814c9ce0005dc78f3dff2b4c633f53d6beaeeaa50e22e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba230dbb982a8abc3b694114981d55b82253428332849167a77e93830078e91a408a0e853964c1851aa847aca4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c9d41ac52f70733efbc61564810dd4c5df581130161ca57af6aeff6a550f4c87b5ae3e2a5b7373d1f665794f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2daaa4294021a40a29a513155c088af60243eece8583265f24fdcc5a33ff55856f22d97a54a49cfd622e0cc557;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40a4c9e90b325aabb76e9672c48e770a551bb3f4add48ec16dae08713925a0632260e37a498f07419b6377f3fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1971196c2f0f6bccb8977c3decd238ce5597c2f64d98a66ad9c4b5f263acc56e6de087fed4196a4c31e8d79c6c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e21fdf815597400878b60a425addb2c31f221baf8f525ca4f55ef8d3848431f2c7cb25f21e1b659958d7a7036;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b4e0aee8c20e6dd7b97a56411389268a1738ca7e5b76bc784dc6670afd60b4e299a22d438880d43f9bb14f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144e2fcb4e18d920102d6da94abf4eae71e77bb9c74f1283cabf9d1576be40a938fbb64fc25a9a3c3bef0cdac60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91b7b1d662f0d1263e0c2fb0ff86473add2f817f39dac884e6162c7b1f12f0479fd6c82c1a79fe092d34dce6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbf88518932da61a2c54407f10ca8bfb1d9a354a2084e9170095999167f353aa254e3d403b97b650b6c96c4455;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de022bf97b8d0ce1c96d4b2bbe9fa188714fbcc867d8931a9bfe02b6464d4bf1cccd0d3ab6643dee08a8bfdc15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbe1b39c1bd207b1a46f8807e740c218d38a79c2709e07eefb543de685e2f55c8c2364b72561149b03031b191f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12015c35858be622f80a593fd14c3c995107281792f73294479fe72264951c9334e64d6402dbc81ab04b5ae12dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf247ae82d8a715ebb89c951c9f16b0cb917176a7aadd0cb330f72d45b5b5e301aefd891fe0d627d23452b52280;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1585df0bc1325ea0869457d483f7cbd40c396cf12d26bcdb0f80171db8442fa22f1fda43786c0b62a6e296a167d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b350f298a6aedfcee5d223251c2957687f8f076a7d202d2c999fec70134116bb31e5dbe810529e83cc7bda9919;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a7799411b725abfd887eb09aafa2c36418e182954ea2a1d0e9e7caa8812e2cc1b21fa36f590f6adaa82731ca0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12fa09d6a1fb0da3ec84605a188e7976ebb2ff40cc9bab8cb4cd4b0f068576aed3f328726ab7f11c35232c01cba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f38fa1c5027989a3eca1beeb3f0ed6c7dc184ef9e754551f981471828d8b696f413b7ea49772858cba495d96b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19228ecb50140c96ae1e6cfc3086833e089fd6ecadb37cb48054a78a08915b4ba3efa3dec6bc76ae54c97fbb0bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h443290bef452cc4044da5b0c1ba70a9837987d92f055e6a7ba347e4fb968758a0d698e0a38c74f08408ba7a3f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed4d60197299594d35c19a130fb3b429b2890270287ea30f5e6abb23f535d9616f8494e86d93e30e3158c576c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7ec43e52f5e45c0866655e90379b425f1572c7d2c332868215616b3a9d36ff188af1b1e21c5a6177e5bca4441;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f64c2d985f8c65993a5e403f374f8bcf384dde0849a70c93982d4077752ee9ef2450435b3737d7185376c95e2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd98f0d6b38730427e099d8624392b544fd07f0202663e52a505439f35e67e86273a5cd663de540f2f4f588b57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c457414626adbf6963d4c7e62088a70a4b1ea2f83e9eddd0619b400381cdf244b604e354b0e56e6d0fcba3337;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa9e2da970b0cd7b6b28cd56b122526229f483d198d523d802aeb55dcb9be377738d7aa9de843541075476bcc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6357f14dfa837bcd806842d2a0c00494783103cac7952ff71c6c1b52d6b0d1066ecc8538d3f18bd16af1d8574b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7cda73c879d6fa5151c4a816bcb0d8847866f3e25675a581fb2452e07763245447ac897287e2376f29dba2c39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111899e413252019c3a290dc9f996d747bc140246236fb5b39360d2795e86f64375885a1fa0c6bb61cdc8c09298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16328dc053259eca54571a86a2f7a0fa2a44f39b35f45ad01084b42a8fccd039352b5160bc21b5ac63ee8dbc20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc030e6eb5400465794a880a9bb66c649e96fc9a29f8ab55f84410d404296be9d69a27d88cfb6eeb6bd76d3c08d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d85c71786d1a8f11f098a7247ac63013f6f27721985c023240f657ecb0b892860723bc0e499b46d0aa200d6db1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159b2084b1d6a6761b52e97e7e0aba3d5ac6177a3a3024f307eca0abc93ec000e5859a72dbf65411fcb53fdb636;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3296fa164fde7157fec5f12b39bbf5b56aceef933083e343502d98832c2d799e9fa93fb4dacf469bd337faad3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb6f56403815a3f072d2ebed1b7be7fb44cf1269922d6b560e56a418c63a7a74ec4cff5c57229b43980b4c2410;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b54297d84ec85c64b149847dd088afe89b27207500d26bb44bba2d9bf112172814e5b8e1e0bd26f0df95f4e894;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h691ac5cc0c88ae06e65096536ba7988523e6b922c42cc4d091b5b6fd6d6176ce6f912d6486544361d221c950d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h21c9e2320cbb44b1ee8b1acab4b0d011d9b6e33a6d384510d43fb1d4184c1db8760d4f700716811f06d18579f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb750671f2b11d33491a150876a39a3102615c048ed87cc9f1b8d01e4a2768cf3e60c91b7f62a9e2c14fc3e51eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6cf546887a711e96cd2ad73dc5e7796c565319195aa4995b6a36d6ac6a0c5e32711ed961129fe9edacb6e7e69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c449049676a9867f3f398f12708c75305543f18e8a2aab0fba176f9e0129518ea133e40f486e80fc1ec85a4a40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d3854cff77822fd3d7f77137b4f1e2d7f74e2d98eec24460186113701de3ef6dd92fd68b2cd48bce282bbf6df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e1fbb76fd4438421cdabf6e6d2475ac306768beb09dc4a022ef4b516b37ed63562fb683ca863788e542f664ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17be2daa741d1bfd6990bf7038e49a0ac333e8cc3fa18a36f1981fe24dea799c076482f61ac4a7e3c04b1c89d72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82dc2db190dc39ecf9e8e71ba67168525edfc1bf398245819f204432cd390c1365ff72ae79dcd60cf2904ffdf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131056b3c6e679aa410ed96fc5d3667da2f3bcc57640ca55e96877e2e1dd9d5385cda0e7d8a02342710b10d2be5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha16c507cf81d5192c41fc6094400ff4d8ac0098c0247ed2127636fbedae90feee56683773d41c0c1d5d45a048b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbb6efce85384aafe0f9912f5356cd398aeb39d97b5d555d7074642c3b4e95b1869fc5ced4e26d3733936eda5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18400deba79c68efab7312f50b51c7b0eb5ca7ee542cfa287e194748ec14d0858ce41b2bcddac78767266dc9a04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc51925376e69e49a508660b28192a405eddfc38c8017845ef2332d4b0215205b5cf3aaaeae3a750c2c8fbc7d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13807af0b4856abfc524d1f0527481fd4169555e0e5d77f8cb061ba2520654d7eba7095bb1954038ecc052d7d14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb4039928cf8a4e49db81480e4b1a5328e51984a479e9de8135481c59c16d696e773fa31abce433ad87550b557;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19231c1c0f36e3111193da377af06359ca6057827d50051c2bd7cbd4ae111c5cb4decf46b9dbd7f450d0038942c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d8f7cb794dde9d79b379455d190e082121b33f3a1e32f1b266425a4a8d643ae382d2c7abdd6db2df76fd5a43d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d112eb2915351018690cd4e9fd7cffa64cc0fc0b48601aff68435b7e3dcbed745bee5bf21278eeacae7d3b394;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3b91c143dc063b9b51372c21e57e466bf9d8623f16704f70ea1c2fcca9a85b7c9fc64d77355edb30ce2682a02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136e3d41ebc5eb805f1ed31fce2c5ce7596e615df8942624dddf24d8f750641545e05a19132abb6fb5c2e84b97b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195e336cc74ce42cf30715e643283b20a04673ea8e70ac2d86d6bc363265fb63615cbcb8ad2287ea6b9c972c545;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1604aa0ca3490240f714bf1f016d68f13234734b30b7372027e109e496602ca5eb0b28ac46133d4e64ccf66d15e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1936812e470ce2722a3d0132b833ea9c408940ce70b9a1e38be126d950e8d08d265844a5b02933fb682a5f7bc88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168519337f7017db82c88d8c51caf639f330bdf266a54de2f7cfdf5c7e03b8c01558976bf858db26ba868146824;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78fd30a39a8bfcea596da4ff0c1b17ccd72282a64c2f88343fb770db395bd760a1bfc48e0aed277f6ee80df701;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h615336a6889a722780e0e03bc777c22c499f9b970ad3b74634a9ae5ff1c8fc2903d5f1b294eebba583ee3fae14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0644023c23b193541edb33b2328ba5f5de1d5699562786981335adf95fdc6fc716ef2f03218e20f5e782224ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19fe14236d4a5b6012c15ee95646f55216ef34a24799be67005d2d302a31a0a0d61644f18b3b78a359bf93c8bb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178152cedb4198ee7a763646ff40930c5a4be694d7d41f72255c1b629669dc769b0c213f710600e5c82e33ea55d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff015091dc43661bbc7b4a66d2cd28c26b0f483bed1329b8f39f63ac5e270abe121967e0bae0c57cc62b0016ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f1c0df3d8059a78c769bece0a57cd380b7b385dcf3d587c17492e257e0b802c09a08c6869cfb71dff622724;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5b094cd2e4fa37d9832bd46bab4b1f2ea810b63324f8ea675ac8e881f38c652809fef6145b30f978a063e8430;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e98c48893c9a19d538d4b4a12feff3a0e545d607a6c11819d5125e71b5aa147771279454ea529c258f8bea6c02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he239613d3797bccd0aa0ce4eea025a595c8ea28616976172db0b8fa895929be3a88496ccb3afb9e80457229871;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7406c024ce3970467db7176b00f041a875ed7863d5bc684e0f4358793bcd202a83b5e4ab25efaeab5e7360927;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8fadd0f1488ae43046b08e0163236070f409c7f2d5b4d17b3f9b167ad15fac4814d93252e9920ad0e3a6bffe0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda88079cc58319d911b2b5da27c02503eb9c5f252ccc3241c344d1e72e624e995d5b36d464d9d4875b62898ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2815ed5c4d23c604f4ed04a6aada94d8ebc22d43d30ace35dba8ffe25c1fc4eaf7f77871ab587de5c4aa33d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f94f48965648e04464e86d9aa638e90d15a46901a04ce4854af935188ffc52936d62032d9e34209236a3108c5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5469f481e5ddffeb08a7d3886a53fbf9aab71ea9d501a765dea8be92ddd2643d8515d783d474e66c0e7fad8fce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h888a511f516cd93f574fd47ff3beb046f77439200eb34764d819f2990e09f0c361b3cfcd37e329feed82d5899b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1162c91e49936ec148671a6636cace12da7a478bf85270d26a4fc365baa44aa43b0e0f3c5165f38cc14d4d3b045;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20c28f4fd27654afb936ea199fc34b0b6b386ad78b1bd3463b9e7be1b06b19ad491499dfbc4b7e43f3b11f6553;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1445a3b6c51eef56daf1588053d27076fdc929d49d4bb5f9be5fb9b2f49efc924016c3eab6df1944e15559c272e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d92d9052664da61e75876871d3423764f63d859878ddc4f4b4e0bb08723ce60ddcf2fdcf800c41e03a5a7ed2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7d17621a58003eb033be9c5d1e89a58347bf50f73b95192cc776c820b8a302ec7bbb146ddb2bb1c2bf736651e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44c4015d54d4f1bca3e684cc896124900f93170388f04d46ad3d436ac7f510af2058708ea7af55db2812ef872a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f1dbb60d6a333ee6fe12d895f0a08110fb9388a62fd375dc45788341df718c18519b8bb46061e295723711b2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178f5a58fd6b38094142427518f4cd1d34bd0dd090417a422d88c15c90cd293356856d1d714aa95f47f2563fb9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h744cad4b0dc14a4efeccf2a753915ad6174b32099e1810374af362834dab2b64729e19dbada574c4bff7e9b948;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14676b24e5c881e8dd144a2728a420bfe810be9731b21482766fe7d72015876febc047874b6bb8c7124bae649ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161deceb78f4fee54df7f8ee7e045633237d981908ba1f01332f88e411a7af9ba5d65905afedf932e438d599cf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7bd0047b6482f656c1c617061f75242eb36526b9d303a26758e01b6ad9c4d38f6a792264d4e9c7486b9d67387a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1266b8e013b1316c8f1af049a37a49986c562ecd0d93e2734fe361886ff1c7440d873f44251af5e91d5c2042c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4672f655d11ec9341b0c2b6ed3dae287ced58c0598ae5231dd68f68b98b0721d296407067e8a8520ad7aa74d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4436818bee0dc093840a898277271b9840f72a36bc9eddd00aaa3c0d7e08067ef7d0dc529a2d5d52e2d8ef9bf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b085d068d9123e903c7172fe9fb92ff290b2ccaea3c67f9126ae615f6f223497b939687a618a27777115451dfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0583298bb71a8e06b75b5cd32789064db4bda40c3c3cf01c86e60e06f8b5d88b29359c66c41c64692d189e4d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3dbec38bc501aa6bd2cd538c72240354ac64a4a32c1e1acb5eb8a4b9faa7bfda114cff56f21cb545fc27e0c13e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfafd26fe535dca4c8682af3dd46ca42a115e8db6930158c77d61abc53488ee3b7fd986b9037bca1d46c3fec782;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb3e08f68a84283688ae8167645e82dc7efec1c1ccbbc5465359e5252fe5b10dc90dd210d4edfc443b29ade35b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe4b77fcefe92684ec1eb45525f2bce6a33e6961739c8a879020d30355e0de1a059b45814a2db45b846b994b0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d866b695b74704c37fb9cee949c6a76cee49f8c41249a19552fc815f80be8fe28224aee5225d97618518bd12a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd263d35731b6ec8e623a46a1682c0fa93af36ecc22399d59a9161ad8925e706f596161708ca6f5e9eff91afd4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1327a7b65cc732f7c80febcc0f0c1c23a16c23b9acd19924a998c08d30d85314387404516f5c91c6296db98637d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0adf92a7f50ad47fa5aa1116ddfeb77ea30975761efd529454210acbbc2f52e2ffcf019ac317e2164ea0d658c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4789f20f6fe317e9997d473849e0cc05f95861ff3625341682171686a5977fe936888b58939376d151aa44fd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55d7f76cd57a03d522d554ea7a4f0bf2268f812d8a0b4b2213adcf09d80d4eaf13bc91045e1474f6c5dd676ce5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78adef6da86b759e3308996f64978f8981ed13b39d81c11475e11913b497c1d7b1fb3bd952fc256c18c6226bf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb0997c0eeee2f217108f594b07bb091addf6e21b4e1810a719173bff057f07b163ce2109d023c3c4dfb906d94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3761b1ebe7f0f414034571ef78db2f5bfbafbf48e974f309fdc9b8dc959b230fd2977fef921dae281453002be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb37877b20861d4214c030726597d47e8b4c09ea797ece5228717b47d26bd251cfc133a4aeea5bfd9e323095192;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156737ab6ce358c2f2eac82fd8d5d1aaf229d07e0bf07c3dfce2e70d5b75f75d2837fc690a9df771048253c6773;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac11b4fa377617161183ec98bb811aba09afc623676122181a1dfea4cb5eb9e6aeac1b7b75e091dd6962cf15e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f3184ef3d1a8240a465aa5ed92d88bb2417d65b7e04774c59d7939561d4ce571307f8e291683873e8c3336e67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb34bd920a8540b077417695c5eaad4067154b94a736b6b060fd37b0d45ef59e5d28548272d8ff725958c73080;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c4d12ea06fa34921b1914d15fb33fc59573056be6801a8b67a4c46e99126961f259dd550106d57c3931fefd57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h867091e7b914caa8e6d10384a42fd296c78261cde68bc6724a1cf564c1b13fbde30da0e01817acb8a525402957;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae3b3c8f58641244ce867e8c6b11373dab7fcb7915a82b51be84a5bef4e7633f98af3cc7f15941faba63729aef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h340a384c15a646fe996ca0eada4b214eeed349b669cfbd312c7c2793cc8ad2c9583e970c92f482586437d6c2f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c74234dbb0b3bd30b51fe26f39cf9f4f0402236f8171e5d78faae3cb9d49474c9b4cc0e12f11f2989b2d0120fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140c079dd7e0ff71665dd5ffa506bfba316dc09042fc2b9fa2baa8f373fb682fecbd4e214fc5cecf03f193df518;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f648127fca55351e3bd797869f1c33ff704d9c558f3ca767e0a27bf600c4292839991e0c1f5065d4639e6c876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c861a0814ebeb57541e588ebc4407b9109fb955a5abf7e5dab0cadc325434df9b2be854a720225133ecaedd599;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bcf5549f0f6d146dad8dbb0c41df15253f6b23706ba81c59cc0fa1f7bdde1fa17c740c07f18e05ca36ce1a1942;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0051ca4f0e05f3accecbb14e32af901a961cd4866380bd611aa1c2876f5a8527b4755bc6d84ac20195c3f5ab7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha82a7ccff02324430fc857f1257116c8960501da079c38eed254a16750e48190502fce56b0f00d9ec62cf60f98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a05cd0aba7e8a2dbfeb633c0d41d5033f805299c41f258aff68ad9f71f55c8669e849ed83098a4d45c903c15f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce5fb0c6c26adcb4eca12c02ebbdd90c26dad71bd24f06b8917b6bb9419350dbce1141913c8ad316cb2d74c10d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0e23d9d8d0b67c1c71035172b4244551666bb18386fbdfc5cb11c5d347cd561d470c6a071b3efb81b8ebf31c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c5bc8e04734055a182c57f02a8cd7114387b5de38896eda16f63ff2ae3cbd4ec69a74f800f8069d4bf8969543;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1847bc58320580eff8449b74641b9af783af5da3d0354f9c6b9ccea0feb4eead876999ca41f762be3a8f80339b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfad3bc3fee90df6aa735bee3c0b7d2019e9e90e9c664e457da09c034d987d6350ede1a6d1c469684a155d5a5ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98537880f58b31e77d5a87acf0346374a386231f5e8b33fa5860826cfb13b5b93317bf2612b68c53f22ce0ee22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18488a4d9970e148c7da8bfc656deaec884ea9046b7040f98770e1e20e7855967eafcc13766545823580ad34afd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0d06bed056ac93cdcc9a89ac030871315580bdaa1e2b27f1b3a47668c37c9ab8b3f6f467eefa47d3eb4699646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e02df610beb2b7f8ca46c174c562de41131c11931b97b4ff7d7c17a8e28520ba778a1e05a0ff9a5a1802e1d97d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69f28b201331ed13fdf02f6b24fc6b16de4f7282627cd45e26c86086e8d42109f72197c3502863a8c190293873;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1525f82d21afc3bf79ad1fb6bae354dab8a67a85f474abb99f1022a459eb974959a8197e42628a6655ca2e36d83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d9c26648e6d38d07f5dd23594eb57e471adae8be400af3ffe6e95e12ec7147dfedaeb3d9110d0503587fbb0c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1648f84063f47a82ae9ead7f2614b986006cdd2e9436d6d5bddc6b638c53f6065cc3115ae30e95a10942d1a9b9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2ecbc6a68b858dc7f379a30bd8940e3f221245147e0c4f149c55b5245e98a471f11652f5fe3364b2540408f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae80862a1d79b0e7809a541587dc00b96a2ee38513236c9d3226b320ecdad58e908724e88825530711e2a69c96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fcc2658ed4283b11de575d29dff36bd27d5d9a5c9e3a8e153700ba9fe41ed9a9b35c0d7298360e40245626072;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be2d355c4175ead63bc052b9013a61876e698c5ec779b189c985898ca45e95406535d5d36a48cb8edfd06d50a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1063a53a06b96353e21c5d0d2632b61503adb6358487cc6685a04c097264863e47abc61697f6e6f6c61743d28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3700f76a1dec0be3a3728d146d4624f2c65367dded4777f4a34a2ea91477d6e538b3731172c8c0970633cbcf5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h304a49510accedf2d1381fa68e3621e12ed6aa1f4dd1490a1de4adcad3d44fe2e4f1189400ce3b0c7f78ccef16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15193a9263cd0f482e23cbba1338edeb2c35afc2a31baf091fc2d0d9b5f8266c794cc53d6ab6f463af6f5be5b3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h410a626e0cec971eb340d55e8ccd1b080aad4f7c3b7ff43aa54fc1a8dac19b1edb5a8bdb9a5a53513cb9a1db97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2705e224b95ddda24d0b9defd900d136b744f10368492ea0a41d132ee7ebd429be88a39f8157658655789858b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha896712477407223562d91cc9e8c49c2d8d5ea67f54f6a5b2b3453c37194fb66f4d9557866f8e188be31e8f81f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95fed617cc7658f94c3ec338fed8ca31d626fd066e26bbeefc266b4a94122b79daf6f13f20e9cb85c7fc519e49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f700bbb8d820180a394c7fe9e328c00ac4a9db3c5770d3aa3a916935442fa6f8ff28d213935fc2e7968b91e739;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17988a30f151e89ff83b5da8491dfd6ff2868e04f3d2e58f2a01bfd5c98997b0cf1d98e699e9db254e21ea750ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha583d3898f7f3920fead5fc8884d6d49fbb6f6c1d2209f5b6d260345958504206194fbf612e3c23d9f7943ac8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bcbfbb45a3eefbf4b6a4cf2111af00d01ce28f71237b73da1de9dfb3075098e36b1af5c33977689fc855c31567;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d96313da5258a52cac5ac36a8d116f4507597c040bedea97d05075e0164521dd0be6ebf2f1c721d0c1877e739;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h702264c2736b5a441a79c8c87569e284b8948a24012e5bd4342687deaa301a92bddc02eaf7efe1da2ab4d1c942;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136398ec734a90f70114af9eb59eb8aa1dacb1b3ba6aff328e092105008b17be1f93f76db0072be4a0ba5a36b1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed8870746e20532284a9e431fffba45140e59f93595d67dec75e2d694181e668286f4df0120ee87417c0fd7a8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e3b412149baf9e5eab5f9dbc62cb29f7dcbbd4c2686bd02dff54ae2d0d6a6c4fbcff5b1596bdd46ebceaf6ba0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4181ba97897e2a24de1c2cc94d7f39969b2203fcf8fe6d7129fa69fced9de136067fc0fab7370b8e844b6d98bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bdd69457cff415d9f44abef504093fd5a29504291041bc77fed35d86817832e7f3bf503fe774fc957031e4f52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71e56b7b176749ee688dbd5b0a1c5f9b7f617887f16063c5e7b156df43027e9604d26eed73b5d6cb315e0597d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b7be3f73d90592e58ab49ec020896237730bfe4e8ee9123a3771cc6e5eb589b6a6654e405bdc5d2e9b908a610;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha627772206f9a3e55d72261be2c610e3cf316d313b038003cbd66a0beef001ffc7869bdc9c509ca2b614cebda9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb04da3b1f6673c4e6f60a8c15412c955598e93f252862e3917ca9e7e3b328c444d1984e20c13ca5569068e9213;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1076234df29704c074db459814e564370a10aceaf260c37df59058df1e01aca1cbddd45e3c2c2746a47e0fb6a94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14804641947e79df30d1a86cd285a789ebb0e6460fb5b0bfae56ff92552a2b960cf4813b0dd0516e3906a8459d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15652b5147a0691eac62b5b111fcbd19c951648bf15289b0982a0be9bc77e62ac1469963f12e090f1fbe87287e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167b8b5eb619e9b7a904bbef0df0c729ce301f1573210af0a7ac5357d0027103eff8c8973d61ccf09475fbd3358;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198bca071343a6551205fed1a3836074c4395bc5abc71235a380f9016e31929f17329ab9f1dfe23c25360efd8fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8c88af69d71248dd04e86ff44a159829e4cd3439a9342df90f693f396ecb84aab374d528f2c9e6290dafd7407;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10258eda2a35f53aeb72a3ddf5930ff31fde319201dd6754d58ed7998779f3225b621c1f56606a0355d68df4706;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdf26aa0deec89abd394fadeea8a6242886470ae01b4988ce3ff6ecf527826c7f8a3d3405f2c7d316f07f7d034;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191778c62efa71fd51b35fec5cf129d372e3f8a1dff5cd09b6215fbd209a74e3fbe8818b272cf65fc67d570454b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c07e5b92bff741daed9c8bc8faffeef3c61fed2c9d2ef722690b1e205c3c30f4909c933af899d04a77a0e62d13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38974b92376f9e04010ad5693fbdd88818cdfd5dcbc11e2d43c0fddf78c3232546f1622c26d44c17859a083582;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heabe852809c696f4672984ee6aa9bed633bf585719f24a4a042f160118945f982de7a1428fd1fc38befefc1465;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165d1d6d6a1d92f11cd14c502cb7b681062867f2e9b9f42769ce07d8e5a2671fc42580a5961019f6d473e2a8953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37364d41a9101c22d0fd46debfbb0bbd0f4391c1a2cae4321e2c42b82436a35d53b1d3d35517b09ce1865a3b58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d1310c811964aa8bdd847ca00c6dd6f506596ada0d2e88a5eae739b9ec7d00f72d54843b01a6ac456e81cd76c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c02d79fa12205ebbdc48f99038bfd8f1dc65b8a8ce65b7ccb76bf06033b1dfa39c575eb1520defc449f8acace9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a51a5931b536dfdcd8a63b6af3f19287af1fedf8ae1b883f0b2653fc994263ad0a838bd64e4c35d72c04c47c1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4af9f035a4d596c28073e816b10447b3f576a1316af4fbc0d62fdacde7d8403e0d9901717e26436b480bbf3d29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7328f2fa944ea87c73d649b6ae909572f7179963069c5a01a68d145e97216aa52408d23c895d27af35df0afc1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ba15b3ec2e4cd5d5a1bd5a9b9892d9e9d59aa1a25138610382144d8ed350d380c9d841ec6d189cc4e62b59135;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88748d0b49ec1c6d8c020e98cfc71ca2d563afaff5bcabda8e3aa1c452c6b32ad5668fc61ca3d324007cba6e19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb887edbca1395d574a2e92694fbfebbae134d9edecbc9363ecaff9ef46bbcd5d8cbec75c0c1365edc89d59de7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19defaabd1767e5d65c987640f77c0d83db46deb6a7b9101737d3f69b286591f72012b6f689a1bd0417a31d3a64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c268091231cf01256b5db0e9a7e47baacba4692c7588e7631215843cd064039d5097a4cc879c13407d30a97be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b9e8ffa45a4a68e91380006ad8f70f9ac120b58b38b7bb010b9d0f57d102717840feadd28ef32cf6342b63c10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166b9a69d6683b9b7208c767182f9515f2dbc3b0566e9a744b17cacda82e4dfdaa8e9331db24b8ba838f43986a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45f233bd49bd24ce969899b630c2606213f17c36041bfa6d8f317e2f4a79781744ffa6060a20865e6d4c29d44e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha03493b0e904d36de00fa05f79f7c33a876a5ed0ecc228a14805daecf10fd9bc3694c7f15888e64d77225aa56e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81fe8098bd8eb8946ecbcd8661dd7de3985d2d6e51980bf37a731349d9281e91c899e59c15ecb33fccb37569b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e43adc62b372d5f40db5bea42f6c399a5f363f689c760df15c3fbb186429c507fd61425c4c86e2ecd40afe0a3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37bd20014c668d0bd42b1a20d6e5a6c3ef82df2a482c549baf8495031e288aaf2c501680686a8c88b1635d1e25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5bc57c07c69eda8f5da4583d89ac23fe67a37218657f1add817fefeb83e9fa0bdae9de58bcb7553aba2c25f8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16313ba0045fa42cd1796f4581c21b11a402b9155c29e9bb7392f98076a22b3bcf03511ac90b64828fdc186b6ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8351298086cba93053a911d0e506e4838e0a3069c41f08469e369415e3d6fccf396446d90bf398107b59a49d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1b84f0a1f1b727f660de12f41dde287b3b471b4ec14e11c48dd15b10eccf022e36eb6b77c50098414c0e56325;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9604ac2ad038e52d93046ad79a38cc4cbc4d6af20247760008f6720270f2545e4856721bac367568447e47ec04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82dc66ed7211ede7a461a972a2ae2242fac0b1126f65023a432d51fdfa5d229f2b9e47290f40025797cf8c80b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h421ef148254f83d4498b05dea06d2ceab9595a487399ffb350f2632bc05d73351cb85e77459469489f0b8e6832;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd232705706912e6609f72e71bf08716429a26e8f42d1af6c21a735d2a2c810f539b151d825a796eb60830e444;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1671bf43f398f80ff605c3d3e11a5061e3f1bba4c3e6298ad8fd358d50d6a785a0e9e09a4836f1b5a449786e289;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6bbbcd7f032dc8136ad1482f4c86603cf59de656162af6734b7564b2edacf0e4b23a2be624dcaeb47c311169e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90418fadd480571a23ca56063ae0c1c21d1c4eab58204e7a92bd53a100192bcfa11572231d778278471494166a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e747d40d580c20b7cfa344c7f2ef5fe82d2e12241dce3fd507b7498098159c749152bd0a689ef3075b09e098;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6731d1572d49534a796677bab967c20362dd4985d6b7a524e40e6664d86de65cebf8a0e760e0d588444ba57344;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb2dd9a43f6439b29939a3265d5793ef3bbfa06c284a0c1ba1f513f754a158e63ceb5ffd74086760e383851649;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16331ba6e944689f4a656e0d4ba836fd5cdcd205a1c06ebe6bc017349a92070de974dde858a3782162bbd826f23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4f55b24cc8f56bf8a7bf7a580ff2b1ccc9ee3f2d36440cdbcd2ca5613127da783a11ef22984951d567c2a6cca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52703b89e78b7e8bc3e248e604c24310fbf335f6dcb00c449fdf7a99e789323eb22829fa7ea0c0f5685af4ebf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h73254ed81d6af91c3f8b191dcc7cbc8211fd29bd5fdd824dc060c1a6ce14202d0987e330520206c36bdbe10e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3a782b59c4fcbd1b79bb61570e373abad468a01c6c2d4dfd524bd3642a4725f55e13f063dd624aa717a6ff3ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ab71f93442e05bc263f332a3c487b31fc3b401f9e4e6085a38439c134fc27a3fd9c589219f08df74acd65e0f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19292664901c8b676f452b16b46ab1a0cbd72a0227c095829f285bfb39a3428696865cff0e51a189252c8c58bb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153e721dd73592e3b83dc770b49b1a34470e569bb23b0ee3555c95b2f625f2323d547d8587bcf4f7ceafa267819;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb3cec8bc93262f5824575896607d4e8bd6d198a7c46eb27513beda3631dbc07a90682ec2a8117d744919d6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14eeb28e650e4e146f348762e33ff48e7e599a45c8857534c031008a876dbf715cb53d7bd501da2468d1e03aefe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1315e23504d5f5896abcb5229793c5230df0a17d97922774c8d73524d6ef3e06f8ab32b332fd40767caa5f45d8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f4b973e9ebf47110db8581ee0524a758fa3816372f5fc21ed43cf4c723e090630a4f12a6e45edbe97e157692a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h800cc5f828222e2613d5a5a423751d67d35b9c544082a7f6c2608efa6986787d33d93ba7ddacbd0306ad5f2892;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b40a28a9bddd3f61ed4bfada5040dc0ae0ba5b523e39b55cc3e47a355f6bf3dc51369e025e360c5bc856e28569;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb2c2724e7464939490239fd9a7538021c0319ec006a552c28e77c7cce74756f53af24d30955f4824d834b1dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2ebaea7d6aa5f01400576c09032c01c4ffcbc84b8bd1174217826e5159dd2932d01aaec6e3a857056f0796541;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10082b0a10d288672ee2b24de54cec244a4c123ad9ed8ff45a3c06fa1966c46b59a8eabe6d0bd6f6dce5cd66be9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha39d27600f1d6a6cbe28e7d3f30faad0d9256bf1fb9b5d203a8a06c2b8d69b828520a19a51aa8b6833ae14bb76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63af734d064075cee2d863969bd4f603af9c957f8a294d94c8b8bf0031269caf73635b8e84c40623b733e4e0b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3b3e7e5e6efd28a18a25acfe40a806cdce8fd5f72d59f9dbe3ad3da8acb343420dd80fe8ca3435e17c2ead5d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152622c972f94daf17028215df5629741fb3b437455441b4fdc84f8f1882d9efa7f68a68c8a56e84d1a0ab2a36f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd349b741ed8f75dcb35b9ad9dbb69c324cc81c4bf30a64c80dc29493281535a59312f05386e088534e7bf5593e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81b6b1e5e4046026545f94c940489042b96ba393e263a78e9d80971157506f94de3b2ee75d745ce6edba1300e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a66e9e1608ac0704e022c42e254f46ca9434a9d50171a61fb99bac64b2c8b43ff41ed488160ced4f7f1180cd6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1134925bd028e5669d80e6b6ce23c2b96d5571c2727429cb399609c930ac7fdd6ca091648164f4613be250f0a0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab83851e97dd7bf8644f14c91ce2fd3a9f8cdaa617e4521a387cd7d5d882d0aec985b52ff3b0c8e250cc4a92fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he56890d4a3b68df2bc255b0f24a1f1c1adee2a7f98d1e894b12f8ec4949f5ad713bb9a5fb1eea7a1aee2050d43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf71e985cb071b750b9899b64503c2dd3677127c8cca15dad5a2a254907e6fd5db87c0d16ca265e0598db85bb3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4033b9b7abd029ad37bb9eac83dd9d75f2121d7993f5b3c15d73a5b4b5895f130d9d518d5904f60e619931c96b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a9312f4ef9d32b2e90b1740811a39ca3d14b93aff467b6e6d6b30891301ac0cc926c2cfe426bd47565d2b0ddf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c80bcfeba00545017f34d9254396e26a0e80e61be4be4cc3526d2f5d43f467ff02a53002108fd9bffc4c622b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haedc31714165a815a78f61e0e1e0e510f3fa8a3d8d7a8ee58107df95b8c8b26bffba18d1a7a2ff38dc2ebebb0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126811fb00b25b1147c6cc2def834d5c54a1066f5b2d0ff8ff2d5327ad8cb6c4c78b7f0ef1bec8748b8aebe49a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124dc3e980be6aae81d7804d98307451275495bdc0b0201111c587918c079b0e5fe878642d8ff4b24121634cd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13074b4da618da62f7ad3de3aeb7ea7909a006f21337141ee7cc0b0f8d78c6be0fa684828c20b4f04f8c5d02433;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18de1a79a256fa27e0411a8ff69bafa13096d506c71cd272d3a9ea125b19f1f984f035bc73a4e05ea8950b87d52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3a1bcf20c4063e190142b73124666846a59c9c075e06ab57763e51de3861117aba7fe11f71e39301164966fcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1795077d05b25e2b57cd78d62b4eeea34d734edf0a90a5c919dcf5aa88decc89948e257fe0ac4bb51e48ba38eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfd55d9728b0ec2b92598ad1350fab848526280305b763bb346948ebd610018e2a24961654dae9fd997327c88f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cf49f3406ef7c93c8f259771e2763548edad4e661297eb8e9f6d3d3e74602bd3d539b551aa98666735156a960;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1387918502cef805c09f7e2df4ae63e0a9d68314b1c1c453cc006bbac878cf1a22bcfb419684c51f85a87cc3079;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50fbfbe5075b5f429ab0efc4de2404918febcb52096a6bb4b318f0ca44aaafcdc96093295f6c4874dd9c0b5ea1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdee95bb1da0fea73544e539055f2b25fb1e78f8f74c688bb582c9894176e23568983194413dfb95800b0565d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e0ab00154552246047fec56797f75641d072623530fdc69bb4a48ff5f2c59128be051718f8ed5fd3f4f7a23fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16342e58164179dd7f646d6675a1351add3688a793a47e40a8bc357e8b33748bb2c9e5eda317f4259ef83821443;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1164447c720304bcf562f29ccd9268bcb26eeedc895a541f394b1f04404ea6cbc444ff2eecc49c7df633a39e24e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdef59b42a805566f57adc241df822f804eb8c62183d708b4c2c0646e4a91a5d20f404e44e722e81ae4a16014e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fec0dc72acd72f945535781c7ce04ade79db0e50b58d31951e12caa31acdf1a78235de3d6fd3c485e062e52e5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fdfc258a8d1114c7ef4cec58e1707b637ea9eff99f739864384c8ce74286e4db21c923f7c8266cd2d363895ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee5c498a855302a7cd1cdc5bb355a9b73b0e451e48a2a2dc72f919a599476629a426a736d66d459880ba5d269e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185fdbe3abf7f4c744fb85bc71aeca57ef79db1e835d9b4368a4d009c23fdf23e2dc07ca542403c998fe4f941e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb55dd87fa428aecffd39872216155891c6ae4024a5d41656b8ab818035b0ccceb7c6a3a505e0c1205dc752413;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17569874d890e3399253177b336ac3b466340e4d469f7eafba6b871a81154b41ad0d9b882ce5b239963acc0a0b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92c128eeca70a04cd58d49362f08b27986445804363662a15c8ffab870da7327d592b0da5370db5d4613c4f87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3c8d938243f33dc071c3e25aefa2c1a6d4a4fc37b94301efa795e3d779b3953fdd0f82f71dc9d65d611f342e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a238dae6ddba7094cc44dbc55fdb53f62a08cc68aab50adf1b7d214dbf9bea14f188987ee905c864e0cbd1b90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde6e961bc74aef2ef275980e413eb4d08280e48f9434bb1acd051e5cdfd92faf110aff450727830f1b2719a63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d462efeaee7ffd6d36bbc1ac7db6e820eb47635caddb514bcb7b8e4a1e6ef080c0df7a7674512455282670d3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28081b239a39877e4e6a59d108be6d5376eb1f34a13cd6ff7f1e4f249045b6dd86ac98a042199540d6e3278ebd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175bb0d8d84e77ddeba95c165b3b1b37a9ee3ae2896b91021ba9eea76b71ffcfc5fb44c0511cd434ad19603249;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c53148c3a317029a6f0b749f57e9c33164669d51fa2dab0c89a9d5e41ffb3719ed398aab3c879decef98726d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef1cf602488a2a802d6a3bb1e32f3db866892b1e05edb70a01d0c52be1ea693e1c6f32a771d6aecee9722a54f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11623bd6375883599529afcacf5d15e2b3acf3173e919df6701b2d8978369d78f0ef98805ef2bf00c176f1aa1ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1075d7e37417cfb902d636c6947ec240d14c7a0c2b2be98c8b26877bda3f7efead1547086b4bca71799f155fae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133533b87661697d96d07e443fbc5b65803214a7ebef484e29e1e568d789d456a5b4d52bf628e985b8a29d9dd5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b17f2dc0561a78fb0b4f457efeaad27e6d9c9db9d0ba6d2a32c317947dbdcd465219553addc8dd9d1c687f5ad5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6768935e4ee9126c7060ddf3b0685ae41338663298c3e9f67675d36c681b955a3202c19265e218ff86200546b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f2d32dca296fef1475b90e6dd154c6d570a38de97c65956c624f90632ff417c76449bded38eece07ad69a9bad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ad61476786994fca1f18c29a7f736a453913e4da9088f691b0feafa9b46a11a97025a4f9b60d7a1c91f80e35a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1edd85767723c9caea4d17d6159e1d7e4e596bb7ec7ec1507f61d928cdaabc10d1bd7a384617a25fd6e03701496;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h353a4c553bb230c0a4b263612beb6acbaa76d5f006e54187578f631d6040efe49785b90a159dbe089c79702ea6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b6dc2b29c8c528d0d7af481accddcc17103f06fc2286f843979b4bf909b6f3fd9e63c91a17ec4282b8b568354;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163ec98364b11b9dc1d59f2edfb10d59ef84d70c706604aa629586ef97e55c39d73146fe41d3e73b0f1f46ccf18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b601674ba5b0c8bb082711b3054d1941a94ddce41870cc99394deb44752ff9822ea301a01a7871dbd7116d84e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2f5003dd30d1b5a4b2e6b52b249cb16c5bad5c97afe7a78f3beb30c43e56a55fd0126b27e5714b80a09ae9461;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1efbd24a0c49a41eeab742323d0a86215d477f600b67fc7cc38ae6c535e7f229b8ce9b2dbffe3833c837df43d56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a0b36c7cb8bd783660de8e7f99f0b56cdd2d2f82bff685d61dba34fa31fb42b7552656e0a62eabef8afa47107;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78a05cdd536b55d8072992bc9fecf864b2e048d42f638196ae9b81b79422ff6d58bde6f605aa3f816bae3532ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1707bbb7946dc417e5abd309c957489f6194e7cb949747fec2b8ea03aaa3082cac1fa678792dbcc606b9d20aabe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65000db4eced32b46ef52422d79f095baddd9172630745473d3fdf013bda19d3e43ea30b43cb2f8cb1e0bd88f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1662163300517313503f7c72ca549591118429d02e935fa8946ac2c1118555b64d0c95c7506186daeaf36bb2dff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195219ad60634e8487ac090c6bd625a7f6e15a0530080e7eabec050f84b42e30b9faf4baf1a4e09fb96011be3e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d71ab82e80b51bc0e41cac6b6c26a52f7696c2796d8f7f57d1b17125026e4f7928097da443b42be272fd411d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14812062d261ce02f5df81b293ae943bc519b242a751c5ff8ddd508db1b46043ca554280f18c884332119b684cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120e71ad6f71e79675f52c46ed78b859a437b38e36e190060390bde449592f679b26652b3eb5b4046e2f328d7b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8de81a5e9b4ee16fa9b6eba26470034b3b3f56f30b90d2c899338c3e53050862d833328233d648890be9042d8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c38cd95b1e250f1ae0cc546de8481f12740705aa3c4dd75978dac8285622715b3652fb65e4e1cc627b40c6b5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b58438f1061c485a1d15bd4e08e058ab2d77e8c831abc7960e739010bd5b02790f53c6f77218ccfc20a344a55f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1588a569ddfc7279cd991cf7b9c8ea9f29bc54738d6dea118d3d6a52ab211184e4c793655606702ba4300ec574a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccdfb0bcc97ab5ba6a38fb45e1f52c40c07e3ad68e0f15bb8739e31d1a2c76bd222b3f48aaa59f61cd2b435270;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1326a014518e617fa13832657616a5d664d989856221c230a473dcb2d5eb78120a50dfa72f7e7fb95d187cd1bee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36ab462ceb52d31affe9eb4ad4bb429f0ace17b9e8f4c3811846f57da7435aebcd1c6c5d6c224189f0d935f2a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c5268898639cbd689f3858f10b49d81f8cbd73cb9888285b5a1479d93aef93034b8b16d9063582bd4bd9a0432;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19636eabb569c9bb62d7b27b482a5518328734f1512897d90fe616d251844b45fa7920bfe03e91d09f85c8e3a10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a883b4f1037bbf9c9ca3c28274eac1cdcb602f99e09587e323a9458c43df8ffc52c5326e2b7384e45619979035;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba6f490807fdc86d8924c1ef2b604ba02a698e65ff5b81f5e0152a8fd6f4ed3bf9e024c60670bcfd8880db83b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148192281cb14a2b0f8ab84fe9f64ffc3441da0f3ecb0588cd3417fc480a948fd714b1fc720494a1562764f6ff6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5bf3da5b840e13556d2023980af340b0cd68872cc3a548bf4548d5bd8c1386e502a03ee6cf5259e5bdf1020b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h264b36e7989857c90a22991ff870f0ad1b6f1673bc83746814675faa214d04ee99cdd7d84ada61c216a9dc1f88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199ebe2e2090b2a2d62c719539a4b2cbcd0d3718eda67b80cb5260aef5e6c409c0b4203e5e768f5216c58d14bf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2269a92d12fce935535e49893cb5dc46aeae07360cbaa08a2e18407cf1db4e3c7fa48fb843eb711d7e1027086;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84465dea27e2942bc1bd21286d59785034833fd536f92b1a67b3a8726c4c010e971fab199232a5966b99323e3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67efcda69eec79419ad987af011283daa5310e94d6a66bee84f585ad9cdc358aae445d02538155e9adcb22c71f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18daecf5a0a1382488f1ccdcfc944fd9c842a67b947be08f43a9671d5f99b59bb4b22e60d4face0f00079138575;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89c181a3187784e6f0033e981e0cc2bdd02fbe0e755a9d59bbc92d3ff4d97366ab213244de18c8f64ab40b903e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ba2a039b747ad06b78bc6bdcc556617d67cdcfddd7a2a16780d35babbf9927ccf5ba32fb911dd5bea50e227f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1317ad7875ac8246645677bb19ac5234e5a2ce26aec631e476f0bbccec7027af963de78b39fd112d5aa48cc7abb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1899d81b920dc5f6063177434fdb1b226186a578e43032ed0af3c30d6eafdf9cdeac2b98a334a1f08720bb95c29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101e85508ef84c06e527fd052b5d7165f4782270c256d5b37c869b398f484852ff485cf6aa35668fa926c7524d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1119d8d8ac8bdad342de4c6ccc1ccfc3b2c92e30d54736fb0d7fe33b0a188c9a7c135342067c6ba5e7c361b2023;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa70c7a12ddc2bd05a373f1cce0d1d9e4eae2fd85887e7f0863864af04fdcc39140bf83f1773ea8e04020932eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffa012180f1a2d399fa28af5cf70d3fa589402b4f9e2c69310f2c31f2da15d3c0cf600b1399868c73a01f9edc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c454701ee83c0be88aceb59f1a4a9bbb2e041bddd3ffaf38685549e048e575cfa7fde00f6b20fec05891b698c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ee1c3f719b361faf22c8d2c615f91cc68d7190616e7283e9e06077ccd9116ba39d83fb3075e5abefe0e12a50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50d214337eb90e34240aa5d3c34037f2e57000ab45276c78344cfab2e62bf04043120c25f4353fd63f049a961f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6cfa4b6bbc0343a62fb73c6adfce2fa8ca38e380d8c1ea6c35c021591d0e8cf261e1b44bf60ce672c2b9864a70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbfdb7cabc574fe5d23246b65cf3acd92bf6de3bc7f9485a45909c90547c0fc4a3e15ce0b959aa0e9a4f2d9500;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ecf85e927210691a2070074c9c7cd2763e1c89543c7e9c384e7124ffc6433942751ddbb51114b370ab5a945839;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1b6efe1adef85b7490c8ebf496d4c0101e7e0ec8c26d7263fb3a89c7b8827881804eaf3df900e6789b8f15e70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9450146bdc2e5290efea5b3fe18ebc67a266a18cfe7b638c5a14851c8fc2264a68da501b14b732cbffbc819272;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf4844aaf13e5316f1510593155b4b3e109c7dc82de876be36b26ad00b60d0f5768e9fabd658327455ed0a436a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dada46edca334635a540fbafe1f516f5bc668865c6fe4f8519d3970ef15ec03f498914149c822572ce65137a04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdeaefb6abc161ff85a88f4c69dca7273c4a7bd2b3c5eecc37c64e99c6844095152ff989c8c73c24ac4e59a85b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c362ee83ba639ef6785c3323ba02ef7858ea526c905640111a691c41199d60e35104603bde720697aba342e3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ff9953ca87fd1991ae6e109f478e77e3e15133424c7c30b81e491339426f71689481c6dd5d050a106460b22d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d4707124d69ad6922138f36a47612c923ea1a6ab46b60ea07d0eb514a3cdd52c4e1c5d1e48ed0bc00c5db3ea1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b623269d2665de6ba4e6f73db433c10d2845b75ee08fd88f70592542cb746cebb425999fa561e7e7bdddd81364;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a19fc021aa8d08ac3a4a712d4bcbf988ff11cd08a903242a1443baecb021a847cbf6360d086d96f3f626c415c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1259e2bd8d87cef20e65e79bbe85cdb1a1541bb97920479ab08477108fd7fa97edd02b9fbc346a2131d496b37c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3367ae2cd443338f0d28ad516985915c59d3422a4721bccf53dd3666e357e86404698cb77097cccc4c06aa473a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1320e42cacfb6fea52411f0ad83a7a79cc81c6f0c8ee9b450fa33be50a9fbdbb4301add6469a951506772303821;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b402fee0679658cdbcdce853670d56f65e38d58cc7712c249a41db99b77d1356cf57f909aad8b7f93ebf6a1bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb74347101c9fcb705f864141354640aa388394d110faa712025c4f47b34d241f49a76d65f5e2d0542577d23920;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ba8061d6b3b54d2da3aa99f16d8bbf902e1cc8ef2fc4cc6b03c465e0e430b276337a03b1c34185c889218b8b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3d44c2f3bd79089b0908ea6401287b53dfefd7aac488210888160cc8fe4d77581611a3888f7cd9738f114fb97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd25160a402f394a92b1629dc98b68a40e434deacbbb6ace0147683f3977f5f0dccd1242387e6da49fe412da1db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2f1ea078f2cf47d6563527dd4283f6206add7f3909cc9734f9e48089bbb0767ee65dc6977a9f83af1ec0f0909;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a56213d705d1ad4de36790b15969ac7f1507540c4f70132bf7266824a80deb747e825fbf00c35d5fdb7941536;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155e8c54cc4cb866030ac5f04249160b02e401b0be32cacad9744a2eec091b94de69c64972c3d032b2a1d710990;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1604ab1232e1c189ef04f9043d39c173d6cacc2606ed30f4eca26b1ae6626eb139b4bd87f55ed4a8c34b30ef261;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a733050ac51a3fe174c05d5d49a12361b9215aab87e195aade8b6b2b5adc7fc72f24812e80e8d60ecd577a707;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4d9815a673376938a10d8066bc3cccc45e789658473e20d522e9b04b406d24e4414105f6cf3ab1bd3a17559c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70c70b1eaab349b510195b0219a409f49878fa06bbfbb0421c88a5cc410fe3e157db8e849262d2aefec17351aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bcce81ba7c66b416cec6575b54c006a74f0b11ef75f6b7c7cfb9d2efc92c6daaec540bd6a434770a44e7126cfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17df0f8232a3715cee1aa345f29dbc908a681dff687647c7f29578a2190a09ba8bf6cd89acba5608a8960f7ecda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc67588ae9864781824fea2c33a8380563c434f49443ecb9e703e449e551abc8ba403ff926790ede7e13655511;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12171d80369af6f48d4e45c58544d74f3f1fe3d0d37b731f1d9670a30e596585fefd2c85228bb828bee7b71750;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1360d12d149bfb4ff7ff937d5f935000fd587aecb935e88091a11df5f8a77f9b59b4bd00df3f600dfc6e2dfc47c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130f564845fb96b5a66216b90b9c0c5e394388a35827bd516c8fd43c1e53b27062da881fb0c2842d25238a0f0fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e173186f5f3f0d60c03b571db70e6b91743c38aa4b4e1b0b730452cc83b61242898c7ca03572bcde1ba645f51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1694137bd3e7aa60fbb3b2f5338ca2ac7572cecc097fe9a75785d7067662f5b10b92cb28c4182998397e252fa2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115d708d8bcb4d352042cf26c8bf73b9dd77510151e9a76493405cab2523ffe5f659822ce269e9ca66ecb4c4e41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18103afc06372e2a2f7220388d4c7eb2e6392f6a8c7036adde64ec64180b488300de081085f4a5168c5d8dcc417;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41d7c8cf8a3a668a8aa236fe2782ebc92535876ac2f11a0979f18e386e7d72414320d82093e1797a174b7f1172;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b80911bfbc6894d2ce680a36f90ad67ddcb97b21dbd3dcd48dc0c147940a0d17179ef9d4e80361960bcd5a871c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha70cb9cd0482cd119aa2cbc248dd7920ff90f7d88eac72e40e610f9fc1f709e0c00b3a9b619c87fc4149bfeb4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc86bdde97f8525cba82cdcbc9a7aae071fa464fc24510160d74eb21a7cede629f861c67119136c8c6f184a98b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134857c64a1f175532d458e4192dac544fe00c3a86cf54e37cba6d6196f79fb983fde2a45529e47a84bedc4aad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdff278c5255e4301bba50db95c5580f7eb35fc6873e93e10bd5ab2edd6ea4c8b843b58871912db9f5e1779a308;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3b5942bb548d075748689bc5f923dd60e6724f28dab925ddad850c5e6c7c7f743706e71fa74bd4ba1723372f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebb4c2dbf672a873a87418b0a860516307e74e2c14e007913b3ee1411770d5c0239193e03c4c09773a87380706;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19670d2bfab00a4c77f313bd161e03b2563414b55e12514b6abacc7fd628dca83fb676ee0620a2a412f3d7de57c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c29907c697c49773c4cf2f33461a7ff71fc800d2f243caa8596d10c7b3686993d5d2aa8159619990b7db016693;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbf22ce5cfc70c4aef35b9d014bf14b75d7aac30f521e3d2c2f6f07f4c831c5f94b7bcbe20f65c772e921cb7d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec11924669963fc611a4bf4dec468fa40da1d4cc4977e4321643c20cf23f4b09d80ba6fb57f6ece499bb5182a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce3a2cea9732e644878c97d0de5859e14d83b66d36acd948b99f4cf1415ee46d262549ac659cd40e4f697a27b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefee132739544be850046d33950fac88d9814bcb7fb303d67794b552294f60c6f1a04df0d01b9818f96c635105;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5974e640ff6fb091247234378e7763a3d7b9ca4e0b94c541c61fe2861d1861fa968cb246ffee5fc7024f9a02bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61d1ddef7302da66029b3f0762bf012073a01407d101d68b6d03c3eb2027e7d40a50afc1453efdd18a19fa9ae1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6bf16c1735093c4930e82cdb5c70bc4b0271c24577a6c32a7f0bd7417a81462955c803e497f7da4ef0e1cdd9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d7401c164e8cf72d53c9a008f1c2c2c0e78df0ed5c97e9db295c785834f02a5dffcc114f80c0cf107c1b266e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7c0ace5595d18db5aacbc578e8f4586e559061092858bb2ff5fecec1dbc5de37756e9814a2b0e9502752aa0f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12fc95d6a0e958b2847e407ed906af55457d424ac6a8045728abf64a62120cd866dd7af0de4d6589608532db014;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc57599cfcf11de24c22863f506a16d6ae76bb843c2667b63d0a7fc2d8d0bce6262c31ad06d83da87c4b0c0cd12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161582d5896483ab771a5e1a07b8146eecfc91a6bb38471b6e869ae4f50a00d466bffe8bdc9f29df38e59e5ba6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1052f34bc03537568dfe89474ed9561743854fce97ffacb0bb5e7e92d7d5a08820fb14d7c8d87262c4009fd79a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b40d8c12584e6e556625c29c2a1cd47fb6924585348ac43b9d4156eb86ce95b953e7ae46c7166c3b1e9d766b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dbb6916687c2ae77577354d7a86d39fd77daa501b4d4b598268e65fccaff9c1adef0701615ce10c53f8019aede;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c50ea4753ed1934d7752efc505988b4d03d4f4c66c2d40fafed7ab7539aa140ca98eb461090d651d64f7ad7432;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1336dd5c846f31d7b19fbef6447c8259005b5ce09ff3847bc0044fcb26313c65e66ee26f03a3a3d5d3e1f9d46a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cd318a739e09171639cc5b906561047240e6e6979ad8f3dbbb21c0f4b981d1c699565698c845bd986a5e5abc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7777932237a7ded8bbd13068eca0a4522eb4d138d8ca35d501f73ccf11710fb9e71ecea131347de7ccddf78c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc155faeb286c61f0d77b982a5ddb601b39d3ce4da27f81af63796b6cc12ddd26c298881dc577bb26423908b153;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14978f71c087f7fcd3878b161a9b5a421cbe4d9bed5aaba1a6df4482f9296828a1bb458d46667095f7f3f264561;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1c5b211c0ebb33ee76de7fb450ef863f858e7855c1c5819ce8e758a514b50b827f990a3a2fe5640f9f9290b7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d34a1cfe37d1a9b6d8bc4bfb930d425e3228ce86517a202793801c20931dcee3b2fecc0e66b1991b593dcd0f17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5b6ddd434a9d45b8a9290d4c60b66659c8a88a23da6505b59970c15188d291a448fe0dd0663a840e3d1f2e0e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c815bb63801a0437ae172b55a1b2575deb5c1372395eda4c4433c55719958fff1a7418576f2dfead512359807;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b28fc0092f6f020828aef6bb05a1e74c7c9fe84c4ba41bb8300d9ec7c04d65a955c25a159b0774c1ffff486ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f18ef0b10a2aa97a2db156857a5964b7cf5e688c052fa39eefabc55aced18151771907b364c0578d40357a439f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1c2e1d2a3d4aecfd92738bbdcacb4a04629031bfe490d914a14323543ad50eef861eab0ec9bf0c1cb8a4bdc2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1ceb0dfbd94df85d4d2758f8e1cb56a146fc7569d598e9c21832b3fda9e8551d0bd38ebcf5ed0451bed403823;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e1ec0312fc865c1b720043beffe2a900da356ea63607a0ec6fb0c11afd4ce219f9a7798b480ea5d74d4eb99b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48959c46c41204aca620824cf3e1135685aa59ed243d21729d2e33050280509c57d228056a550aecb2e10b29ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6cf331731dc5bc1bcce1be378db60957b2439ca320dc426c769cffa61d2f9cc44f62a2cc0a3fa6e259eebf741;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd058a7bce4c07e57b72f7b17960c43d8dd79fd6676b73037aabe61c95cbe74388a17ae66fee074316d3866b70f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acfcb8a71693de193c723ad3ab96fd5786a90d8753834fab93cb835089e9ac10f2e8509a56e29c41334a1300e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf42b12e985dae93b0022695c1b1a7eac6db68c67b226fd386aab64ddba95d931ff31af3ff8046d5431f2eddbcc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8af07e7a8c61cbbbd2c61f60f63dec69a96d04f8bc07d17eee2f8f82e2e7600829d50aee9443f6b69b2faa8ab7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd27d581ffbe4bb061e9552a4db6f0dd73da5e070c4cb250732640365a26fc52ab2a7297ec59eb5798ae1df40fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h606980dede922fa34b23cb935f790d8ad57cd076a61be49698863f24a184342136a14daaac3efa4df805cafbb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1484cae00affd889919780921beb1b460bfd8f7c83c081de872106f4cd2b0346869f8f60bb7ed6f56561df0eab9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f72c42f7a326068e24766d4159600f054358fec41228974a9a56ebeaf821f13a56d30ee69fb643e0c8aeaf3ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9f5def0248e229da44e1bb1fcbbb445be39502911b1a5a2274cc53c42ead8ae6729d03cf98f7a2374224474c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1064bbc6cf106f44ea6841009448f955cafd2d6b096923f20e6234831a6d578eb7d9cc1fded0ab51186b4d4d601;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0a6cd50f33389a66e6b55cef906ce7895c256a2ad78ce4d3c3d5c9e68b331d562038e78abd699d1131d4ec783;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h73cd54e71553a2f3f6ed35f05a16bcc3b696fb8faacb2bddd42f7f7cb09f848a9a92d6a9d649e266a346559246;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c1e3d649df370d9b966884b33e74a7a5fb0a58ae24b211d72937dfdd7b9b6dc2d02dce7d1d3f62b354efb9696;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e2d930305f581367544083de7550dd8c90fb7c21c30decc2d535770feae03ccdd6f3f022bd243268c730dfe05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f785ee914ceaef090cad3e79e3a40360b6d872adcd9d0700b7dc6424e694f2ae13602272e2285eb449debb54e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2244c0c25ddfeaca6c5b5a905f61f964ebb9201e36fbff6edcac290b31796f992807635448aa65d7215317168;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd27640f7423dbc7873a2b26bfe8279c8801d1e5bf6280a4dc992501255c7cf37552fbaa00c5354cc4a405eb22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39f59b79ba4fecf35489486b2c3720ed50b9f4e42cc1135be1f84d0c0772e1c3965046cd43bac52b6fe7ed1ced;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75da27851f1ba0815f1c29bc8dc3dabdae2a3eae2368ec7de5cefeee3297d97a2c0164d4367d6702a16bba5555;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3765d9430f55572bebe91f523cd37e6670ee35a1c41810ea135bbf1a491529b3d92a95f566682f30d48134c63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a2b9f550b37b55247c7c5dbd593d3429883088666858b3329c411a1585cf0e7175192d5d08b3b4cf2cde521ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bd3309ec7b5ce32f58bd955bfb7d953dfa8fd2f6c169de368f0a2ec5a0d6defcb375a83fbf8c8914ca94c31af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c6e57890e647bc77fd216122e2dd3331e331a1287a8ec5a4d7d50601bb98c0c8c845200276f97bd8f0f5e335d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd2b6e6b5cc546a64c6c776921be96ff31a887fa9395d0c4793ddf26185415df6a5f015e92c5a235ab73111b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd9c53c6f50277518f4f385f3ffad75a5695d517f195d8e25f56a112045b5ff6f38f9c1ff387f868ea54a0750e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f719f05a93a389bb1acbdeb3a376953b426f55280843eeb2f159853fbd55fb6e2fcf1313eb8c24085f9a5c02d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b58861e7a03c4ce9ac9ac523548daadce781c00b7e6f64788a0075d81057df3837d590979373246bf196511bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h818f52b3061c223795fdd6465a3cbffcf022954c0e1764858a8257b62ad3742fb8b5b43869572e9210d3f37e68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he879fff3a2a40e4f78e851bc318bd6e56095253448e059f6e8e0342fcf4a261cbed761c5745514956cd019e2dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127522689d8d3d046a9cef224649daf023d2f4593557d1a2882588a82b29f9c61fcfa3e17560a3d23e0dc014820;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea2e8cf2ab7b5e31cd0b5afa76185e08d78c9e6d11e0b4231928deb66c7c7b316b5f68806fb9d3052072c8fbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91b9104c37a159eb77c898fc3ff41ebcd33ac5f751cde19c67f5291f97f09a5b989a51f89d7be6f54b4710e3cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ba98124160325ab5336b92d6b9c65ed9bff6dc5620f6af82b643d3d86fecac4008e688dd826903853bc6bbaa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b567499ebe154035a5d1bad10f84626234dc32a80d6d4ebbbf3712d98de8344f9f3138cd9d58eb50ce2eab7bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7a125690aae5034911376e0f8691a09dc1de3e33ef1cd011f804618e286b8c194e653d384976f6a4c4e0ee29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9cb6a9d1d3657f6ce9c488d8b1b3643ed0c745aec23c82e329d720fe6a1a5ba6ba1537e47efba40e0042a2cb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h517e613c6d4b8c6fad638cf6927c172ba73b5a28ed0ec0ae6919a0e533ebc93fc75dfae0398ac59adf794bb4d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192dc22cef01874389fb48e2b5247ec1f29b8d4226e38c538c80da4a74d6b7c2823dfd6940895c55d3cace01b7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4097a1fc057b550b415475974de4e4da8016956636064ff332042374f032fae225927826d79ea97a4d813c2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e8624ee204a64916974333ca0bbd034e5c565e765f3b9963a8c7566be8b2f37f7084f9d598e97c62908c83094;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e45f40004be752dd6f66f181430a3b734b990786ef1ff7b96adad71cc99cf1529137ef647704521c6214016b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c62022ccbdd74a39d01cd9059764075275f52baff2c42cf75361a47c974ec86380bc2949e4b9e1ad4856270fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e94d47323b81a84427188e8d80333a27692476ad48eacc110e575b5a07448ea25adaad03b6707f30ac8dbe04b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1539aa21ec19f8688a792672915c4d912d8b543d7a124e9e0fe1c39f298b88644355c56dad0883b4772deca3aa6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154bc0aa18a14384ff9b2195fd32a44adaae1541e5bcc4bbb364ed3f8020b44ce0c64d412241521a1f86557868e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h558285ba5d834f5438ddacf6dc16023a3b518fb8a4f49121e47db063fc53bb7e2fa9f8ea3ff6a55eaad280e5b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34d43b41d76c76967b014f4d30c661b73cd717e3e93c2c1283b14890aa6133c05f473c3ae79142553e9e6381c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he51b4f254bbc7fd1f353d3446753063083fcd6cc7f019f6ba2eb01c2d58b9b8e2b1ba0e482c012a24534048db2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1690dd60596c3bbdbd3d87fee6000c45848b4ffb5004417dd19a5a1cc2ce0badf4445831b68fc171004e8dda27a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b83c9802e2cd765bfd5011bdb7216d747b2450b70256443a3236e003ad7149f7cad9b2fbbf3b20877c9b3192f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a9368c74ea155a800e8151ba99d5aac3b2052bfe547479563ced2371b89757dcf4a5f382bf2940cf937642bfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b429855bf3ce30902f01947905dc32eab8f3dad1ad05cdbd57c39a4ddaa50dbcc4506a0f536143356474aa81a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3deb37cabab9393bd9425196213869639e8c34d840121cc5ecc886dcf4546d88df815972c44ec4e4c48878940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f2d6c80bf96fa0e51626a8b9ee7b522265737c88f1394f2e26160f137c38b83802ec1d0dc9efc12ad05ec8a3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d862ac180037ae343bf3bc1ac0d02378cf05c49a536fcb29c4bfcaee279d8d4c9318060dcd6364d7b56202b51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18303b1f3ef5d4f2a1ad70912f42ef8ec86557a661a9a6c0f7ca9ff8ff8bb254d9851344ec747f8c5438d0ca386;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7ce5a15ab201be9e30e2f0d9c405fa6e8d0c4c678df48840efa41f08449845c70d4c65514a77965c16dbb9bee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb76152d075d66a030f932a13921ea9ed9f0b15d3decaa0d62b7928e200e1451a925b48aca07369e56cb50eddfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc3b0997340e561edea700ba6cc826970a4b5fd3d638141ab3ea7c18d191923a0d57663c0bc151b1fb66b55c5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102c4da4b3eaebcc041efc4b934f656f3ca518345a372222816fb2f559974de95a8bccc3df4e6f1e13095ae633f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h331a3b416b71926408585bf14c2563648fcf1b18a7e5ba4f36c77c1c23ccdfbff8fa2b1f255c0609d10810fa8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5d694ee7234142b753297660a6712df0337e388ec03f3768b77185be9e20d214af1762898e1946fd02a453368;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d8ccd9d584f12a90f925bd1448bb6150010e9162203212e050c2b828e70fe032fb697fb03a8642c6464731dab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b89c5c704214280f738a027219cac4c02ea7275cd726bcb37e956db1177cd58a60d7deebf9abbc982ff7f24cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d08d4af33cc7545353841ca9431cbded9ccfa8083c2e4804c4bfbc46ec716e6853c20ad9bd1b9efd3d11f36578;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b1795a2c6e62d021f51452582ed62194ebfa3d8ee1477f9199513c57aff512a7d9a4868cbb96cf501715ce440;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3af3ac2a69519a0fd53d25ab7cfd38f6bf263c9a99d81bd05597c6ac955ee24a44f8e035245183f142e5919c04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h306ffd1ebb8ae6b626ed2eefc4bba53e1ec4c83c86ef4ea2608be6fd99c5f4f3c03e282a754bc716a929e4f723;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197255d2466c2770c35bc46705bbdaff4c9ee591e17b27045d326a14f3f485ebfaffb553331c258aac1fa73b2e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8240cb12bf8542e12e5f89ee191301af8d1d2dfb831f2f2526335c59905bc6e4b87854d2617b9536c0222b0134;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0401623b76252ece62b52c9e72b0cf9334a07d7e009198f087b2871046ca395a3c85232d6745563d46f621b4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1dc9e8b0e3854a29cbd63afa19ea50558de74f2246e3c9e11fdefde981db948b52a5ca084e475ee2e9b45f53d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11df07735f8ebb163bb277d9ed5b62609871b0f84c49886e6a7288d2655a1dbdf6892ffb3d9528faa023cf4be7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b1edf6355e164281e83c2850804a1ffc26e97c61a6fd3ebfaac056b082a0e3c329589f2bbc6946fde7b8bace1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a481226350464c579fd4348287952945b1d87bdb4c9d06ccc74524aae7c19de106a146ddf9596ec5438ca2fe42;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87f16f4791ac0a36da93cda9394ac31e6bf2ef0a0834d8a5f3d0be5081a2c60050ad1d5e9ae2d6c91dd3eb1756;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1799bf88250262cba6269bad49025e1143425e3c2d133992911b2003e5d4f042d21f51a36ef8e4f00ddc423e77c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d60759cf9f6ef081eaa8982d2c3bfa2c609bea580bdd8823a0e422307326148cd77562de160cf8b855aecb9e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca17e6ed8ee4cc257757be986167697cac723b0fa3e35ce247b78b6343682363bfa633603250189954c2e1ef7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ad3e1c133ffcfd681b700b9843706f47e126f771c6495ea7e5f00484db04189f8abe543e6a8659b2976f600d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c25b9a070f10d8cda0005f011afa01f24656b75f8ac47053a1c18e0c640f4c3c6bfec5808e1c5165391fd8778;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a519adeb68df672c532ff415f1e71c3a9693406adbc2493570ecd182c65b8f9ac2ad726c8193096f7bf5af2d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc581d865569d314b109a4ecb8622826d39b500819c1ef466e62ca23fdfcc6a19a90f67447311852a64ff1154c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19503b45bd032a375536f138629f868da10d984dfaef8fee54881dcc92d32075722f557c0f1b89e540b21a74f6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110c4b5f5846267422591f89d8bc40236331ed4eaa944dd85ec636ac43a5212b687d8c203c9b46be391aff02301;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he24fb871e64841a75e7da4e09fbfcd7a51d4c9a8dab387e222a69593e74cfd9029f6e7a12b4297a073bf78d60d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112ae115ef4a1f1da1f002aed2a0c324119225d8f64de745a0f28ee132f98cc4873c5c6d764569c552f24188640;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59443c12da1b9840289a17372a53b91c4fc090bb5934d6c3a7aeab69e967684914dd665e37848d99143d3ae6e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d89c4717a412fcd5609eaf440c40cdacbe82c3d649fd260e9fb814273e540e766a204db63c5fc2d922aa95db2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1861e76ceb1b31919550d73ff06eb7628af98044a8a3bad84b995ceeffbac49fe83c6a19994547766bc7b44ee51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3af5827b8edb2a44d5978e1c132c60205a236af80b0f5b489cf6b231d3df78ae42a244811296852b4766ea344;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h659346cd0e4fedcd0f63a62a706834f43dfb8561dfee6919b21abcf5f602ccd10901b14adc64b7c07cd660e6bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd772976ad2b6231a4743d06207682d813e662f990a43e7e57f2d048f175259e025934ce9956e191c8d7daa125a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b72ef08b1f776463af517b93a3cc33628ca663a9df8393dc65fc3e09694d2119f34170a409f6e799d4d108c5c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1115eeb4fa44021891b38f4c20ec1af0c44a69337033d2aacc2fa0f0bf1641a156beb5c85a398ff343ff0c1c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8a53f157a3d0946b58ee5c4ef38194fb09be179664c34526dd5901e81ea578e6330706e109cb7ae9dab8d199a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3393938bc7419c15a31330d0854aaecd43e70ca2fe1fe2106dce230840803e31d9f53b15dda70017ed54a27e0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7a0c422aea41fe3dd8e5b0259ae04b25055d62d38d1201e35aec73d35832fe0d71a81fbf9474c0dc0def47267;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193ade915d026bfd777e1100bbebf5cb4fce510b73e1484c603e21e5855304b1e080201ea869834ae0599f52d4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86a628e5c976476777289053a1b6c15f0b5b21f5f6ea28cf69995d42ca26d1c446fce9b49f67d5fc4265c3bd32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h803921445ab87be8e87282b92d0b1e7d5a015a7924c062c59b1de49b910301eec3c64d5dc8290d8f8e689ea39c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3dab11eca9365408abe4b1e5242c51713c110e99597f5c2a3923bfc66407ea74096b18f35f351f2b16c57dca0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a63ca9488bdfeb4b601339bace7c1b96193811609d4bbf12491c3ed03c6aa4c0b1146e34b8cb02eb990538b001;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114cfd5542f8325bcaa42da8dd3387e873182cd96271390a60be49b3b42612989a1c302ac35b6bcfea967a6d71a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dcb4b0c3a16e5c6d7a32e9e2e4a870c84318438803c0d576f71881fe23b9714e97fd59c06f2497c2903ae281e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151eb60d89a9d0c55fe884cf2f830a56b196cbabc93d1eb2442199555c667d98c65878ad327d7748793a161a00c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b27746de20f05f536e24410e338d180bc564dc92b03da7b64fe4731168d8e687d151c299872b70c7863b93bda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h809da90fc547c6235bacd7fac7c6719ddc5d1ba87d3447ba85f42083e16e647adeb0eb6130a3e229fdaecafe39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc86b0453cc39bdd7ee486c80c5ae95f36b92806058c829665d0ae134c5561b0eb3988a9a00ce789a7aed1bde82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ec2351150cbb1e1d2c847299effe262b2bc2d8efe689c23e78fae3d480ff677da799c43fc01df9a33b797c69c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66e7258af89c59392a36ca16294dcf7de69151da4c30e1ae22ed2d7d06d70932ada9185a688a20fd82bbe9da9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ec055d0769e2b010c4e04b7b5793b4e9850db1db0ab14e66fcde3b578bc378141278217ca76b2180495d7bda9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87d259ae5ae6bbc8d19269a9b9eab841ec34eafe141731a01f3ae982e42f59b4260a9391686d3c33eb1a0b0442;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h767294e908bef477ac355a2b32516bb19770beb23c8d0339517d465f4ec82f076cbb294556bb202a0c1c715253;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2203ac81bd94c856bffe1b2fb55e8d936905df0c8fce6937e0e83d7ea6c9836c9e7decf0b5b9f53f52a4470ee9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c11512953c252f1a09f2e17d4bf655087b9ddb5056d9783da75577ac073df0d8f92787cb8fa0fa212a5ae8f162;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f9e1617878a3455cd7e9c5a346da7b71a2a691fcc7fc375d215c5e378a8c234b62367884585e1c64b7692c5f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10764720d370936358867bbfa3d3b197f6896d2560e5e5ea25a23572af91e13e913b263f6f897a615f2dd4f0d76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d812a1edd7c04df9d46bb2f510f19499c21b2a19ec691c5fa7af5f54655637c03f974592ddb8b4ccc471a05a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0c3818d9dd77a986718254b05b1b2c4bbdb32dd15b32b5b8b529803cf8aa3bb4567fbd44654ca96c8ebd13ecc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170b707e02b863174058cc1fcfdb5f2dd3ea3cc976555a4a101df2a12d0cbdd3d301d7d2710045e2773ddd93d71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfbe2a8914d1f66b310e219d9aeb7ee48d83f5a0659d8ac07535d2e4d617ee1dd1096e292136ae269a5f88bca51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b70f70cac83768e2f55c7ffed407e73cf83a92fd5a3f7ab6ce3432c32bcd14db1bccddbadd909795acd10679ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f331ce763bc365156a61b503a6b7742ed4142355feb7554b1dc4dbc2bccac519a4c4bb2a141286c8b1bac39ee9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b3444c6df863f469403c23e2efeefc2f31b1309f7c065c831ab575fd7ab3ad2128c15aca9d165a67d1f46c4b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46d84c24b8a756340a7ab123b926ca9259974538b6151a9bb69a84d753248a637107c6107c5c876a2d94b41341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7c8aa080da68d8fbcd204a6b73851d8808542244710296a19d739b49c24a91e9e03c816451cf45b8211eb36b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9135e48da5403ee57ad37320d54edd80ff67b692b87caba8bd1aa9ad074bac2c5148f38483dfaf5cc214a30c9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f952aeaa198aac18ec28111dba382b242042688767f2bd6bf8c11cb59ea94390a1ad91b42d83f898e6f17051f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7602bc2e33d6d247a37a5bef47f9da80d4b0971d3cfd3b68c1327628d5034b70be4ceff334bee622e3ffb9122;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1284a185af0abffcf4b6ea25c30eb6725024ceddc04a85be73da7c7f5c52d31d8c479433bfca758835f49fc50ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b91c31d4d6b668e334cb753aafba4d8806f9ee8b91565686293b082ec31532af0791f08a6d0ab0c03ad3ee2f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae450ffca37e120bd2e53a445b3d1995440ac3348759f3439101340b070f51ed4b1ddcdc101d6c07d8132e6091;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d11fbb357bc4647bbc2c468648700b30003e46af2b74a994efdf1177dd379055a5fd4307acfab21740a17473e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f3f201e740ade2e3cf6f2343cdea6929fa237f68e7ca7bc6148a1ebc7a9bbcd8197b2ae746a0f4651367041ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106e42d89c106deb1f1acfaa619c4d3868855897a663719b7b60003a353ded194297ce9451cae52bae69f882bb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117717764c991abae471af198d128ea57aebf8b68a7bed56dffbfedac2c5a7458be240eea76e7e1a7d460875f1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hacb26141c4436102c0d616792e9982ca67b37ad396fa086d999913ede9dbe146f53113bc2dcd5a278a7990d12c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198e7a13497b8932368426f3814b56ee00896006cdce8e204e27929a756442fdea4670580fc7a83b9cc9c3ddae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d20ff37059f7e8d13a32425b1929736a5c21d79c7cf921d2e0d29ec9280d8e36a9fdd463d67c13f419dbc75b55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ebb4591752fd89edb15e6eb4a02b9f0db2cc97c707c84840dcf473bdaa5d872e42d3cbb8ae73cb68e0674c9a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb2914d84545d1b90943bd9ea2381ce79af890a332925c570b56a57004aaa265b41c65c3d28787f9cd88279ae4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4966bde4ce8defaae865f6bac33681bbb2f8a26baf6c43c47b0aff0b1dad45e7fe2f4d1f6e0404c24fda1d0342;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154db104e2c27a971c865f9e8c4fd7840b187beac1f7751a711d1ae45c97fe4f6c5b874b7904e6100068a0b3dd8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195d63e09fc7cca3ecb1ecd69fbbf306f208a1b18a650423188220441735bee36364909d7b6c62b40e57c26d06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bda88483d68e6b2205a1e6f8c76d6e3ec2d931729fbcf354b2a34364093b6684ac643b5081d0688359714a00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4b2c5f1cf4a502aad47272af446ba6e17d6168e0bbf136c67e393773ddceb9528478fa491dc4bdc73f677fe93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bd6dee7a9aa945a8b053ebb5be67f7442f9d8515b2ab90a4487d9f393a0e12eedc12e10d3fac1c0a04cba5799;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6a7766fbbb139acba2534206060e2154874214cbe7e7bc8538e6530c7118a543873288c967314df8951a1f1d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b41fdde1b12ba2c02244fd56a1efcf7f842360b440b5a56ac1fc143a22448750f59d704f13741fbe14f5616fcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4fc547b9e19e6d31320a5dc77c3fb829d10544959f2e78ce540cd7c349949c8ffd41083a579ed4752f5799f2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1a7cecd840398358ac5ef1d7dd63c5fa087d63065881a55a85b4ab021db8439eeb06cc2a91dd7b87a99fcc34d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc960913f6a6d4c62c481c24a9542c195e0cbf1d045eccee8a17676f4c3851e67e6672743c62111a07f66fb32b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1871f448b6cf8cf81cfb7885d2d3a2ea71086fe9177b5d230043d4c6397164703ff2cd430c123c6307e723fa704;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee75e8b7969b007e55bf9a7f5dac89b31f0a790b4da0a9a55b1783f4d08dacf0ebba9fd7983734220946bcfa52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eebbf0bded07ac1df89fffd50bac85d2b1feecc9950aed0c4524b6d234cf54563bd9e30971f40a9dc8f9dc1fd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17257b18e78aa61b6bd6d3cd387042a4a148f71fed6e331dd90025984d7480b9a04298413bece0879f4a9dd202d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0fd5119816b2bc3377e64358bdd6cfeb01c9d2a0600dbc1501019dc6acc2925996a2f64e8ce25b8870c07681a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb444ac08f7a0d4ae67b3d9d8a0bc68450c772c7a2793def94573ae6f55c3bcb9cf98830df08417ffd4886fa86d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9476c810de97c10515d5721fd4814994d68dcb2fcd6fd9697928f63fc1a3bc191770bd001a44ab054dffd58f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1624eef2c18de0df904b603d6cbf8705b2b06380587ed49ef3abeeb27ae205d0fe40b371099315b515d9652d18c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3d7b2402c8d54f8dd740706fe46b07b65d0570570c60cc888a55d36d1e339f7c2b3e49236ba1b9c4a9a70f87a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196836c9f87cec77af3912b249aedf4901a39a3c196b37e0aa8d07e216a830ea82caf5d61119d31eb4e9a2c3621;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50610ba9853bfea68d753798f47939d4f0efa524d81d4404903e4eb8ba9b5e6addc64af8470a951455090452ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haecd48742bba2f9841d1c5bb4b8ff16fc5ce33af55fcb72347b877feb7debd06f807fcdb3d737b0546f4a40d2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he855e3324f799c772578e61d1f8bd465e3138ebffe8aa8bbfc9af894170f3d340ca8f23f72bc43220722ee714c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6e376e5d60b0ce38b419c8b86132221904c4d32787c72a3d9408950b92727b7f70cff5861d6ad31f346b600b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8510125391b511be95db9a3db3e4115c85c02e6153c670170577213cd4a76e51c87e857973aebec30596e322d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h314a676efc2452374cf1f5dd0552afc5c687e81526cfaeb2e022638b4bfb91a8f76e6330d9ad67542684f915b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bac46a802143a913106e4b2ae6c635c8a63c6a4c6bcda8b51b6d4f45c4e8f63e3dc212f16a09ee96e8c392242;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165e7c99995590189c4af4d6750878eec581274be1681664d62b335563a818d362f275f6f2c4bdef051aee40b9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d71c0f270692c9a44018ec411c9a30881448d74d1af32744e91008b9d2c22726b86d4e7e21cf4f7407a4d9c013;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe939e55f6693cbeef9d0895b132290cf366bcfbe2512b82ba29f828271c0755f00a65a920ccbb4f6e35f5a641;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he019b5a903a2b30c068543673a9df54f279f40adc7afebcca52ae512cc550fb3c4936d3b17534808e3247a311f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf945411ac1856edb040c260edd711d1aa130aeee2cc26da392f7797940b36f1f02e1c342d6186fa6c34c0fedfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47b536c59718dd944ad3ba5f2984a362c9c14f620d4914fbb28a3b0834434363d283d06763c5916c1bc54ff045;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb383aa89273d865268125a23b8064eb0ca4ea8a546246cdad2c7661ca19e73ddab88fd4a56c83486b53cd520cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108e64115815a9388e9ab3cd7460eb3cdc33ca3fdb9fafcaeb38a86bee24b769da4c0450bbf4d26feed3bd96398;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10aaf203780409e1828060a468425b0b36b143cd2847ca5b2ac6af8f9ab28a878d54edd781d38b46f5e4498509e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebe796566bdff56e80ada3025d815e1947c76476235b6b91e0c9960bb65fd590596a875a773fa38877005995a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d0b28229bee9087507bca1b492eb0cc15bcd0b00f0aeb79940679a2902589d78244087d618a488f2573cb43a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17022c71a5936a0f71774828fadc737e55370e295bbea93209a700530d92f7a81574de7da29d9e996f76800275b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hceaea62263c80f2521e62f48f709f1016be9eccf56185a8941a11c23865675760919bb0089500a8dd216f6184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199ed83f0228bddff24a823338f6e9f9a091b5da66f2d9e973cab9a0aed53c674d8597af5a5fd9a3c6e4638d940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h643ca2497582d057c7d7ea7f0a2cc16581dd5e84dbd8f585919378d16c4671002c7a731e515d611e68b7924db4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7f389f0ff26890e9af459d5b7155a91392bdfefda0bcb8ce41b2d75fa24d95a1f3091478ae87c5cfbe744a45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8324ec1d465cfc588e72d28cc3883e17e421ff2007172fd5f4a150704104bf0a2be7bdd1e8be6f9c04d1413b46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ae9bd96b2cfb647c2bb901993227d6bbcb0583d6cbae4d0810ba4a47c743d89d1ab1eda5a6c7fe253bdbff392;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a1a0e0cb88a98d4613c3ccdec5758533cbb0a7eb6fbe682f422b5d1aae20ea2f408e1cbf39820837367b2779d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa17efa203f87d67053524ff104e6871fb8cfb27bcc5725ceb65f7159bad7da33cfab9eec71eb786b21ca3fd95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5992c002640b8895a89657d8cfa90661f61923a7cb0981a36d7b0b26cf7ad8fe5d7eb07c6f1cc690da6b36c76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34f445a19d1239c5b30d1c35150491eb17e98fa6667ed1b36d3ec701e1817d00dd73be7053453f19426e6d059a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4c921df6ddda51672b9cfcbf8268f46e712f20a55e56ea430ebd77b608fe772c3e73feeecb8439ae94a5b914f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141b49b28bd4c5cfd1cfaa251edd62410456a4a5c758ad6249fe70ace6a09ea16c56111d04d4db2ac51edeafddf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4dc695ccff7ff955b8905628c3d38b8319d9dcabc6eeed359b082fb5110a963d4013fc85fc1120580b852e23e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100185d536327bad052068e1b567617772142c70c0665a44cfbccb4bf1d252f753182be47b33ab2b7ca1800d656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17574ff2884acfb9dbe6ec2e3e8ceb19fa138fed85e1a42d272192c16ec53dde5c870ab857cd15ed87141adcde1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160d24e43d3ad1b09dd09ad4f6cd8f5eaf3b5ec4854cf9b6eeaf903367b35f1d8f122c84b8a0e5a69c69e7f2624;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb5f58a9042e1d0f4155982d257b807494e0be0f79a30182a0fb0308982228e10a447bc6610ebebf51ba9c782e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163b1c35d4a1ecc2d10f38b428778499a3f2461c7c8457682f103f246074c9a5376bdc2d14d0ebd9f10779043d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ed64e81231074a9d54dfec61ac97666bcca6e846f8617468a9b2c47d2b034d4453a0973f0aa354eeca0c44fb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha64a339884922cdff535c0c3ddd7b6ed0732e8f7469f6dc0822c8d320f7b70dbfcb242946949395bf11fdfcc7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c3aedb2e46202d7586c8595d65a414d7f6798fed4230380f135b57489f36e1cd0fc40355ac7f4604862bd677;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138cec8dadceca69908e326a63d67f963d94142093ac4310da74c2992e042070ae499ecdcecff3ea01c7612946c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14cc59b010d17d2f59f5f0fc1da743dd291b49bf6aa458483e4318cf00c4dae29b9f63e080451584dd912601956;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bfe27747b27f218f31451d2ee1ab52be49a876fd615bc823b46ca0dc7617e0808e7d14cd2deb010fb886eabc90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142d349bb4f90a55d10e7450504eeb27daa576704600920c0832672329e3a8615e246c9f7fc9efc6cd03ea5fa4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he47939f7f9492efc29fe8f489b33020b8a8b93c752da243836c76a0df3b12c4b34cee9b6a847a50157b63c9a76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac41f289199b3bf7245e40a579a51493346b851a0e1c6590352864ab99e7405a9729d3e432ec4aa5d0e8ceeb02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143008f46daa738b1565f8e561a444ee7d5654b39af785c3f865deed5363d9f6c257028c05dba7beb04c71c9ee4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffdf88832736a8ad0f3722d8992295b14a0be5662b3e6090114bb3c47f78b9df2d18a8646a0363f6474d162f05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2fbdd75e6fa9055dd63750e765873a389a4620fe71c850bc264674c644ead44df5353811de340e341eb58b819b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdedb6a8bbf7410c0daaff910565c57e676cd8ee99ca30905360214301d69cf139652436b5cc85c203833f3519;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed002fb050e7a1ab100b25ac62872bddf59ca2b8e313c63f34460df6a39780cf3140a7d274b1e03cfff0d1d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14772d8b137f761a67422c5ee80f3466dc5b9d8e292d256ddfad51f04737375645da4699d881679ebdda1d183d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb68c62514abea4342387b62d85cdae56b3dd0eb16b1028ee32c09be4af8d3746da7d386a9cb5e295367768846;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda860c71b8a72bf4a4331df64dd7a177dd2c4a1030ec0562b7f03495499ea89862a6358005012d6b6de90b7be5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c7f226527af9020d20e20030fa3171e770b8b437f8a9ecfb5bcf248d64bfa0f450e36a122597d81bed3ab4d78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed705c80dfd3cab8fafd117d8ddd64831f13854803c0d2bbbd316cf2789ec5f5de485530a7089ddb762f0cdcd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fe0ae58dd56067adf4765367ddd0e6da9db70c4702e35928d7b185c05bdf066ce393ab1f3ca026ddb6044677;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29ce94df237898c3667be6b0f8136598c32af57013595db87760fecd438ab40231b6f20bc476ba85e24d8ccc76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb68054a9fbbe2f332efb019d88ac8f27689921814cc25db42b6ced6a3480bc11267fcce71f62b97fd7ce4a5315;
        #1
        $finish();
    end
endmodule
